module tt_um_alif_dual_unileak (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire params_ready;
 wire spike_out;
 wire \system_inst.leak_cycles[0] ;
 wire \system_inst.leak_cycles[1] ;
 wire \system_inst.leak_cycles[2] ;
 wire \system_inst.leak_cycles[3] ;
 wire \system_inst.leak_rate[0] ;
 wire \system_inst.leak_rate[1] ;
 wire \system_inst.leak_rate[2] ;
 wire \system_inst.leak_rate[3] ;
 wire \system_inst.leak_rate[4] ;
 wire \system_inst.leak_rate[5] ;
 wire \system_inst.leak_rate[6] ;
 wire \system_inst.leak_rate[7] ;
 wire \system_inst.loader.bit_count[0] ;
 wire \system_inst.loader.bit_count[1] ;
 wire \system_inst.loader.bit_count[2] ;
 wire \system_inst.loader.current_state[0] ;
 wire \system_inst.loader.current_state[1] ;
 wire \system_inst.loader.current_state[2] ;
 wire \system_inst.loader.current_state[4] ;
 wire \system_inst.loader.current_state[5] ;
 wire \system_inst.loader.current_state[6] ;
 wire \system_inst.loader.shift_reg[0] ;
 wire \system_inst.loader.shift_reg[1] ;
 wire \system_inst.loader.shift_reg[2] ;
 wire \system_inst.loader.shift_reg[3] ;
 wire \system_inst.loader.shift_reg[4] ;
 wire \system_inst.loader.shift_reg[5] ;
 wire \system_inst.loader.shift_reg[6] ;
 wire \system_inst.loader.threshold_min[0] ;
 wire \system_inst.loader.threshold_min[1] ;
 wire \system_inst.loader.threshold_min[2] ;
 wire \system_inst.loader.threshold_min[3] ;
 wire \system_inst.loader.threshold_min[4] ;
 wire \system_inst.loader.threshold_min[5] ;
 wire \system_inst.loader.threshold_min[6] ;
 wire \system_inst.loader.threshold_min[7] ;
 wire \system_inst.loader.weight_a[0] ;
 wire \system_inst.loader.weight_a[1] ;
 wire \system_inst.loader.weight_a[2] ;
 wire \system_inst.loader.weight_b[0] ;
 wire \system_inst.loader.weight_b[1] ;
 wire \system_inst.loader.weight_b[2] ;
 wire \system_inst.neuron.leak_counter[0] ;
 wire \system_inst.neuron.leak_counter[1] ;
 wire \system_inst.neuron.leak_counter[2] ;
 wire \system_inst.neuron.leak_counter[3] ;
 wire \system_inst.neuron.refr_cnt[0] ;
 wire \system_inst.neuron.refr_cnt[1] ;
 wire \system_inst.neuron.refr_cnt[2] ;
 wire \system_inst.neuron.refr_cnt[3] ;
 wire \system_inst.neuron.threshold[0] ;
 wire \system_inst.neuron.threshold[1] ;
 wire \system_inst.neuron.threshold[2] ;
 wire \system_inst.neuron.threshold[3] ;
 wire \system_inst.neuron.threshold[4] ;
 wire \system_inst.neuron.threshold[5] ;
 wire \system_inst.neuron.threshold[6] ;
 wire \system_inst.neuron.threshold[7] ;
 wire \system_inst.neuron.v_mem[0] ;
 wire \system_inst.neuron.v_mem[1] ;
 wire \system_inst.neuron.v_mem[2] ;
 wire \system_inst.neuron.v_mem[3] ;
 wire \system_inst.neuron.v_mem[4] ;
 wire \system_inst.neuron.v_mem[5] ;
 wire \system_inst.neuron.v_mem[6] ;
 wire \system_inst.neuron.v_mem[7] ;
 wire \system_inst.neuron.v_mem[8] ;
 wire clknet_0_clk;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;

 sg13g2_inv_1 _0727_ (.Y(_0085_),
    .A(net106));
 sg13g2_inv_1 _0728_ (.Y(_0086_),
    .A(net165));
 sg13g2_inv_1 _0729_ (.Y(_0087_),
    .A(net158));
 sg13g2_inv_1 _0730_ (.Y(_0088_),
    .A(net112));
 sg13g2_inv_1 _0731_ (.Y(_0089_),
    .A(net167));
 sg13g2_inv_1 _0732_ (.Y(_0090_),
    .A(net154));
 sg13g2_inv_2 _0733_ (.Y(_0091_),
    .A(net169));
 sg13g2_inv_1 _0734_ (.Y(_0092_),
    .A(net192));
 sg13g2_inv_1 _0735_ (.Y(_0093_),
    .A(net102));
 sg13g2_inv_2 _0736_ (.Y(_0094_),
    .A(net4));
 sg13g2_inv_1 _0737_ (.Y(_0095_),
    .A(\system_inst.loader.threshold_min[5] ));
 sg13g2_inv_1 _0738_ (.Y(_0096_),
    .A(net201));
 sg13g2_inv_1 _0739_ (.Y(_0097_),
    .A(net213));
 sg13g2_inv_1 _0740_ (.Y(_0098_),
    .A(\system_inst.loader.threshold_min[0] ));
 sg13g2_inv_1 _0741_ (.Y(_0099_),
    .A(\system_inst.leak_rate[2] ));
 sg13g2_inv_1 _0742_ (.Y(_0100_),
    .A(net161));
 sg13g2_inv_1 _0743_ (.Y(_0101_),
    .A(\system_inst.neuron.leak_counter[2] ));
 sg13g2_inv_1 _0744_ (.Y(_0102_),
    .A(\system_inst.neuron.leak_counter[1] ));
 sg13g2_inv_1 _0745_ (.Y(_0103_),
    .A(net205));
 sg13g2_inv_1 _0746_ (.Y(_0104_),
    .A(net215));
 sg13g2_inv_1 _0747_ (.Y(_0105_),
    .A(\system_inst.neuron.v_mem[4] ));
 sg13g2_inv_1 _0748_ (.Y(_0106_),
    .A(\system_inst.neuron.v_mem[1] ));
 sg13g2_inv_1 _0749_ (.Y(_0107_),
    .A(net212));
 sg13g2_inv_1 _0750_ (.Y(_0108_),
    .A(_0006_));
 sg13g2_inv_2 _0751_ (.Y(_0109_),
    .A(\system_inst.neuron.threshold[6] ));
 sg13g2_inv_1 _0752_ (.Y(_0110_),
    .A(net208));
 sg13g2_inv_1 _0753_ (.Y(_0111_),
    .A(net202));
 sg13g2_inv_1 _0754_ (.Y(_0112_),
    .A(\system_inst.neuron.threshold[3] ));
 sg13g2_inv_2 _0755_ (.Y(_0113_),
    .A(\system_inst.neuron.threshold[2] ));
 sg13g2_inv_1 _0756_ (.Y(_0114_),
    .A(\system_inst.neuron.threshold[1] ));
 sg13g2_inv_1 _0757_ (.Y(_0115_),
    .A(\system_inst.neuron.threshold[0] ));
 sg13g2_inv_1 _0758_ (.Y(_0116_),
    .A(net104));
 sg13g2_inv_1 _0759_ (.Y(_0117_),
    .A(net108));
 sg13g2_inv_1 _0760_ (.Y(_0118_),
    .A(net144));
 sg13g2_nand2b_1 _0761_ (.Y(_0119_),
    .B(net145),
    .A_N(net1));
 sg13g2_nand2_1 _0762_ (.Y(_0120_),
    .A(net181),
    .B(net106));
 sg13g2_nor2_1 _0763_ (.A(_0012_),
    .B(_0120_),
    .Y(_0121_));
 sg13g2_inv_1 _0764_ (.Y(_0122_),
    .A(net134));
 sg13g2_and2_2 _0765_ (.A(net1),
    .B(net3),
    .X(_0123_));
 sg13g2_nand2_1 _0766_ (.Y(_0124_),
    .A(net145),
    .B(_0123_));
 sg13g2_o21ai_1 _0767_ (.B1(_0119_),
    .Y(_0125_),
    .A1(net134),
    .A2(_0124_));
 sg13g2_and3_1 _0768_ (.X(_0126_),
    .A(\system_inst.loader.current_state[1] ),
    .B(_0121_),
    .C(_0123_));
 sg13g2_nand3_1 _0769_ (.B(net134),
    .C(_0123_),
    .A(net166),
    .Y(_0127_));
 sg13g2_a22oi_1 _0770_ (.Y(_0128_),
    .B1(_0126_),
    .B2(net144),
    .A2(_0125_),
    .A1(net104));
 sg13g2_inv_1 _0771_ (.Y(_0004_),
    .A(net105));
 sg13g2_nand3_1 _0772_ (.B(net134),
    .C(_0123_),
    .A(net156),
    .Y(_0129_));
 sg13g2_inv_2 _0773_ (.Y(_0130_),
    .A(_0129_));
 sg13g2_a22oi_1 _0774_ (.Y(_0131_),
    .B1(_0130_),
    .B2(net145),
    .A2(_0125_),
    .A1(net150));
 sg13g2_inv_1 _0775_ (.Y(_0002_),
    .A(net151));
 sg13g2_and3_1 _0776_ (.X(_0132_),
    .A(\system_inst.loader.current_state[6] ),
    .B(net134),
    .C(_0123_));
 sg13g2_a22oi_1 _0777_ (.Y(_0133_),
    .B1(net128),
    .B2(net144),
    .A2(_0125_),
    .A1(net166));
 sg13g2_inv_1 _0778_ (.Y(_0001_),
    .A(_0133_));
 sg13g2_nand3_1 _0779_ (.B(net134),
    .C(_0123_),
    .A(net150),
    .Y(_0134_));
 sg13g2_inv_2 _0780_ (.Y(_0135_),
    .A(_0134_));
 sg13g2_a22oi_1 _0781_ (.Y(_0136_),
    .B1(_0135_),
    .B2(net144),
    .A2(_0125_),
    .A1(net152));
 sg13g2_inv_1 _0782_ (.Y(_0005_),
    .A(_0136_));
 sg13g2_nor2_1 _0783_ (.A(net108),
    .B(_0119_),
    .Y(_0137_));
 sg13g2_a21oi_1 _0784_ (.A1(net144),
    .A2(_0123_),
    .Y(_0000_),
    .B1(_0137_));
 sg13g2_nand2_1 _0785_ (.Y(_0138_),
    .A(net156),
    .B(_0125_));
 sg13g2_o21ai_1 _0786_ (.B1(_0138_),
    .Y(_0003_),
    .A1(_0117_),
    .A2(_0124_));
 sg13g2_nor2b_1 _0787_ (.A(net136),
    .B_N(\system_inst.neuron.v_mem[0] ),
    .Y(uo_out[1]));
 sg13g2_nor2_1 _0788_ (.A(net136),
    .B(_0106_),
    .Y(uo_out[2]));
 sg13g2_nor2b_1 _0789_ (.A(net136),
    .B_N(\system_inst.neuron.v_mem[2] ),
    .Y(uo_out[3]));
 sg13g2_nor2b_1 _0790_ (.A(net136),
    .B_N(\system_inst.neuron.v_mem[3] ),
    .Y(uo_out[4]));
 sg13g2_nor2_1 _0791_ (.A(net136),
    .B(_0105_),
    .Y(uo_out[5]));
 sg13g2_nor2b_1 _0792_ (.A(\system_inst.neuron.v_mem[8] ),
    .B_N(\system_inst.neuron.v_mem[5] ),
    .Y(uo_out[6]));
 sg13g2_nor2b_1 _0793_ (.A(net136),
    .B_N(\system_inst.neuron.v_mem[6] ),
    .Y(uo_out[7]));
 sg13g2_and2_2 _0794_ (.A(params_ready),
    .B(net1),
    .X(_0139_));
 sg13g2_nand2_1 _0795_ (.Y(_0140_),
    .A(params_ready),
    .B(net1));
 sg13g2_nor2_1 _0796_ (.A(\system_inst.neuron.refr_cnt[1] ),
    .B(\system_inst.neuron.refr_cnt[0] ),
    .Y(_0141_));
 sg13g2_nor4_2 _0797_ (.A(\system_inst.neuron.refr_cnt[3] ),
    .B(\system_inst.neuron.refr_cnt[2] ),
    .C(\system_inst.neuron.refr_cnt[1] ),
    .Y(_0142_),
    .D(\system_inst.neuron.refr_cnt[0] ));
 sg13g2_nand2_1 _0798_ (.Y(_0143_),
    .A(net2),
    .B(_0142_));
 sg13g2_nand2_1 _0799_ (.Y(_0144_),
    .A(net2),
    .B(_0139_));
 sg13g2_nand3_1 _0800_ (.B(_0139_),
    .C(_0142_),
    .A(net2),
    .Y(_0145_));
 sg13g2_nand2_1 _0801_ (.Y(_0146_),
    .A(\system_inst.loader.weight_b[2] ),
    .B(net9));
 sg13g2_a21oi_2 _0802_ (.B1(_0146_),
    .Y(_0147_),
    .A2(net8),
    .A1(\system_inst.loader.weight_b[1] ));
 sg13g2_and4_1 _0803_ (.A(\system_inst.loader.weight_b[2] ),
    .B(net135),
    .C(net8),
    .D(net10),
    .X(_0148_));
 sg13g2_nand4_1 _0804_ (.B(net135),
    .C(net8),
    .A(\system_inst.loader.weight_b[2] ),
    .Y(_0149_),
    .D(net10));
 sg13g2_nand2_1 _0805_ (.Y(_0150_),
    .A(\system_inst.loader.weight_b[0] ),
    .B(net9));
 sg13g2_a22oi_1 _0806_ (.Y(_0151_),
    .B1(net10),
    .B2(\system_inst.loader.weight_b[2] ),
    .A2(net8),
    .A1(net135));
 sg13g2_or3_1 _0807_ (.A(_0148_),
    .B(_0150_),
    .C(_0151_),
    .X(_0152_));
 sg13g2_o21ai_1 _0808_ (.B1(_0149_),
    .Y(_0153_),
    .A1(_0150_),
    .A2(_0151_));
 sg13g2_and4_1 _0809_ (.A(\system_inst.loader.weight_b[2] ),
    .B(net135),
    .C(net9),
    .D(net8),
    .X(_0154_));
 sg13g2_a22oi_1 _0810_ (.Y(_0155_),
    .B1(net8),
    .B2(\system_inst.loader.weight_b[2] ),
    .A2(net9),
    .A1(net135));
 sg13g2_nor2_1 _0811_ (.A(_0154_),
    .B(_0155_),
    .Y(_0156_));
 sg13g2_nand2_1 _0812_ (.Y(_0157_),
    .A(_0153_),
    .B(_0156_));
 sg13g2_nand2_1 _0813_ (.Y(_0158_),
    .A(\system_inst.loader.weight_b[0] ),
    .B(net10));
 sg13g2_and4_1 _0814_ (.A(net135),
    .B(\system_inst.loader.weight_b[0] ),
    .C(net8),
    .D(net10),
    .X(_0159_));
 sg13g2_o21ai_1 _0815_ (.B1(_0150_),
    .Y(_0160_),
    .A1(_0148_),
    .A2(_0151_));
 sg13g2_and3_1 _0816_ (.X(_0161_),
    .A(_0152_),
    .B(_0159_),
    .C(_0160_));
 sg13g2_nand3_1 _0817_ (.B(_0159_),
    .C(_0160_),
    .A(_0152_),
    .Y(_0162_));
 sg13g2_xnor2_1 _0818_ (.Y(_0163_),
    .A(_0153_),
    .B(_0156_));
 sg13g2_o21ai_1 _0819_ (.B1(_0157_),
    .Y(_0164_),
    .A1(_0162_),
    .A2(_0163_));
 sg13g2_xor2_1 _0820_ (.B(_0164_),
    .A(_0147_),
    .X(_0165_));
 sg13g2_xnor2_1 _0821_ (.Y(_0166_),
    .A(\system_inst.neuron.v_mem[4] ),
    .B(_0165_));
 sg13g2_nand2_1 _0822_ (.Y(_0167_),
    .A(\system_inst.loader.weight_a[2] ),
    .B(net6));
 sg13g2_nand2_2 _0823_ (.Y(_0168_),
    .A(\system_inst.loader.weight_a[1] ),
    .B(net6));
 sg13g2_nand2_1 _0824_ (.Y(_0169_),
    .A(\system_inst.loader.weight_a[2] ),
    .B(net5));
 sg13g2_nand4_1 _0825_ (.B(\system_inst.loader.weight_a[1] ),
    .C(net6),
    .A(\system_inst.loader.weight_a[2] ),
    .Y(_0170_),
    .D(net5));
 sg13g2_nand2_1 _0826_ (.Y(_0171_),
    .A(\system_inst.loader.weight_a[0] ),
    .B(net7));
 sg13g2_a22oi_1 _0827_ (.Y(_0172_),
    .B1(net5),
    .B2(\system_inst.loader.weight_a[2] ),
    .A2(net6),
    .A1(\system_inst.loader.weight_a[1] ));
 sg13g2_xor2_1 _0828_ (.B(_0169_),
    .A(_0168_),
    .X(_0173_));
 sg13g2_o21ai_1 _0829_ (.B1(_0170_),
    .Y(_0174_),
    .A1(_0171_),
    .A2(_0172_));
 sg13g2_nand2_1 _0830_ (.Y(_0175_),
    .A(\system_inst.loader.weight_a[1] ),
    .B(net7));
 sg13g2_nand2_1 _0831_ (.Y(_0176_),
    .A(\system_inst.loader.weight_a[2] ),
    .B(net7));
 sg13g2_xor2_1 _0832_ (.B(_0175_),
    .A(_0167_),
    .X(_0177_));
 sg13g2_nand2_1 _0833_ (.Y(_0178_),
    .A(_0174_),
    .B(_0177_));
 sg13g2_nand2_1 _0834_ (.Y(_0179_),
    .A(\system_inst.loader.weight_a[0] ),
    .B(net5));
 sg13g2_nor2_2 _0835_ (.A(_0168_),
    .B(_0179_),
    .Y(_0180_));
 sg13g2_xnor2_1 _0836_ (.Y(_0181_),
    .A(_0171_),
    .B(_0173_));
 sg13g2_xor2_1 _0837_ (.B(_0177_),
    .A(_0174_),
    .X(_0182_));
 sg13g2_nand3_1 _0838_ (.B(_0181_),
    .C(_0182_),
    .A(_0180_),
    .Y(_0183_));
 sg13g2_nand2_1 _0839_ (.Y(_0184_),
    .A(_0178_),
    .B(_0183_));
 sg13g2_inv_1 _0840_ (.Y(_0185_),
    .A(_0184_));
 sg13g2_nand2b_1 _0841_ (.Y(_0186_),
    .B(_0168_),
    .A_N(_0176_));
 sg13g2_xnor2_1 _0842_ (.Y(_0187_),
    .A(_0184_),
    .B(_0186_));
 sg13g2_nand2_1 _0843_ (.Y(_0188_),
    .A(_0166_),
    .B(_0187_));
 sg13g2_o21ai_1 _0844_ (.B1(_0188_),
    .Y(_0189_),
    .A1(_0105_),
    .A2(_0165_));
 sg13g2_a21oi_2 _0845_ (.B1(_0176_),
    .Y(_0190_),
    .A2(_0185_),
    .A1(_0168_));
 sg13g2_a21oi_2 _0846_ (.B1(_0154_),
    .Y(_0191_),
    .A2(_0164_),
    .A1(_0147_));
 sg13g2_xnor2_1 _0847_ (.Y(_0192_),
    .A(\system_inst.neuron.v_mem[5] ),
    .B(_0191_));
 sg13g2_nor2b_1 _0848_ (.A(_0192_),
    .B_N(_0190_),
    .Y(_0193_));
 sg13g2_xor2_1 _0849_ (.B(_0192_),
    .A(_0190_),
    .X(_0194_));
 sg13g2_nand2b_1 _0850_ (.Y(_0195_),
    .B(_0189_),
    .A_N(_0194_));
 sg13g2_xnor2_1 _0851_ (.Y(_0196_),
    .A(_0161_),
    .B(_0163_));
 sg13g2_nor2b_1 _0852_ (.A(_0196_),
    .B_N(\system_inst.neuron.v_mem[3] ),
    .Y(_0197_));
 sg13g2_xnor2_1 _0853_ (.Y(_0198_),
    .A(\system_inst.neuron.v_mem[3] ),
    .B(_0196_));
 sg13g2_a21o_1 _0854_ (.A2(_0181_),
    .A1(_0180_),
    .B1(_0182_),
    .X(_0199_));
 sg13g2_and2_1 _0855_ (.A(_0183_),
    .B(_0199_),
    .X(_0200_));
 sg13g2_a21oi_1 _0856_ (.A1(_0198_),
    .A2(_0200_),
    .Y(_0201_),
    .B1(_0197_));
 sg13g2_xnor2_1 _0857_ (.Y(_0202_),
    .A(_0166_),
    .B(_0187_));
 sg13g2_nor2_1 _0858_ (.A(_0201_),
    .B(_0202_),
    .Y(_0203_));
 sg13g2_a21oi_1 _0859_ (.A1(_0152_),
    .A2(_0160_),
    .Y(_0204_),
    .B1(_0159_));
 sg13g2_o21ai_1 _0860_ (.B1(\system_inst.neuron.v_mem[2] ),
    .Y(_0205_),
    .A1(_0161_),
    .A2(_0204_));
 sg13g2_or3_1 _0861_ (.A(\system_inst.neuron.v_mem[2] ),
    .B(_0161_),
    .C(_0204_),
    .X(_0206_));
 sg13g2_xor2_1 _0862_ (.B(_0181_),
    .A(_0180_),
    .X(_0207_));
 sg13g2_nand3_1 _0863_ (.B(_0206_),
    .C(_0207_),
    .A(_0205_),
    .Y(_0208_));
 sg13g2_nand2_1 _0864_ (.Y(_0209_),
    .A(_0205_),
    .B(_0208_));
 sg13g2_xnor2_1 _0865_ (.Y(_0210_),
    .A(_0198_),
    .B(_0200_));
 sg13g2_nor2b_1 _0866_ (.A(_0210_),
    .B_N(_0209_),
    .Y(_0211_));
 sg13g2_a22oi_1 _0867_ (.Y(_0212_),
    .B1(net10),
    .B2(net135),
    .A2(net8),
    .A1(\system_inst.loader.weight_b[0] ));
 sg13g2_nor2_1 _0868_ (.A(_0159_),
    .B(_0212_),
    .Y(_0213_));
 sg13g2_a22oi_1 _0869_ (.Y(_0214_),
    .B1(net5),
    .B2(\system_inst.loader.weight_a[1] ),
    .A2(net6),
    .A1(\system_inst.loader.weight_a[0] ));
 sg13g2_nor2_1 _0870_ (.A(_0180_),
    .B(_0214_),
    .Y(_0215_));
 sg13g2_xnor2_1 _0871_ (.Y(_0216_),
    .A(\system_inst.neuron.v_mem[1] ),
    .B(_0213_));
 sg13g2_nand2_1 _0872_ (.Y(_0217_),
    .A(_0215_),
    .B(_0216_));
 sg13g2_o21ai_1 _0873_ (.B1(_0217_),
    .Y(_0218_),
    .A1(_0106_),
    .A2(_0213_));
 sg13g2_a21o_1 _0874_ (.A2(_0206_),
    .A1(_0205_),
    .B1(_0207_),
    .X(_0219_));
 sg13g2_and3_1 _0875_ (.X(_0220_),
    .A(_0208_),
    .B(_0218_),
    .C(_0219_));
 sg13g2_nand3_1 _0876_ (.B(_0218_),
    .C(_0219_),
    .A(_0208_),
    .Y(_0221_));
 sg13g2_nor2b_1 _0877_ (.A(_0158_),
    .B_N(_0179_),
    .Y(_0222_));
 sg13g2_xnor2_1 _0878_ (.Y(_0223_),
    .A(_0215_),
    .B(_0216_));
 sg13g2_nor2_1 _0879_ (.A(_0222_),
    .B(_0223_),
    .Y(_0224_));
 sg13g2_xor2_1 _0880_ (.B(_0179_),
    .A(_0158_),
    .X(_0225_));
 sg13g2_nand2_1 _0881_ (.Y(_0226_),
    .A(\system_inst.neuron.v_mem[0] ),
    .B(_0225_));
 sg13g2_inv_1 _0882_ (.Y(_0227_),
    .A(_0226_));
 sg13g2_xor2_1 _0883_ (.B(_0223_),
    .A(_0222_),
    .X(_0228_));
 sg13g2_a21oi_1 _0884_ (.A1(_0227_),
    .A2(_0228_),
    .Y(_0229_),
    .B1(_0224_));
 sg13g2_a21oi_1 _0885_ (.A1(_0208_),
    .A2(_0219_),
    .Y(_0230_),
    .B1(_0218_));
 sg13g2_or3_1 _0886_ (.A(_0220_),
    .B(_0229_),
    .C(_0230_),
    .X(_0231_));
 sg13g2_o21ai_1 _0887_ (.B1(_0221_),
    .Y(_0232_),
    .A1(_0229_),
    .A2(_0230_));
 sg13g2_xnor2_1 _0888_ (.Y(_0233_),
    .A(_0209_),
    .B(_0210_));
 sg13g2_a21o_1 _0889_ (.A2(_0233_),
    .A1(_0232_),
    .B1(_0211_),
    .X(_0234_));
 sg13g2_xor2_1 _0890_ (.B(_0202_),
    .A(_0201_),
    .X(_0235_));
 sg13g2_a21oi_1 _0891_ (.A1(_0234_),
    .A2(_0235_),
    .Y(_0236_),
    .B1(_0203_));
 sg13g2_xor2_1 _0892_ (.B(_0194_),
    .A(_0189_),
    .X(_0237_));
 sg13g2_o21ai_1 _0893_ (.B1(_0195_),
    .Y(_0238_),
    .A1(_0236_),
    .A2(_0237_));
 sg13g2_a21o_1 _0894_ (.A2(_0191_),
    .A1(\system_inst.neuron.v_mem[5] ),
    .B1(_0193_),
    .X(_0239_));
 sg13g2_xnor2_1 _0895_ (.Y(_0240_),
    .A(\system_inst.neuron.v_mem[6] ),
    .B(_0191_));
 sg13g2_nor2b_1 _0896_ (.A(_0240_),
    .B_N(_0190_),
    .Y(_0241_));
 sg13g2_xnor2_1 _0897_ (.Y(_0242_),
    .A(_0190_),
    .B(_0240_));
 sg13g2_and2_1 _0898_ (.A(_0239_),
    .B(_0242_),
    .X(_0243_));
 sg13g2_or2_1 _0899_ (.X(_0244_),
    .B(_0242_),
    .A(_0239_));
 sg13g2_xor2_1 _0900_ (.B(_0242_),
    .A(_0239_),
    .X(_0245_));
 sg13g2_xnor2_1 _0901_ (.Y(_0246_),
    .A(_0238_),
    .B(_0245_));
 sg13g2_or2_1 _0902_ (.X(_0247_),
    .B(_0246_),
    .A(\system_inst.leak_rate[6] ));
 sg13g2_and2_1 _0903_ (.A(\system_inst.leak_rate[6] ),
    .B(_0246_),
    .X(_0248_));
 sg13g2_xor2_1 _0904_ (.B(_0246_),
    .A(\system_inst.leak_rate[6] ),
    .X(_0249_));
 sg13g2_xor2_1 _0905_ (.B(_0237_),
    .A(_0236_),
    .X(_0250_));
 sg13g2_nor2b_1 _0906_ (.A(\system_inst.leak_rate[5] ),
    .B_N(_0250_),
    .Y(_0251_));
 sg13g2_xnor2_1 _0907_ (.Y(_0252_),
    .A(_0234_),
    .B(_0235_));
 sg13g2_or2_1 _0908_ (.X(_0253_),
    .B(_0252_),
    .A(\system_inst.leak_rate[4] ));
 sg13g2_and2_1 _0909_ (.A(\system_inst.leak_rate[4] ),
    .B(_0252_),
    .X(_0254_));
 sg13g2_xor2_1 _0910_ (.B(_0252_),
    .A(\system_inst.leak_rate[4] ),
    .X(_0255_));
 sg13g2_xnor2_1 _0911_ (.Y(_0256_),
    .A(_0232_),
    .B(_0233_));
 sg13g2_nor2_1 _0912_ (.A(\system_inst.leak_rate[3] ),
    .B(_0256_),
    .Y(_0257_));
 sg13g2_o21ai_1 _0913_ (.B1(_0229_),
    .Y(_0258_),
    .A1(_0220_),
    .A2(_0230_));
 sg13g2_and2_1 _0914_ (.A(_0231_),
    .B(_0258_),
    .X(_0259_));
 sg13g2_and3_1 _0915_ (.X(_0260_),
    .A(_0099_),
    .B(_0231_),
    .C(_0258_));
 sg13g2_xnor2_1 _0916_ (.Y(_0261_),
    .A(_0226_),
    .B(_0228_));
 sg13g2_and2_1 _0917_ (.A(_0100_),
    .B(_0261_),
    .X(_0262_));
 sg13g2_xor2_1 _0918_ (.B(_0225_),
    .A(\system_inst.neuron.v_mem[0] ),
    .X(_0263_));
 sg13g2_nand2b_1 _0919_ (.Y(_0264_),
    .B(\system_inst.leak_rate[0] ),
    .A_N(_0263_));
 sg13g2_xnor2_1 _0920_ (.Y(_0265_),
    .A(\system_inst.leak_rate[1] ),
    .B(_0261_));
 sg13g2_a21o_1 _0921_ (.A2(_0265_),
    .A1(_0264_),
    .B1(_0262_),
    .X(_0266_));
 sg13g2_a21o_1 _0922_ (.A2(_0258_),
    .A1(_0231_),
    .B1(_0099_),
    .X(_0267_));
 sg13g2_nor2b_1 _0923_ (.A(_0260_),
    .B_N(_0267_),
    .Y(_0268_));
 sg13g2_a21o_1 _0924_ (.A2(_0267_),
    .A1(_0266_),
    .B1(_0260_),
    .X(_0269_));
 sg13g2_xor2_1 _0925_ (.B(_0256_),
    .A(\system_inst.leak_rate[3] ),
    .X(_0270_));
 sg13g2_a21oi_1 _0926_ (.A1(_0269_),
    .A2(_0270_),
    .Y(_0271_),
    .B1(_0257_));
 sg13g2_o21ai_1 _0927_ (.B1(_0253_),
    .Y(_0272_),
    .A1(_0254_),
    .A2(_0271_));
 sg13g2_xnor2_1 _0928_ (.Y(_0273_),
    .A(\system_inst.leak_rate[5] ),
    .B(_0250_));
 sg13g2_a21oi_1 _0929_ (.A1(_0272_),
    .A2(_0273_),
    .Y(_0274_),
    .B1(_0251_));
 sg13g2_o21ai_1 _0930_ (.B1(_0247_),
    .Y(_0275_),
    .A1(_0248_),
    .A2(_0274_));
 sg13g2_a21o_1 _0931_ (.A2(_0244_),
    .A1(_0238_),
    .B1(_0243_),
    .X(_0276_));
 sg13g2_a21o_1 _0932_ (.A2(_0191_),
    .A1(\system_inst.neuron.v_mem[6] ),
    .B1(_0241_),
    .X(_0277_));
 sg13g2_inv_1 _0933_ (.Y(_0278_),
    .A(_0277_));
 sg13g2_nor2_1 _0934_ (.A(_0190_),
    .B(_0191_),
    .Y(_0279_));
 sg13g2_nand2_1 _0935_ (.Y(_0280_),
    .A(_0190_),
    .B(_0191_));
 sg13g2_nor2b_1 _0936_ (.A(_0279_),
    .B_N(_0280_),
    .Y(_0281_));
 sg13g2_xnor2_1 _0937_ (.Y(_0282_),
    .A(\system_inst.neuron.v_mem[7] ),
    .B(_0281_));
 sg13g2_xnor2_1 _0938_ (.Y(_0283_),
    .A(_0278_),
    .B(_0282_));
 sg13g2_nand2b_1 _0939_ (.Y(_0284_),
    .B(_0276_),
    .A_N(_0283_));
 sg13g2_xor2_1 _0940_ (.B(_0283_),
    .A(_0276_),
    .X(_0285_));
 sg13g2_xor2_1 _0941_ (.B(_0285_),
    .A(\system_inst.leak_rate[7] ),
    .X(_0286_));
 sg13g2_nand2b_1 _0942_ (.Y(_0287_),
    .B(\system_inst.leak_cycles[3] ),
    .A_N(\system_inst.neuron.leak_counter[3] ));
 sg13g2_nor2_1 _0943_ (.A(\system_inst.leak_cycles[1] ),
    .B(_0102_),
    .Y(_0288_));
 sg13g2_nor3_1 _0944_ (.A(_0093_),
    .B(\system_inst.neuron.leak_counter[0] ),
    .C(_0288_),
    .Y(_0289_));
 sg13g2_a221oi_1 _0945_ (.B2(\system_inst.leak_cycles[1] ),
    .C1(_0289_),
    .B1(_0102_),
    .A1(\system_inst.leak_cycles[2] ),
    .Y(_0290_),
    .A2(_0101_));
 sg13g2_nand2b_1 _0946_ (.Y(_0291_),
    .B(\system_inst.neuron.leak_counter[3] ),
    .A_N(\system_inst.leak_cycles[3] ));
 sg13g2_o21ai_1 _0947_ (.B1(_0291_),
    .Y(_0292_),
    .A1(\system_inst.leak_cycles[2] ),
    .A2(_0101_));
 sg13g2_o21ai_1 _0948_ (.B1(_0287_),
    .Y(_0293_),
    .A1(_0290_),
    .A2(_0292_));
 sg13g2_inv_2 _0949_ (.Y(_0294_),
    .A(net124));
 sg13g2_o21ai_1 _0950_ (.B1(_0294_),
    .Y(_0295_),
    .A1(\system_inst.leak_rate[7] ),
    .A2(_0285_));
 sg13g2_a21oi_2 _0951_ (.B1(_0295_),
    .Y(_0296_),
    .A2(_0286_),
    .A1(_0275_));
 sg13g2_o21ai_1 _0952_ (.B1(_0284_),
    .Y(_0297_),
    .A1(_0278_),
    .A2(_0282_));
 sg13g2_a21oi_1 _0953_ (.A1(\system_inst.neuron.v_mem[7] ),
    .A2(_0280_),
    .Y(_0298_),
    .B1(_0279_));
 sg13g2_xor2_1 _0954_ (.B(_0298_),
    .A(net136),
    .X(_0299_));
 sg13g2_xnor2_1 _0955_ (.Y(_0300_),
    .A(_0297_),
    .B(_0299_));
 sg13g2_xnor2_1 _0956_ (.Y(_0301_),
    .A(_0296_),
    .B(_0300_));
 sg13g2_xor2_1 _0957_ (.B(_0300_),
    .A(_0296_),
    .X(_0302_));
 sg13g2_xor2_1 _0958_ (.B(_0286_),
    .A(_0275_),
    .X(_0303_));
 sg13g2_nand2_1 _0959_ (.Y(_0304_),
    .A(_0285_),
    .B(net124));
 sg13g2_o21ai_1 _0960_ (.B1(_0304_),
    .Y(_0305_),
    .A1(net124),
    .A2(_0303_));
 sg13g2_nor3_1 _0961_ (.A(_0108_),
    .B(net118),
    .C(_0305_),
    .Y(_0306_));
 sg13g2_o21ai_1 _0962_ (.B1(_0108_),
    .Y(_0307_),
    .A1(net117),
    .A2(_0305_));
 sg13g2_nand2b_1 _0963_ (.Y(_0308_),
    .B(_0307_),
    .A_N(_0306_));
 sg13g2_nor2_1 _0964_ (.A(_0246_),
    .B(_0294_),
    .Y(_0309_));
 sg13g2_xnor2_1 _0965_ (.Y(_0310_),
    .A(_0249_),
    .B(_0274_));
 sg13g2_a21oi_1 _0966_ (.A1(_0294_),
    .A2(_0310_),
    .Y(_0311_),
    .B1(_0309_));
 sg13g2_nor2_1 _0967_ (.A(net117),
    .B(_0311_),
    .Y(_0312_));
 sg13g2_xnor2_1 _0968_ (.Y(_0313_),
    .A(_0109_),
    .B(_0312_));
 sg13g2_nor2_1 _0969_ (.A(_0308_),
    .B(_0313_),
    .Y(_0314_));
 sg13g2_xnor2_1 _0970_ (.Y(_0315_),
    .A(_0272_),
    .B(_0273_));
 sg13g2_nor2_1 _0971_ (.A(_0250_),
    .B(_0294_),
    .Y(_0316_));
 sg13g2_a21oi_1 _0972_ (.A1(_0294_),
    .A2(_0315_),
    .Y(_0317_),
    .B1(_0316_));
 sg13g2_nand2_1 _0973_ (.Y(_0318_),
    .A(_0302_),
    .B(_0317_));
 sg13g2_xor2_1 _0974_ (.B(_0318_),
    .A(_0008_),
    .X(_0319_));
 sg13g2_xnor2_1 _0975_ (.Y(_0320_),
    .A(_0255_),
    .B(_0271_));
 sg13g2_nor2_1 _0976_ (.A(net125),
    .B(_0320_),
    .Y(_0321_));
 sg13g2_a21oi_1 _0977_ (.A1(_0252_),
    .A2(net124),
    .Y(_0322_),
    .B1(_0321_));
 sg13g2_nand2_2 _0978_ (.Y(_0323_),
    .A(_0302_),
    .B(_0322_));
 sg13g2_nand2_1 _0979_ (.Y(_0324_),
    .A(\system_inst.neuron.threshold[4] ),
    .B(_0323_));
 sg13g2_xnor2_1 _0980_ (.Y(_0325_),
    .A(\system_inst.neuron.threshold[4] ),
    .B(_0323_));
 sg13g2_or4_1 _0981_ (.A(_0308_),
    .B(_0313_),
    .C(_0319_),
    .D(_0325_),
    .X(_0326_));
 sg13g2_or2_1 _0982_ (.X(_0327_),
    .B(_0268_),
    .A(_0266_));
 sg13g2_a21oi_1 _0983_ (.A1(_0266_),
    .A2(_0268_),
    .Y(_0328_),
    .B1(net124));
 sg13g2_a22oi_1 _0984_ (.Y(_0329_),
    .B1(_0327_),
    .B2(_0328_),
    .A2(net124),
    .A1(_0259_));
 sg13g2_inv_1 _0985_ (.Y(_0330_),
    .A(_0329_));
 sg13g2_nor3_1 _0986_ (.A(\system_inst.neuron.threshold[2] ),
    .B(net117),
    .C(_0329_),
    .Y(_0331_));
 sg13g2_a21oi_1 _0987_ (.A1(_0302_),
    .A2(_0330_),
    .Y(_0332_),
    .B1(_0113_));
 sg13g2_xor2_1 _0988_ (.B(_0270_),
    .A(_0269_),
    .X(_0333_));
 sg13g2_nand2_1 _0989_ (.Y(_0334_),
    .A(_0256_),
    .B(net124));
 sg13g2_o21ai_1 _0990_ (.B1(_0334_),
    .Y(_0335_),
    .A1(net124),
    .A2(_0333_));
 sg13g2_inv_1 _0991_ (.Y(_0336_),
    .A(_0335_));
 sg13g2_a21oi_1 _0992_ (.A1(_0302_),
    .A2(_0336_),
    .Y(_0337_),
    .B1(_0009_));
 sg13g2_and3_1 _0993_ (.X(_0338_),
    .A(_0009_),
    .B(_0302_),
    .C(_0336_));
 sg13g2_nor4_1 _0994_ (.A(_0331_),
    .B(_0332_),
    .C(_0337_),
    .D(_0338_),
    .Y(_0339_));
 sg13g2_nand2_1 _0995_ (.Y(_0340_),
    .A(\system_inst.leak_rate[0] ),
    .B(_0294_));
 sg13g2_xor2_1 _0996_ (.B(_0340_),
    .A(_0263_),
    .X(_0341_));
 sg13g2_nor2_1 _0997_ (.A(net117),
    .B(_0341_),
    .Y(_0342_));
 sg13g2_xnor2_1 _0998_ (.Y(_0343_),
    .A(_0264_),
    .B(_0265_));
 sg13g2_nand2_1 _0999_ (.Y(_0344_),
    .A(_0294_),
    .B(_0343_));
 sg13g2_o21ai_1 _1000_ (.B1(_0344_),
    .Y(_0345_),
    .A1(_0261_),
    .A2(_0294_));
 sg13g2_inv_1 _1001_ (.Y(_0346_),
    .A(_0345_));
 sg13g2_nand3_1 _1002_ (.B(_0302_),
    .C(_0346_),
    .A(\system_inst.neuron.threshold[1] ),
    .Y(_0347_));
 sg13g2_o21ai_1 _1003_ (.B1(_0114_),
    .Y(_0348_),
    .A1(net117),
    .A2(_0345_));
 sg13g2_a22oi_1 _1004_ (.Y(_0349_),
    .B1(_0347_),
    .B2(_0348_),
    .A2(_0342_),
    .A1(_0115_));
 sg13g2_a21oi_1 _1005_ (.A1(_0302_),
    .A2(_0346_),
    .Y(_0350_),
    .B1(_0011_));
 sg13g2_o21ai_1 _1006_ (.B1(_0339_),
    .Y(_0351_),
    .A1(_0349_),
    .A2(_0350_));
 sg13g2_a21oi_1 _1007_ (.A1(_0302_),
    .A2(_0330_),
    .Y(_0352_),
    .B1(_0010_));
 sg13g2_nor2_1 _1008_ (.A(_0337_),
    .B(_0352_),
    .Y(_0353_));
 sg13g2_or2_1 _1009_ (.X(_0354_),
    .B(_0353_),
    .A(_0338_));
 sg13g2_a21o_1 _1010_ (.A2(_0354_),
    .A1(_0351_),
    .B1(_0326_),
    .X(_0355_));
 sg13g2_nand2_1 _1011_ (.Y(_0356_),
    .A(\system_inst.neuron.threshold[5] ),
    .B(_0318_));
 sg13g2_o21ai_1 _1012_ (.B1(_0356_),
    .Y(_0357_),
    .A1(_0319_),
    .A2(_0324_));
 sg13g2_o21ai_1 _1013_ (.B1(_0307_),
    .Y(_0358_),
    .A1(_0007_),
    .A2(_0312_));
 sg13g2_nor2b_1 _1014_ (.A(_0306_),
    .B_N(_0358_),
    .Y(_0359_));
 sg13g2_a21oi_1 _1015_ (.A1(_0314_),
    .A2(_0357_),
    .Y(_0360_),
    .B1(_0359_));
 sg13g2_o21ai_1 _1016_ (.B1(\system_inst.neuron.threshold[0] ),
    .Y(_0361_),
    .A1(net117),
    .A2(_0341_));
 sg13g2_nand3_1 _1017_ (.B(_0349_),
    .C(_0361_),
    .A(_0339_),
    .Y(_0362_));
 sg13g2_nor2_1 _1018_ (.A(_0326_),
    .B(_0362_),
    .Y(_0363_));
 sg13g2_a21oi_2 _1019_ (.B1(_0363_),
    .Y(_0364_),
    .A2(_0360_),
    .A1(_0355_));
 sg13g2_a21o_1 _1020_ (.A2(_0360_),
    .A1(_0355_),
    .B1(_0363_),
    .X(_0365_));
 sg13g2_nor3_1 _1021_ (.A(net132),
    .B(net118),
    .C(_0341_),
    .Y(_0366_));
 sg13g2_a22oi_1 _1022_ (.Y(_0367_),
    .B1(net116),
    .B2(_0366_),
    .A2(net133),
    .A1(net170));
 sg13g2_nor2_1 _1023_ (.A(net140),
    .B(_0367_),
    .Y(_0022_));
 sg13g2_nor3_1 _1024_ (.A(net133),
    .B(net118),
    .C(_0345_),
    .Y(_0368_));
 sg13g2_a22oi_1 _1025_ (.Y(_0369_),
    .B1(_0364_),
    .B2(_0368_),
    .A2(net133),
    .A1(net164));
 sg13g2_nor2_1 _1026_ (.A(net140),
    .B(_0369_),
    .Y(_0023_));
 sg13g2_nor3_1 _1027_ (.A(net133),
    .B(net118),
    .C(_0329_),
    .Y(_0370_));
 sg13g2_a22oi_1 _1028_ (.Y(_0371_),
    .B1(net115),
    .B2(_0370_),
    .A2(net132),
    .A1(net160));
 sg13g2_nor2_1 _1029_ (.A(net138),
    .B(_0371_),
    .Y(_0024_));
 sg13g2_nor3_1 _1030_ (.A(net132),
    .B(net118),
    .C(_0335_),
    .Y(_0372_));
 sg13g2_a22oi_1 _1031_ (.Y(_0373_),
    .B1(net115),
    .B2(_0372_),
    .A2(net132),
    .A1(net191));
 sg13g2_nor2_1 _1032_ (.A(net138),
    .B(_0373_),
    .Y(_0025_));
 sg13g2_nor2_1 _1033_ (.A(net131),
    .B(_0323_),
    .Y(_0374_));
 sg13g2_a22oi_1 _1034_ (.Y(_0375_),
    .B1(net115),
    .B2(_0374_),
    .A2(net131),
    .A1(net180));
 sg13g2_nor2_1 _1035_ (.A(net138),
    .B(_0375_),
    .Y(_0026_));
 sg13g2_nor2_1 _1036_ (.A(net131),
    .B(_0318_),
    .Y(_0376_));
 sg13g2_a22oi_1 _1037_ (.Y(_0377_),
    .B1(net115),
    .B2(_0376_),
    .A2(net131),
    .A1(net177));
 sg13g2_nor2_1 _1038_ (.A(net138),
    .B(_0377_),
    .Y(_0027_));
 sg13g2_nor3_1 _1039_ (.A(net131),
    .B(net117),
    .C(_0311_),
    .Y(_0378_));
 sg13g2_a22oi_1 _1040_ (.Y(_0379_),
    .B1(net115),
    .B2(_0378_),
    .A2(net132),
    .A1(net175));
 sg13g2_nor2_1 _1041_ (.A(net138),
    .B(_0379_),
    .Y(_0028_));
 sg13g2_nor3_1 _1042_ (.A(net131),
    .B(net117),
    .C(_0305_),
    .Y(_0380_));
 sg13g2_a22oi_1 _1043_ (.Y(_0381_),
    .B1(net115),
    .B2(_0380_),
    .A2(net132),
    .A1(net153));
 sg13g2_nor2_1 _1044_ (.A(net138),
    .B(_0381_),
    .Y(_0029_));
 sg13g2_and3_1 _1045_ (.X(_0030_),
    .A(net136),
    .B(net143),
    .C(net132));
 sg13g2_nand2_1 _1046_ (.Y(_0382_),
    .A(net143),
    .B(_0365_));
 sg13g2_nor2_1 _1047_ (.A(net131),
    .B(_0382_),
    .Y(_0031_));
 sg13g2_nor2_1 _1048_ (.A(_0140_),
    .B(_0142_),
    .Y(_0383_));
 sg13g2_inv_1 _1049_ (.Y(_0384_),
    .A(_0383_));
 sg13g2_o21ai_1 _1050_ (.B1(_0384_),
    .Y(_0385_),
    .A1(_0144_),
    .A2(_0364_));
 sg13g2_o21ai_1 _1051_ (.B1(_0385_),
    .Y(_0386_),
    .A1(net207),
    .A2(_0142_));
 sg13g2_o21ai_1 _1052_ (.B1(net148),
    .Y(_0387_),
    .A1(net207),
    .A2(_0385_));
 sg13g2_nor2b_1 _1053_ (.A(_0387_),
    .B_N(_0386_),
    .Y(_0032_));
 sg13g2_and2_1 _1054_ (.A(\system_inst.neuron.refr_cnt[1] ),
    .B(\system_inst.neuron.refr_cnt[0] ),
    .X(_0388_));
 sg13g2_o21ai_1 _1055_ (.B1(_0383_),
    .Y(_0389_),
    .A1(_0141_),
    .A2(_0388_));
 sg13g2_o21ai_1 _1056_ (.B1(_0389_),
    .Y(_0390_),
    .A1(_0104_),
    .A2(_0385_));
 sg13g2_and2_1 _1057_ (.A(net147),
    .B(_0390_),
    .X(_0033_));
 sg13g2_nand3_1 _1058_ (.B(_0141_),
    .C(_0385_),
    .A(_0103_),
    .Y(_0391_));
 sg13g2_a21o_1 _1059_ (.A2(_0385_),
    .A1(_0141_),
    .B1(_0103_),
    .X(_0392_));
 sg13g2_a21oi_1 _1060_ (.A1(net206),
    .A2(_0392_),
    .Y(_0034_),
    .B1(net140));
 sg13g2_and3_1 _1061_ (.X(_0035_),
    .A(net95),
    .B(net147),
    .C(_0391_));
 sg13g2_nor2_1 _1062_ (.A(\system_inst.neuron.leak_counter[0] ),
    .B(_0143_),
    .Y(_0393_));
 sg13g2_a221oi_1 _1063_ (.B2(_0393_),
    .C1(_0140_),
    .B1(net125),
    .A1(net109),
    .Y(_0394_),
    .A2(_0143_));
 sg13g2_o21ai_1 _1064_ (.B1(net148),
    .Y(_0395_),
    .A1(\system_inst.neuron.leak_counter[0] ),
    .A2(_0139_));
 sg13g2_nor2_1 _1065_ (.A(net110),
    .B(_0395_),
    .Y(_0036_));
 sg13g2_o21ai_1 _1066_ (.B1(net147),
    .Y(_0396_),
    .A1(_0145_),
    .A2(net125));
 sg13g2_inv_2 _1067_ (.Y(_0397_),
    .A(_0396_));
 sg13g2_and3_1 _1068_ (.X(_0398_),
    .A(net99),
    .B(\system_inst.neuron.leak_counter[0] ),
    .C(_0139_));
 sg13g2_a21oi_1 _1069_ (.A1(\system_inst.neuron.leak_counter[0] ),
    .A2(_0139_),
    .Y(_0399_),
    .B1(net99));
 sg13g2_nor3_1 _1070_ (.A(_0396_),
    .B(_0398_),
    .C(net100),
    .Y(_0037_));
 sg13g2_nand2_1 _1071_ (.Y(_0400_),
    .A(net187),
    .B(_0398_));
 sg13g2_o21ai_1 _1072_ (.B1(_0397_),
    .Y(_0401_),
    .A1(net187),
    .A2(_0398_));
 sg13g2_nor2b_1 _1073_ (.A(net188),
    .B_N(_0400_),
    .Y(_0038_));
 sg13g2_xor2_1 _1074_ (.B(_0400_),
    .A(net185),
    .X(_0402_));
 sg13g2_nor2_1 _1075_ (.A(_0396_),
    .B(net186),
    .Y(_0039_));
 sg13g2_o21ai_1 _1076_ (.B1(_0397_),
    .Y(_0403_),
    .A1(net131),
    .A2(net115));
 sg13g2_nand2_1 _1077_ (.Y(_0404_),
    .A(net196),
    .B(net137));
 sg13g2_o21ai_1 _1078_ (.B1(_0404_),
    .Y(_0405_),
    .A1(_0113_),
    .A2(net114));
 sg13g2_nand2_1 _1079_ (.Y(_0406_),
    .A(\system_inst.neuron.threshold[3] ),
    .B(\system_inst.neuron.threshold[2] ));
 sg13g2_nand4_1 _1080_ (.B(\system_inst.neuron.threshold[4] ),
    .C(\system_inst.neuron.threshold[3] ),
    .A(\system_inst.neuron.threshold[5] ),
    .Y(_0407_),
    .D(\system_inst.neuron.threshold[2] ));
 sg13g2_nor2_1 _1081_ (.A(_0007_),
    .B(_0407_),
    .Y(_0408_));
 sg13g2_xnor2_1 _1082_ (.Y(_0409_),
    .A(_0006_),
    .B(_0408_));
 sg13g2_nor2b_1 _1083_ (.A(\system_inst.loader.threshold_min[6] ),
    .B_N(_0409_),
    .Y(_0410_));
 sg13g2_xor2_1 _1084_ (.B(_0407_),
    .A(_0007_),
    .X(_0411_));
 sg13g2_nor2_1 _1085_ (.A(_0016_),
    .B(_0406_),
    .Y(_0412_));
 sg13g2_xnor2_1 _1086_ (.Y(_0413_),
    .A(_0008_),
    .B(_0412_));
 sg13g2_nor2_1 _1087_ (.A(_0017_),
    .B(_0413_),
    .Y(_0414_));
 sg13g2_xnor2_1 _1088_ (.Y(_0415_),
    .A(_0018_),
    .B(_0411_));
 sg13g2_nor2_1 _1089_ (.A(_0414_),
    .B(_0415_),
    .Y(_0416_));
 sg13g2_xor2_1 _1090_ (.B(_0406_),
    .A(_0016_),
    .X(_0417_));
 sg13g2_xor2_1 _1091_ (.B(_0417_),
    .A(_0015_),
    .X(_0418_));
 sg13g2_xor2_1 _1092_ (.B(\system_inst.neuron.threshold[2] ),
    .A(\system_inst.neuron.threshold[3] ),
    .X(_0419_));
 sg13g2_nand2_1 _1093_ (.Y(_0420_),
    .A(_0014_),
    .B(_0419_));
 sg13g2_or2_1 _1094_ (.X(_0421_),
    .B(_0419_),
    .A(_0014_));
 sg13g2_a22oi_1 _1095_ (.Y(_0422_),
    .B1(_0114_),
    .B2(\system_inst.loader.threshold_min[0] ),
    .A2(\system_inst.neuron.threshold[2] ),
    .A1(\system_inst.loader.threshold_min[1] ));
 sg13g2_nor2_1 _1096_ (.A(\system_inst.loader.threshold_min[1] ),
    .B(\system_inst.neuron.threshold[2] ),
    .Y(_0423_));
 sg13g2_o21ai_1 _1097_ (.B1(_0421_),
    .Y(_0424_),
    .A1(_0422_),
    .A2(_0423_));
 sg13g2_nand2_1 _1098_ (.Y(_0425_),
    .A(_0420_),
    .B(_0424_));
 sg13g2_nand2_1 _1099_ (.Y(_0426_),
    .A(_0418_),
    .B(_0425_));
 sg13g2_nand2b_1 _1100_ (.Y(_0427_),
    .B(_0417_),
    .A_N(\system_inst.loader.threshold_min[3] ));
 sg13g2_nand2_1 _1101_ (.Y(_0428_),
    .A(_0017_),
    .B(_0413_));
 sg13g2_nand3_1 _1102_ (.B(_0427_),
    .C(_0428_),
    .A(_0426_),
    .Y(_0429_));
 sg13g2_a22oi_1 _1103_ (.Y(_0430_),
    .B1(_0416_),
    .B2(_0429_),
    .A2(_0411_),
    .A1(_0095_));
 sg13g2_xor2_1 _1104_ (.B(_0409_),
    .A(_0019_),
    .X(_0431_));
 sg13g2_nor2b_1 _1105_ (.A(_0430_),
    .B_N(_0431_),
    .Y(_0432_));
 sg13g2_a21oi_1 _1106_ (.A1(_0098_),
    .A2(\system_inst.neuron.threshold[1] ),
    .Y(_0433_),
    .B1(_0423_));
 sg13g2_and3_1 _1107_ (.X(_0434_),
    .A(_0115_),
    .B(_0422_),
    .C(_0433_));
 sg13g2_and4_1 _1108_ (.A(_0420_),
    .B(_0421_),
    .C(_0428_),
    .D(_0434_),
    .X(_0435_));
 sg13g2_nand4_1 _1109_ (.B(_0418_),
    .C(_0431_),
    .A(_0416_),
    .Y(_0436_),
    .D(_0435_));
 sg13g2_o21ai_1 _1110_ (.B1(_0436_),
    .Y(_0437_),
    .A1(_0410_),
    .A2(_0432_));
 sg13g2_inv_1 _1111_ (.Y(_0438_),
    .A(net121));
 sg13g2_nand2_1 _1112_ (.Y(_0439_),
    .A(_0010_),
    .B(_0437_));
 sg13g2_o21ai_1 _1113_ (.B1(_0439_),
    .Y(_0440_),
    .A1(_0097_),
    .A2(_0437_));
 sg13g2_nand2_1 _1114_ (.Y(_0441_),
    .A(\system_inst.loader.threshold_min[1] ),
    .B(\system_inst.loader.threshold_min[0] ));
 sg13g2_nand4_1 _1115_ (.B(\system_inst.loader.threshold_min[2] ),
    .C(\system_inst.loader.threshold_min[1] ),
    .A(\system_inst.loader.threshold_min[3] ),
    .Y(_0442_),
    .D(\system_inst.loader.threshold_min[0] ));
 sg13g2_or3_1 _1116_ (.A(_0095_),
    .B(_0096_),
    .C(_0442_),
    .X(_0443_));
 sg13g2_nor2_1 _1117_ (.A(_0019_),
    .B(_0443_),
    .Y(_0444_));
 sg13g2_xnor2_1 _1118_ (.Y(_0445_),
    .A(\system_inst.loader.threshold_min[7] ),
    .B(_0444_));
 sg13g2_nand2_1 _1119_ (.Y(_0446_),
    .A(\system_inst.neuron.threshold[7] ),
    .B(_0445_));
 sg13g2_xor2_1 _1120_ (.B(_0443_),
    .A(_0019_),
    .X(_0447_));
 sg13g2_inv_1 _1121_ (.Y(_0448_),
    .A(_0447_));
 sg13g2_nor2_1 _1122_ (.A(_0017_),
    .B(_0442_),
    .Y(_0449_));
 sg13g2_xnor2_1 _1123_ (.Y(_0450_),
    .A(_0018_),
    .B(_0449_));
 sg13g2_nand2b_1 _1124_ (.Y(_0451_),
    .B(\system_inst.neuron.threshold[5] ),
    .A_N(_0450_));
 sg13g2_xor2_1 _1125_ (.B(_0442_),
    .A(_0017_),
    .X(_0452_));
 sg13g2_xnor2_1 _1126_ (.Y(_0453_),
    .A(_0008_),
    .B(_0450_));
 sg13g2_a21o_1 _1127_ (.A2(_0452_),
    .A1(_0016_),
    .B1(_0453_),
    .X(_0454_));
 sg13g2_nor2_1 _1128_ (.A(_0014_),
    .B(_0441_),
    .Y(_0455_));
 sg13g2_xor2_1 _1129_ (.B(_0455_),
    .A(_0015_),
    .X(_0456_));
 sg13g2_nand2b_1 _1130_ (.Y(_0457_),
    .B(_0112_),
    .A_N(_0456_));
 sg13g2_xor2_1 _1131_ (.B(_0441_),
    .A(_0014_),
    .X(_0458_));
 sg13g2_xnor2_1 _1132_ (.Y(_0459_),
    .A(_0010_),
    .B(_0458_));
 sg13g2_nand2_1 _1133_ (.Y(_0460_),
    .A(\system_inst.neuron.threshold[3] ),
    .B(_0456_));
 sg13g2_a21oi_1 _1134_ (.A1(\system_inst.neuron.threshold[3] ),
    .A2(_0456_),
    .Y(_0461_),
    .B1(_0459_));
 sg13g2_and2_1 _1135_ (.A(_0457_),
    .B(_0461_),
    .X(_0462_));
 sg13g2_xor2_1 _1136_ (.B(\system_inst.loader.threshold_min[0] ),
    .A(\system_inst.loader.threshold_min[1] ),
    .X(_0463_));
 sg13g2_xor2_1 _1137_ (.B(_0463_),
    .A(_0011_),
    .X(_0464_));
 sg13g2_o21ai_1 _1138_ (.B1(_0464_),
    .Y(_0465_),
    .A1(\system_inst.loader.threshold_min[0] ),
    .A2(\system_inst.neuron.threshold[0] ));
 sg13g2_o21ai_1 _1139_ (.B1(_0465_),
    .Y(_0466_),
    .A1(_0114_),
    .A2(_0463_));
 sg13g2_nor2_1 _1140_ (.A(_0113_),
    .B(_0458_),
    .Y(_0467_));
 sg13g2_or2_1 _1141_ (.X(_0468_),
    .B(_0452_),
    .A(_0016_));
 sg13g2_nand2_1 _1142_ (.Y(_0469_),
    .A(_0460_),
    .B(_0468_));
 sg13g2_a221oi_1 _1143_ (.B2(_0457_),
    .C1(_0469_),
    .B1(_0467_),
    .A1(_0462_),
    .Y(_0470_),
    .A2(_0466_));
 sg13g2_o21ai_1 _1144_ (.B1(_0451_),
    .Y(_0471_),
    .A1(_0454_),
    .A2(_0470_));
 sg13g2_xor2_1 _1145_ (.B(_0447_),
    .A(_0007_),
    .X(_0472_));
 sg13g2_a22oi_1 _1146_ (.Y(_0473_),
    .B1(_0471_),
    .B2(_0472_),
    .A2(_0448_),
    .A1(\system_inst.neuron.threshold[6] ));
 sg13g2_nand2b_1 _1147_ (.Y(_0474_),
    .B(_0107_),
    .A_N(_0445_));
 sg13g2_a21oi_1 _1148_ (.A1(\system_inst.loader.threshold_min[0] ),
    .A2(\system_inst.neuron.threshold[0] ),
    .Y(_0475_),
    .B1(_0465_));
 sg13g2_nand4_1 _1149_ (.B(_0468_),
    .C(_0472_),
    .A(_0462_),
    .Y(_0476_),
    .D(_0475_));
 sg13g2_o21ai_1 _1150_ (.B1(_0474_),
    .Y(_0477_),
    .A1(_0454_),
    .A2(_0476_));
 sg13g2_o21ai_1 _1151_ (.B1(_0446_),
    .Y(_0478_),
    .A1(_0473_),
    .A2(_0477_));
 sg13g2_nor2_1 _1152_ (.A(\system_inst.neuron.threshold[1] ),
    .B(\system_inst.neuron.threshold[0] ),
    .Y(_0479_));
 sg13g2_nor3_1 _1153_ (.A(\system_inst.neuron.threshold[2] ),
    .B(\system_inst.neuron.threshold[1] ),
    .C(\system_inst.neuron.threshold[0] ),
    .Y(_0480_));
 sg13g2_xnor2_1 _1154_ (.Y(_0481_),
    .A(_0113_),
    .B(_0479_));
 sg13g2_mux2_1 _1155_ (.A0(\system_inst.loader.threshold_min[2] ),
    .A1(_0481_),
    .S(net120),
    .X(_0482_));
 sg13g2_mux2_1 _1156_ (.A0(_0440_),
    .A1(_0482_),
    .S(net116),
    .X(_0483_));
 sg13g2_nand3_1 _1157_ (.B(net114),
    .C(_0483_),
    .A(net141),
    .Y(_0484_));
 sg13g2_nand2b_1 _1158_ (.Y(_0040_),
    .B(_0484_),
    .A_N(_0405_));
 sg13g2_mux2_1 _1159_ (.A0(\system_inst.loader.threshold_min[2] ),
    .A1(_0419_),
    .S(net121),
    .X(_0485_));
 sg13g2_and2_1 _1160_ (.A(_0112_),
    .B(_0480_),
    .X(_0486_));
 sg13g2_xnor2_1 _1161_ (.Y(_0487_),
    .A(_0112_),
    .B(_0480_));
 sg13g2_mux2_1 _1162_ (.A0(\system_inst.loader.threshold_min[3] ),
    .A1(_0487_),
    .S(net120),
    .X(_0488_));
 sg13g2_mux2_1 _1163_ (.A0(_0485_),
    .A1(_0488_),
    .S(net116),
    .X(_0489_));
 sg13g2_nand3_1 _1164_ (.B(net114),
    .C(_0489_),
    .A(net141),
    .Y(_0490_));
 sg13g2_nand2_1 _1165_ (.Y(_0491_),
    .A(net204),
    .B(net137));
 sg13g2_o21ai_1 _1166_ (.B1(_0491_),
    .Y(_0492_),
    .A1(_0112_),
    .A2(net114));
 sg13g2_nand2b_1 _1167_ (.Y(_0041_),
    .B(_0490_),
    .A_N(_0492_));
 sg13g2_mux2_1 _1168_ (.A0(\system_inst.loader.threshold_min[3] ),
    .A1(_0417_),
    .S(net121),
    .X(_0493_));
 sg13g2_and2_1 _1169_ (.A(_0111_),
    .B(_0486_),
    .X(_0494_));
 sg13g2_nor2_1 _1170_ (.A(_0111_),
    .B(_0486_),
    .Y(_0495_));
 sg13g2_o21ai_1 _1171_ (.B1(net119),
    .Y(_0496_),
    .A1(_0494_),
    .A2(_0495_));
 sg13g2_o21ai_1 _1172_ (.B1(_0496_),
    .Y(_0497_),
    .A1(_0096_),
    .A2(net119));
 sg13g2_mux2_1 _1173_ (.A0(_0493_),
    .A1(_0497_),
    .S(net116),
    .X(_0498_));
 sg13g2_nand3_1 _1174_ (.B(net113),
    .C(_0498_),
    .A(net141),
    .Y(_0499_));
 sg13g2_nand2_1 _1175_ (.Y(_0500_),
    .A(net201),
    .B(net137));
 sg13g2_o21ai_1 _1176_ (.B1(_0500_),
    .Y(_0501_),
    .A1(_0111_),
    .A2(net113));
 sg13g2_nand2b_1 _1177_ (.Y(_0042_),
    .B(_0499_),
    .A_N(_0501_));
 sg13g2_nand2_1 _1178_ (.Y(_0502_),
    .A(net157),
    .B(net137));
 sg13g2_o21ai_1 _1179_ (.B1(_0502_),
    .Y(_0503_),
    .A1(_0110_),
    .A2(net113));
 sg13g2_nand2_1 _1180_ (.Y(_0504_),
    .A(_0413_),
    .B(net121));
 sg13g2_o21ai_1 _1181_ (.B1(_0504_),
    .Y(_0505_),
    .A1(_0096_),
    .A2(net121));
 sg13g2_and2_1 _1182_ (.A(_0110_),
    .B(_0494_),
    .X(_0506_));
 sg13g2_nor2_1 _1183_ (.A(_0110_),
    .B(_0494_),
    .Y(_0507_));
 sg13g2_o21ai_1 _1184_ (.B1(net119),
    .Y(_0508_),
    .A1(_0506_),
    .A2(_0507_));
 sg13g2_o21ai_1 _1185_ (.B1(_0508_),
    .Y(_0509_),
    .A1(_0095_),
    .A2(net119));
 sg13g2_mux2_1 _1186_ (.A0(_0505_),
    .A1(_0509_),
    .S(net116),
    .X(_0510_));
 sg13g2_nand3_1 _1187_ (.B(net113),
    .C(_0510_),
    .A(net141),
    .Y(_0511_));
 sg13g2_nand2b_1 _1188_ (.Y(_0043_),
    .B(_0511_),
    .A_N(_0503_));
 sg13g2_nand2_1 _1189_ (.Y(_0512_),
    .A(_0411_),
    .B(net121));
 sg13g2_o21ai_1 _1190_ (.B1(_0512_),
    .Y(_0513_),
    .A1(_0095_),
    .A2(net121));
 sg13g2_nand2_1 _1191_ (.Y(_0514_),
    .A(_0109_),
    .B(_0506_));
 sg13g2_xnor2_1 _1192_ (.Y(_0515_),
    .A(\system_inst.neuron.threshold[6] ),
    .B(_0506_));
 sg13g2_nor2_1 _1193_ (.A(\system_inst.loader.threshold_min[6] ),
    .B(net119),
    .Y(_0516_));
 sg13g2_a21oi_1 _1194_ (.A1(net119),
    .A2(_0515_),
    .Y(_0517_),
    .B1(_0516_));
 sg13g2_mux2_1 _1195_ (.A0(_0513_),
    .A1(_0517_),
    .S(net116),
    .X(_0518_));
 sg13g2_nand3_1 _1196_ (.B(net113),
    .C(_0518_),
    .A(net141),
    .Y(_0519_));
 sg13g2_nand2_1 _1197_ (.Y(_0520_),
    .A(net217),
    .B(net137));
 sg13g2_o21ai_1 _1198_ (.B1(_0520_),
    .Y(_0521_),
    .A1(_0109_),
    .A2(net113));
 sg13g2_nand2b_1 _1199_ (.Y(_0044_),
    .B(_0519_),
    .A_N(net218));
 sg13g2_nand2_1 _1200_ (.Y(_0522_),
    .A(net172),
    .B(net137));
 sg13g2_o21ai_1 _1201_ (.B1(_0522_),
    .Y(_0523_),
    .A1(_0107_),
    .A2(net113));
 sg13g2_mux2_1 _1202_ (.A0(\system_inst.loader.threshold_min[6] ),
    .A1(_0409_),
    .S(net121),
    .X(_0524_));
 sg13g2_xnor2_1 _1203_ (.Y(_0525_),
    .A(\system_inst.neuron.threshold[7] ),
    .B(_0514_));
 sg13g2_mux2_1 _1204_ (.A0(\system_inst.loader.threshold_min[7] ),
    .A1(_0525_),
    .S(net119),
    .X(_0526_));
 sg13g2_mux2_1 _1205_ (.A0(_0524_),
    .A1(_0526_),
    .S(net116),
    .X(_0527_));
 sg13g2_nand3_1 _1206_ (.B(net113),
    .C(_0527_),
    .A(net141),
    .Y(_0528_));
 sg13g2_nand2b_1 _1207_ (.Y(_0045_),
    .B(_0528_),
    .A_N(_0523_));
 sg13g2_o21ai_1 _1208_ (.B1(net114),
    .Y(_0529_),
    .A1(_0382_),
    .A2(_0438_));
 sg13g2_o21ai_1 _1209_ (.B1(net141),
    .Y(_0530_),
    .A1(_0021_),
    .A2(net120));
 sg13g2_a21oi_1 _1210_ (.A1(_0115_),
    .A2(net120),
    .Y(_0531_),
    .B1(_0530_));
 sg13g2_a21oi_1 _1211_ (.A1(_0098_),
    .A2(net137),
    .Y(_0532_),
    .B1(_0531_));
 sg13g2_and3_1 _1212_ (.X(_0533_),
    .A(_0382_),
    .B(net114),
    .C(_0532_));
 sg13g2_a21o_1 _1213_ (.A2(_0529_),
    .A1(net211),
    .B1(_0533_),
    .X(_0046_));
 sg13g2_nand2_1 _1214_ (.Y(_0534_),
    .A(\system_inst.loader.threshold_min[1] ),
    .B(net137));
 sg13g2_nor2_1 _1215_ (.A(_0114_),
    .B(_0115_),
    .Y(_0535_));
 sg13g2_o21ai_1 _1216_ (.B1(net120),
    .Y(_0536_),
    .A1(_0479_),
    .A2(_0535_));
 sg13g2_o21ai_1 _1217_ (.B1(_0536_),
    .Y(_0537_),
    .A1(_0097_),
    .A2(net119));
 sg13g2_nor2_1 _1218_ (.A(_0365_),
    .B(_0537_),
    .Y(_0538_));
 sg13g2_nor2_1 _1219_ (.A(_0021_),
    .B(_0437_),
    .Y(_0539_));
 sg13g2_o21ai_1 _1220_ (.B1(net141),
    .Y(_0540_),
    .A1(net115),
    .A2(_0539_));
 sg13g2_o21ai_1 _1221_ (.B1(_0534_),
    .Y(_0541_),
    .A1(_0538_),
    .A2(_0540_));
 sg13g2_mux2_1 _1222_ (.A0(_0541_),
    .A1(net209),
    .S(_0529_),
    .X(_0047_));
 sg13g2_nor4_2 _1223_ (.A(\system_inst.loader.current_state[2] ),
    .B(\system_inst.loader.current_state[1] ),
    .C(\system_inst.loader.current_state[6] ),
    .Y(_0542_),
    .D(\system_inst.loader.current_state[4] ));
 sg13g2_nand2_1 _1224_ (.Y(_0543_),
    .A(_0013_),
    .B(_0542_));
 sg13g2_nor2_1 _1225_ (.A(net108),
    .B(_0543_),
    .Y(_0544_));
 sg13g2_o21ai_1 _1226_ (.B1(net1),
    .Y(_0545_),
    .A1(net3),
    .A2(_0117_));
 sg13g2_nor2_1 _1227_ (.A(_0544_),
    .B(_0545_),
    .Y(_0546_));
 sg13g2_and2_1 _1228_ (.A(_0116_),
    .B(_0542_),
    .X(_0547_));
 sg13g2_nand2_1 _1229_ (.Y(_0548_),
    .A(_0116_),
    .B(_0542_));
 sg13g2_o21ai_1 _1230_ (.B1(_0542_),
    .Y(_0549_),
    .A1(_0116_),
    .A2(net134));
 sg13g2_nand2_1 _1231_ (.Y(_0550_),
    .A(net3),
    .B(_0549_));
 sg13g2_nand2_1 _1232_ (.Y(_0551_),
    .A(_0546_),
    .B(_0550_));
 sg13g2_a21oi_1 _1233_ (.A1(net178),
    .A2(_0551_),
    .Y(_0552_),
    .B1(net140));
 sg13g2_o21ai_1 _1234_ (.B1(_0552_),
    .Y(_0048_),
    .A1(_0547_),
    .A2(_0551_));
 sg13g2_o21ai_1 _1235_ (.B1(net147),
    .Y(_0553_),
    .A1(net197),
    .A2(_0130_));
 sg13g2_a21oi_1 _1236_ (.A1(_0094_),
    .A2(_0130_),
    .Y(_0049_),
    .B1(_0553_));
 sg13g2_a21oi_1 _1237_ (.A1(net200),
    .A2(_0129_),
    .Y(_0554_),
    .B1(net139));
 sg13g2_o21ai_1 _1238_ (.B1(_0554_),
    .Y(_0050_),
    .A1(_0092_),
    .A2(_0129_));
 sg13g2_o21ai_1 _1239_ (.B1(net147),
    .Y(_0555_),
    .A1(net194),
    .A2(_0130_));
 sg13g2_a21oi_1 _1240_ (.A1(_0091_),
    .A2(_0130_),
    .Y(_0051_),
    .B1(_0555_));
 sg13g2_o21ai_1 _1241_ (.B1(net147),
    .Y(_0556_),
    .A1(net203),
    .A2(_0135_));
 sg13g2_a21oi_1 _1242_ (.A1(_0094_),
    .A2(_0135_),
    .Y(_0052_),
    .B1(_0556_));
 sg13g2_a21oi_1 _1243_ (.A1(net135),
    .A2(_0134_),
    .Y(_0557_),
    .B1(net139));
 sg13g2_o21ai_1 _1244_ (.B1(_0557_),
    .Y(_0053_),
    .A1(_0092_),
    .A2(_0134_));
 sg13g2_o21ai_1 _1245_ (.B1(net147),
    .Y(_0558_),
    .A1(net199),
    .A2(_0135_));
 sg13g2_a21oi_1 _1246_ (.A1(_0091_),
    .A2(_0135_),
    .Y(_0054_),
    .B1(_0558_));
 sg13g2_o21ai_1 _1247_ (.B1(net143),
    .Y(_0559_),
    .A1(net176),
    .A2(net127));
 sg13g2_a21oi_1 _1248_ (.A1(_0094_),
    .A2(net126),
    .Y(_0055_),
    .B1(_0559_));
 sg13g2_a21oi_1 _1249_ (.A1(\system_inst.loader.shift_reg[0] ),
    .A2(net127),
    .Y(_0560_),
    .B1(net139));
 sg13g2_o21ai_1 _1250_ (.B1(_0560_),
    .Y(_0056_),
    .A1(_0100_),
    .A2(net126));
 sg13g2_o21ai_1 _1251_ (.B1(net147),
    .Y(_0561_),
    .A1(net173),
    .A2(net128));
 sg13g2_a21oi_1 _1252_ (.A1(_0091_),
    .A2(net128),
    .Y(_0057_),
    .B1(_0561_));
 sg13g2_o21ai_1 _1253_ (.B1(net146),
    .Y(_0562_),
    .A1(net195),
    .A2(net128));
 sg13g2_a21oi_1 _1254_ (.A1(_0090_),
    .A2(net128),
    .Y(_0058_),
    .B1(_0562_));
 sg13g2_o21ai_1 _1255_ (.B1(net142),
    .Y(_0563_),
    .A1(\system_inst.leak_rate[4] ),
    .A2(net126));
 sg13g2_a21oi_1 _1256_ (.A1(_0089_),
    .A2(net126),
    .Y(_0059_),
    .B1(_0563_));
 sg13g2_o21ai_1 _1257_ (.B1(net142),
    .Y(_0564_),
    .A1(net163),
    .A2(net126));
 sg13g2_a21oi_1 _1258_ (.A1(_0088_),
    .A2(net126),
    .Y(_0060_),
    .B1(_0564_));
 sg13g2_o21ai_1 _1259_ (.B1(net142),
    .Y(_0565_),
    .A1(net174),
    .A2(net126));
 sg13g2_a21oi_1 _1260_ (.A1(_0087_),
    .A2(net126),
    .Y(_0061_),
    .B1(_0565_));
 sg13g2_o21ai_1 _1261_ (.B1(net142),
    .Y(_0566_),
    .A1(net171),
    .A2(net127));
 sg13g2_a21oi_1 _1262_ (.A1(_0086_),
    .A2(net127),
    .Y(_0062_),
    .B1(_0566_));
 sg13g2_o21ai_1 _1263_ (.B1(net142),
    .Y(_0567_),
    .A1(net216),
    .A2(net130));
 sg13g2_a21oi_1 _1264_ (.A1(_0094_),
    .A2(net130),
    .Y(_0063_),
    .B1(_0567_));
 sg13g2_a21oi_1 _1265_ (.A1(net192),
    .A2(net130),
    .Y(_0568_),
    .B1(net139));
 sg13g2_o21ai_1 _1266_ (.B1(_0568_),
    .Y(_0064_),
    .A1(_0097_),
    .A2(net130));
 sg13g2_a21oi_1 _1267_ (.A1(net196),
    .A2(_0127_),
    .Y(_0569_),
    .B1(net139));
 sg13g2_o21ai_1 _1268_ (.B1(_0569_),
    .Y(_0065_),
    .A1(_0091_),
    .A2(_0127_));
 sg13g2_a21oi_1 _1269_ (.A1(net204),
    .A2(_0127_),
    .Y(_0570_),
    .B1(net139));
 sg13g2_o21ai_1 _1270_ (.B1(_0570_),
    .Y(_0066_),
    .A1(_0090_),
    .A2(_0127_));
 sg13g2_a21oi_1 _1271_ (.A1(net167),
    .A2(net129),
    .Y(_0571_),
    .B1(net138));
 sg13g2_o21ai_1 _1272_ (.B1(_0571_),
    .Y(_0067_),
    .A1(_0096_),
    .A2(net129));
 sg13g2_o21ai_1 _1273_ (.B1(net142),
    .Y(_0572_),
    .A1(net157),
    .A2(net129));
 sg13g2_a21oi_1 _1274_ (.A1(_0088_),
    .A2(net129),
    .Y(_0068_),
    .B1(_0572_));
 sg13g2_o21ai_1 _1275_ (.B1(net142),
    .Y(_0573_),
    .A1(\system_inst.loader.threshold_min[6] ),
    .A2(net129));
 sg13g2_a21oi_1 _1276_ (.A1(_0087_),
    .A2(net129),
    .Y(_0069_),
    .B1(_0573_));
 sg13g2_o21ai_1 _1277_ (.B1(net142),
    .Y(_0574_),
    .A1(net172),
    .A2(net129));
 sg13g2_a21oi_1 _1278_ (.A1(_0086_),
    .A2(net129),
    .Y(_0070_),
    .B1(_0574_));
 sg13g2_and3_2 _1279_ (.X(_0575_),
    .A(net104),
    .B(_0121_),
    .C(_0123_));
 sg13g2_a21oi_1 _1280_ (.A1(net4),
    .A2(_0575_),
    .Y(_0576_),
    .B1(net139));
 sg13g2_o21ai_1 _1281_ (.B1(_0576_),
    .Y(_0071_),
    .A1(_0093_),
    .A2(_0575_));
 sg13g2_o21ai_1 _1282_ (.B1(net145),
    .Y(_0577_),
    .A1(net189),
    .A2(_0575_));
 sg13g2_a21oi_1 _1283_ (.A1(_0092_),
    .A2(_0575_),
    .Y(_0072_),
    .B1(_0577_));
 sg13g2_o21ai_1 _1284_ (.B1(net145),
    .Y(_0578_),
    .A1(net183),
    .A2(_0575_));
 sg13g2_a21oi_1 _1285_ (.A1(_0091_),
    .A2(_0575_),
    .Y(_0073_),
    .B1(_0578_));
 sg13g2_o21ai_1 _1286_ (.B1(net144),
    .Y(_0579_),
    .A1(net193),
    .A2(_0575_));
 sg13g2_a21oi_1 _1287_ (.A1(_0090_),
    .A2(_0575_),
    .Y(_0074_),
    .B1(_0579_));
 sg13g2_nand2b_1 _1288_ (.Y(_0580_),
    .B(_0548_),
    .A_N(net3));
 sg13g2_and2_1 _1289_ (.A(_0546_),
    .B(_0580_),
    .X(_0581_));
 sg13g2_nand2_1 _1290_ (.Y(_0582_),
    .A(_0546_),
    .B(_0580_));
 sg13g2_a21oi_2 _1291_ (.B1(_0547_),
    .Y(_0583_),
    .A2(net134),
    .A1(_0116_));
 sg13g2_a21oi_1 _1292_ (.A1(net4),
    .A2(_0583_),
    .Y(_0584_),
    .B1(_0582_));
 sg13g2_o21ai_1 _1293_ (.B1(net146),
    .Y(_0585_),
    .A1(net192),
    .A2(net123));
 sg13g2_nor2_1 _1294_ (.A(_0584_),
    .B(_0585_),
    .Y(_0075_));
 sg13g2_a21oi_1 _1295_ (.A1(net192),
    .A2(_0583_),
    .Y(_0586_),
    .B1(net122));
 sg13g2_o21ai_1 _1296_ (.B1(net146),
    .Y(_0587_),
    .A1(net169),
    .A2(net123));
 sg13g2_nor2_1 _1297_ (.A(_0586_),
    .B(_0587_),
    .Y(_0076_));
 sg13g2_a21oi_1 _1298_ (.A1(net169),
    .A2(_0583_),
    .Y(_0588_),
    .B1(net122));
 sg13g2_o21ai_1 _1299_ (.B1(net146),
    .Y(_0589_),
    .A1(net154),
    .A2(net123));
 sg13g2_nor2_1 _1300_ (.A(_0588_),
    .B(_0589_),
    .Y(_0077_));
 sg13g2_a21oi_1 _1301_ (.A1(net154),
    .A2(_0583_),
    .Y(_0590_),
    .B1(net122));
 sg13g2_o21ai_1 _1302_ (.B1(net146),
    .Y(_0591_),
    .A1(\system_inst.loader.shift_reg[3] ),
    .A2(net123));
 sg13g2_nor2_1 _1303_ (.A(_0590_),
    .B(_0591_),
    .Y(_0078_));
 sg13g2_a21oi_1 _1304_ (.A1(net167),
    .A2(_0583_),
    .Y(_0592_),
    .B1(net122));
 sg13g2_o21ai_1 _1305_ (.B1(net146),
    .Y(_0593_),
    .A1(net112),
    .A2(net123));
 sg13g2_nor2_1 _1306_ (.A(_0592_),
    .B(_0593_),
    .Y(_0079_));
 sg13g2_a21oi_1 _1307_ (.A1(net112),
    .A2(_0583_),
    .Y(_0594_),
    .B1(net122));
 sg13g2_o21ai_1 _1308_ (.B1(net146),
    .Y(_0595_),
    .A1(\system_inst.loader.shift_reg[5] ),
    .A2(net123));
 sg13g2_nor2_1 _1309_ (.A(_0594_),
    .B(_0595_),
    .Y(_0080_));
 sg13g2_a21oi_1 _1310_ (.A1(net158),
    .A2(_0583_),
    .Y(_0596_),
    .B1(net122));
 sg13g2_o21ai_1 _1311_ (.B1(net146),
    .Y(_0597_),
    .A1(net165),
    .A2(net123));
 sg13g2_nor2_1 _1312_ (.A(_0596_),
    .B(_0597_),
    .Y(_0081_));
 sg13g2_nand3_1 _1313_ (.B(_0546_),
    .C(_0548_),
    .A(net3),
    .Y(_0598_));
 sg13g2_o21ai_1 _1314_ (.B1(net144),
    .Y(_0599_),
    .A1(_0085_),
    .A2(net122));
 sg13g2_a21oi_1 _1315_ (.A1(_0085_),
    .A2(_0598_),
    .Y(_0082_),
    .B1(_0599_));
 sg13g2_a21oi_1 _1316_ (.A1(net106),
    .A2(_0581_),
    .Y(_0600_),
    .B1(net181));
 sg13g2_nand3_1 _1317_ (.B(_0543_),
    .C(_0548_),
    .A(_0120_),
    .Y(_0601_));
 sg13g2_nand2b_1 _1318_ (.Y(_0602_),
    .B(net144),
    .A_N(_0600_));
 sg13g2_a21oi_1 _1319_ (.A1(net123),
    .A2(_0601_),
    .Y(_0083_),
    .B1(_0602_));
 sg13g2_a221oi_1 _1320_ (.B2(_0013_),
    .C1(_0598_),
    .B1(_0542_),
    .A1(_0012_),
    .Y(_0603_),
    .A2(_0120_));
 sg13g2_a22oi_1 _1321_ (.Y(_0604_),
    .B1(_0603_),
    .B2(_0122_),
    .A2(net122),
    .A1(net97));
 sg13g2_nor2_1 _1322_ (.A(net139),
    .B(net98),
    .Y(_0084_));
 sg13g2_dfrbp_1 _1323_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net88),
    .D(_0022_),
    .Q_N(_0653_),
    .Q(\system_inst.neuron.v_mem[0] ));
 sg13g2_dfrbp_1 _1324_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net63),
    .D(_0023_),
    .Q_N(_0652_),
    .Q(\system_inst.neuron.v_mem[1] ));
 sg13g2_dfrbp_1 _1325_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net61),
    .D(_0024_),
    .Q_N(_0651_),
    .Q(\system_inst.neuron.v_mem[2] ));
 sg13g2_dfrbp_1 _1326_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net59),
    .D(_0025_),
    .Q_N(_0650_),
    .Q(\system_inst.neuron.v_mem[3] ));
 sg13g2_dfrbp_1 _1327_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net57),
    .D(_0026_),
    .Q_N(_0649_),
    .Q(\system_inst.neuron.v_mem[4] ));
 sg13g2_dfrbp_1 _1328_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net55),
    .D(_0027_),
    .Q_N(_0648_),
    .Q(\system_inst.neuron.v_mem[5] ));
 sg13g2_dfrbp_1 _1329_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net53),
    .D(_0028_),
    .Q_N(_0647_),
    .Q(\system_inst.neuron.v_mem[6] ));
 sg13g2_dfrbp_1 _1330_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net51),
    .D(_0029_),
    .Q_N(_0646_),
    .Q(\system_inst.neuron.v_mem[7] ));
 sg13g2_dfrbp_1 _1331_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net49),
    .D(_0030_),
    .Q_N(_0645_),
    .Q(\system_inst.neuron.v_mem[8] ));
 sg13g2_dfrbp_1 _1332_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net47),
    .D(_0031_),
    .Q_N(_0644_),
    .Q(spike_out));
 sg13g2_dfrbp_1 _1333_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net46),
    .D(_0032_),
    .Q_N(_0643_),
    .Q(\system_inst.neuron.refr_cnt[0] ));
 sg13g2_dfrbp_1 _1334_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net44),
    .D(_0033_),
    .Q_N(_0642_),
    .Q(\system_inst.neuron.refr_cnt[1] ));
 sg13g2_dfrbp_1 _1335_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net42),
    .D(_0034_),
    .Q_N(_0641_),
    .Q(\system_inst.neuron.refr_cnt[2] ));
 sg13g2_dfrbp_1 _1336_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net40),
    .D(net96),
    .Q_N(_0640_),
    .Q(\system_inst.neuron.refr_cnt[3] ));
 sg13g2_dfrbp_1 _1337_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net38),
    .D(net111),
    .Q_N(_0020_),
    .Q(\system_inst.neuron.leak_counter[0] ));
 sg13g2_dfrbp_1 _1338_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net36),
    .D(net101),
    .Q_N(_0639_),
    .Q(\system_inst.neuron.leak_counter[1] ));
 sg13g2_dfrbp_1 _1339_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net34),
    .D(_0038_),
    .Q_N(_0638_),
    .Q(\system_inst.neuron.leak_counter[2] ));
 sg13g2_dfrbp_1 _1340_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net32),
    .D(_0039_),
    .Q_N(_0637_),
    .Q(\system_inst.neuron.leak_counter[3] ));
 sg13g2_dfrbp_1 _1341_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net30),
    .D(_0040_),
    .Q_N(_0010_),
    .Q(\system_inst.neuron.threshold[2] ));
 sg13g2_dfrbp_1 _1342_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net29),
    .D(_0041_),
    .Q_N(_0009_),
    .Q(\system_inst.neuron.threshold[3] ));
 sg13g2_dfrbp_1 _1343_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net28),
    .D(_0042_),
    .Q_N(_0016_),
    .Q(\system_inst.neuron.threshold[4] ));
 sg13g2_dfrbp_1 _1344_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net27),
    .D(_0043_),
    .Q_N(_0008_),
    .Q(\system_inst.neuron.threshold[5] ));
 sg13g2_dfrbp_1 _1345_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net26),
    .D(_0044_),
    .Q_N(_0007_),
    .Q(\system_inst.neuron.threshold[6] ));
 sg13g2_dfrbp_1 _1346_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net25),
    .D(_0045_),
    .Q_N(_0006_),
    .Q(\system_inst.neuron.threshold[7] ));
 sg13g2_dfrbp_1 _1347_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net87),
    .D(_0046_),
    .Q_N(_0636_),
    .Q(\system_inst.neuron.threshold[0] ));
 sg13g2_dfrbp_1 _1348_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net86),
    .D(net210),
    .Q_N(_0011_),
    .Q(\system_inst.neuron.threshold[1] ));
 sg13g2_dfrbp_1 _1349_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net85),
    .D(net179),
    .Q_N(_0635_),
    .Q(params_ready));
 sg13g2_dfrbp_1 _1350_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net83),
    .D(_0049_),
    .Q_N(_0634_),
    .Q(\system_inst.loader.weight_a[0] ));
 sg13g2_dfrbp_1 _1351_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net81),
    .D(_0050_),
    .Q_N(_0633_),
    .Q(\system_inst.loader.weight_a[1] ));
 sg13g2_dfrbp_1 _1352_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net79),
    .D(_0051_),
    .Q_N(_0632_),
    .Q(\system_inst.loader.weight_a[2] ));
 sg13g2_dfrbp_1 _1353_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net77),
    .D(_0052_),
    .Q_N(_0631_),
    .Q(\system_inst.loader.weight_b[0] ));
 sg13g2_dfrbp_1 _1354_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net75),
    .D(_0053_),
    .Q_N(_0630_),
    .Q(\system_inst.loader.weight_b[1] ));
 sg13g2_dfrbp_1 _1355_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net73),
    .D(_0054_),
    .Q_N(_0629_),
    .Q(\system_inst.loader.weight_b[2] ));
 sg13g2_dfrbp_1 _1356_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net71),
    .D(_0055_),
    .Q_N(_0628_),
    .Q(\system_inst.leak_rate[0] ));
 sg13g2_dfrbp_1 _1357_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net69),
    .D(net162),
    .Q_N(_0627_),
    .Q(\system_inst.leak_rate[1] ));
 sg13g2_dfrbp_1 _1358_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net67),
    .D(_0057_),
    .Q_N(_0626_),
    .Q(\system_inst.leak_rate[2] ));
 sg13g2_dfrbp_1 _1359_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net65),
    .D(_0058_),
    .Q_N(_0625_),
    .Q(\system_inst.leak_rate[3] ));
 sg13g2_dfrbp_1 _1360_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net62),
    .D(net168),
    .Q_N(_0624_),
    .Q(\system_inst.leak_rate[4] ));
 sg13g2_dfrbp_1 _1361_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net58),
    .D(_0060_),
    .Q_N(_0623_),
    .Q(\system_inst.leak_rate[5] ));
 sg13g2_dfrbp_1 _1362_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net54),
    .D(_0061_),
    .Q_N(_0622_),
    .Q(\system_inst.leak_rate[6] ));
 sg13g2_dfrbp_1 _1363_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net50),
    .D(_0062_),
    .Q_N(_0621_),
    .Q(\system_inst.leak_rate[7] ));
 sg13g2_dfrbp_1 _1364_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net45),
    .D(_0063_),
    .Q_N(_0021_),
    .Q(\system_inst.loader.threshold_min[0] ));
 sg13g2_dfrbp_1 _1365_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net41),
    .D(_0064_),
    .Q_N(_0620_),
    .Q(\system_inst.loader.threshold_min[1] ));
 sg13g2_dfrbp_1 _1366_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net37),
    .D(_0065_),
    .Q_N(_0014_),
    .Q(\system_inst.loader.threshold_min[2] ));
 sg13g2_dfrbp_1 _1367_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net33),
    .D(_0066_),
    .Q_N(_0015_),
    .Q(\system_inst.loader.threshold_min[3] ));
 sg13g2_dfrbp_1 _1368_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net84),
    .D(_0067_),
    .Q_N(_0017_),
    .Q(\system_inst.loader.threshold_min[4] ));
 sg13g2_dfrbp_1 _1369_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net80),
    .D(_0068_),
    .Q_N(_0018_),
    .Q(\system_inst.loader.threshold_min[5] ));
 sg13g2_dfrbp_1 _1370_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net76),
    .D(net159),
    .Q_N(_0019_),
    .Q(\system_inst.loader.threshold_min[6] ));
 sg13g2_dfrbp_1 _1371_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net72),
    .D(_0070_),
    .Q_N(_0619_),
    .Q(\system_inst.loader.threshold_min[7] ));
 sg13g2_dfrbp_1 _1372_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net68),
    .D(net103),
    .Q_N(_0618_),
    .Q(\system_inst.leak_cycles[0] ));
 sg13g2_dfrbp_1 _1373_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net64),
    .D(net190),
    .Q_N(_0617_),
    .Q(\system_inst.leak_cycles[1] ));
 sg13g2_dfrbp_1 _1374_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net56),
    .D(net184),
    .Q_N(_0616_),
    .Q(\system_inst.leak_cycles[2] ));
 sg13g2_dfrbp_1 _1375_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net48),
    .D(_0074_),
    .Q_N(_0615_),
    .Q(\system_inst.leak_cycles[3] ));
 sg13g2_dfrbp_1 _1376_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net39),
    .D(_0075_),
    .Q_N(_0614_),
    .Q(\system_inst.loader.shift_reg[0] ));
 sg13g2_dfrbp_1 _1377_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net31),
    .D(_0076_),
    .Q_N(_0613_),
    .Q(\system_inst.loader.shift_reg[1] ));
 sg13g2_dfrbp_1 _1378_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net78),
    .D(_0077_),
    .Q_N(_0612_),
    .Q(\system_inst.loader.shift_reg[2] ));
 sg13g2_dfrbp_1 _1379_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net70),
    .D(net155),
    .Q_N(_0611_),
    .Q(\system_inst.loader.shift_reg[3] ));
 sg13g2_dfrbp_1 _1380_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net60),
    .D(_0079_),
    .Q_N(_0610_),
    .Q(\system_inst.loader.shift_reg[4] ));
 sg13g2_dfrbp_1 _1381_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net43),
    .D(net149),
    .Q_N(_0609_),
    .Q(\system_inst.loader.shift_reg[5] ));
 sg13g2_dfrbp_1 _1382_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net82),
    .D(_0081_),
    .Q_N(_0608_),
    .Q(\system_inst.loader.shift_reg[6] ));
 sg13g2_dfrbp_1 _1383_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net66),
    .D(net107),
    .Q_N(_0607_),
    .Q(\system_inst.loader.bit_count[0] ));
 sg13g2_dfrbp_1 _1384_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net35),
    .D(net182),
    .Q_N(_0606_),
    .Q(\system_inst.loader.bit_count[1] ));
 sg13g2_dfrbp_1 _1385_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net89),
    .D(_0084_),
    .Q_N(_0012_),
    .Q(\system_inst.loader.bit_count[2] ));
 sg13g2_dfrbp_1 _1386_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net90),
    .D(_0000_),
    .Q_N(_0654_),
    .Q(\system_inst.loader.current_state[0] ));
 sg13g2_dfrbp_1 _1387_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net91),
    .D(_0001_),
    .Q_N(_0655_),
    .Q(\system_inst.loader.current_state[1] ));
 sg13g2_dfrbp_1 _1388_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net92),
    .D(_0002_),
    .Q_N(_0656_),
    .Q(\system_inst.loader.current_state[2] ));
 sg13g2_dfrbp_1 _1389_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net93),
    .D(_0003_),
    .Q_N(_0657_),
    .Q(\system_inst.loader.current_state[4] ));
 sg13g2_dfrbp_1 _1390_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net74),
    .D(_0004_),
    .Q_N(_0013_),
    .Q(\system_inst.loader.current_state[5] ));
 sg13g2_dfrbp_1 _1391_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net52),
    .D(_0005_),
    .Q_N(_0605_),
    .Q(\system_inst.loader.current_state[6] ));
 sg13g2_tiehi _1345__26 (.L_HI(net26));
 sg13g2_tiehi _1344__27 (.L_HI(net27));
 sg13g2_tiehi _1343__28 (.L_HI(net28));
 sg13g2_tiehi _1342__29 (.L_HI(net29));
 sg13g2_tiehi _1341__30 (.L_HI(net30));
 sg13g2_tiehi _1377__31 (.L_HI(net31));
 sg13g2_tiehi _1340__32 (.L_HI(net32));
 sg13g2_tiehi _1367__33 (.L_HI(net33));
 sg13g2_tiehi _1339__34 (.L_HI(net34));
 sg13g2_tiehi _1384__35 (.L_HI(net35));
 sg13g2_tiehi _1338__36 (.L_HI(net36));
 sg13g2_tiehi _1366__37 (.L_HI(net37));
 sg13g2_tiehi _1337__38 (.L_HI(net38));
 sg13g2_tiehi _1376__39 (.L_HI(net39));
 sg13g2_tiehi _1336__40 (.L_HI(net40));
 sg13g2_tiehi _1365__41 (.L_HI(net41));
 sg13g2_tiehi _1335__42 (.L_HI(net42));
 sg13g2_tiehi _1381__43 (.L_HI(net43));
 sg13g2_tiehi _1334__44 (.L_HI(net44));
 sg13g2_tiehi _1364__45 (.L_HI(net45));
 sg13g2_tiehi _1333__46 (.L_HI(net46));
 sg13g2_tiehi _1332__47 (.L_HI(net47));
 sg13g2_tiehi _1375__48 (.L_HI(net48));
 sg13g2_tiehi _1331__49 (.L_HI(net49));
 sg13g2_tiehi _1363__50 (.L_HI(net50));
 sg13g2_tiehi _1330__51 (.L_HI(net51));
 sg13g2_tiehi _1391__52 (.L_HI(net52));
 sg13g2_tiehi _1329__53 (.L_HI(net53));
 sg13g2_tiehi _1362__54 (.L_HI(net54));
 sg13g2_tiehi _1328__55 (.L_HI(net55));
 sg13g2_tiehi _1374__56 (.L_HI(net56));
 sg13g2_tiehi _1327__57 (.L_HI(net57));
 sg13g2_tiehi _1361__58 (.L_HI(net58));
 sg13g2_tiehi _1326__59 (.L_HI(net59));
 sg13g2_tiehi _1380__60 (.L_HI(net60));
 sg13g2_tiehi _1325__61 (.L_HI(net61));
 sg13g2_tiehi _1360__62 (.L_HI(net62));
 sg13g2_tiehi _1324__63 (.L_HI(net63));
 sg13g2_tiehi _1373__64 (.L_HI(net64));
 sg13g2_tiehi _1359__65 (.L_HI(net65));
 sg13g2_tiehi _1383__66 (.L_HI(net66));
 sg13g2_tiehi _1358__67 (.L_HI(net67));
 sg13g2_tiehi _1372__68 (.L_HI(net68));
 sg13g2_tiehi _1357__69 (.L_HI(net69));
 sg13g2_tiehi _1379__70 (.L_HI(net70));
 sg13g2_tiehi _1356__71 (.L_HI(net71));
 sg13g2_tiehi _1371__72 (.L_HI(net72));
 sg13g2_tiehi _1355__73 (.L_HI(net73));
 sg13g2_tiehi _1390__74 (.L_HI(net74));
 sg13g2_tiehi _1354__75 (.L_HI(net75));
 sg13g2_tiehi _1370__76 (.L_HI(net76));
 sg13g2_tiehi _1353__77 (.L_HI(net77));
 sg13g2_tiehi _1378__78 (.L_HI(net78));
 sg13g2_tiehi _1352__79 (.L_HI(net79));
 sg13g2_tiehi _1369__80 (.L_HI(net80));
 sg13g2_tiehi _1351__81 (.L_HI(net81));
 sg13g2_tiehi _1382__82 (.L_HI(net82));
 sg13g2_tiehi _1350__83 (.L_HI(net83));
 sg13g2_tiehi _1368__84 (.L_HI(net84));
 sg13g2_tiehi _1349__85 (.L_HI(net85));
 sg13g2_tiehi _1348__86 (.L_HI(net86));
 sg13g2_tiehi _1347__87 (.L_HI(net87));
 sg13g2_tiehi _1323__88 (.L_HI(net88));
 sg13g2_tiehi _1385__89 (.L_HI(net89));
 sg13g2_tiehi _1386__90 (.L_HI(net90));
 sg13g2_tiehi _1387__91 (.L_HI(net91));
 sg13g2_tiehi _1388__92 (.L_HI(net92));
 sg13g2_tiehi _1389__93 (.L_HI(net93));
 sg13g2_tiehi tt_um_alif_dual_unileak_94 (.L_HI(net94));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_alif_dual_unileak_12 (.L_LO(net12));
 sg13g2_tielo tt_um_alif_dual_unileak_13 (.L_LO(net13));
 sg13g2_tielo tt_um_alif_dual_unileak_14 (.L_LO(net14));
 sg13g2_tielo tt_um_alif_dual_unileak_15 (.L_LO(net15));
 sg13g2_tielo tt_um_alif_dual_unileak_16 (.L_LO(net16));
 sg13g2_tielo tt_um_alif_dual_unileak_17 (.L_LO(net17));
 sg13g2_tielo tt_um_alif_dual_unileak_18 (.L_LO(net18));
 sg13g2_tielo tt_um_alif_dual_unileak_19 (.L_LO(net19));
 sg13g2_tielo tt_um_alif_dual_unileak_20 (.L_LO(net20));
 sg13g2_tielo tt_um_alif_dual_unileak_21 (.L_LO(net21));
 sg13g2_tielo tt_um_alif_dual_unileak_22 (.L_LO(net22));
 sg13g2_tielo tt_um_alif_dual_unileak_23 (.L_LO(net23));
 sg13g2_tielo tt_um_alif_dual_unileak_24 (.L_LO(net24));
 sg13g2_tiehi _1346__25 (.L_HI(net25));
 sg13g2_buf_2 _1476_ (.A(params_ready),
    .X(uio_out[0]));
 sg13g2_buf_2 _1477_ (.A(spike_out),
    .X(uo_out[0]));
 sg13g2_buf_4 fanout113 (.X(net113),
    .A(_0403_));
 sg13g2_buf_2 fanout114 (.A(_0403_),
    .X(net114));
 sg13g2_buf_4 fanout115 (.X(net115),
    .A(net116));
 sg13g2_buf_4 fanout116 (.X(net116),
    .A(_0364_));
 sg13g2_buf_2 fanout117 (.A(net118),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_0301_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_0478_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_0478_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_0437_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_0582_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_0581_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(net125),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_0293_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(net128),
    .X(net126));
 sg13g2_buf_1 fanout127 (.A(net128),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_0132_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_0126_),
    .X(net129));
 sg13g2_buf_1 fanout130 (.A(_0126_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(net132),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_0145_),
    .X(net132));
 sg13g2_buf_1 fanout133 (.A(_0145_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_0121_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(net198),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(net214),
    .X(net136));
 sg13g2_buf_4 fanout137 (.X(net137),
    .A(net138));
 sg13g2_buf_4 fanout138 (.X(net138),
    .A(net140));
 sg13g2_buf_2 fanout139 (.A(net140),
    .X(net139));
 sg13g2_buf_4 fanout140 (.X(net140),
    .A(_0118_));
 sg13g2_buf_4 fanout141 (.X(net141),
    .A(net143));
 sg13g2_buf_2 fanout142 (.A(net143),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(rst_n),
    .X(net143));
 sg13g2_buf_4 fanout144 (.X(net144),
    .A(net148));
 sg13g2_buf_2 fanout145 (.A(net148),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(net148),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(net148),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(rst_n),
    .X(net148));
 sg13g2_buf_2 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_buf_2 input10 (.A(uio_in[0]),
    .X(net10));
 sg13g2_tielo tt_um_alif_dual_unileak_11 (.L_LO(net11));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_10_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\system_inst.neuron.refr_cnt[3] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0035_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold3 (.A(\system_inst.loader.bit_count[2] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0604_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold5 (.A(\system_inst.neuron.leak_counter[1] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0399_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0037_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold8 (.A(\system_inst.leak_cycles[0] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0071_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold10 (.A(\system_inst.loader.current_state[5] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0128_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold12 (.A(\system_inst.loader.bit_count[0] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0082_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold14 (.A(\system_inst.loader.current_state[0] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0020_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0394_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0036_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold18 (.A(\system_inst.loader.shift_reg[4] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0080_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold20 (.A(\system_inst.loader.current_state[2] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0131_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold22 (.A(\system_inst.loader.current_state[6] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold23 (.A(\system_inst.neuron.v_mem[7] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold24 (.A(\system_inst.loader.shift_reg[2] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0078_),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold26 (.A(\system_inst.loader.current_state[4] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold27 (.A(\system_inst.loader.threshold_min[5] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold28 (.A(\system_inst.loader.shift_reg[5] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0069_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold30 (.A(\system_inst.neuron.v_mem[2] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold31 (.A(\system_inst.leak_rate[1] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0056_),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold33 (.A(\system_inst.leak_rate[5] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold34 (.A(\system_inst.neuron.v_mem[1] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold35 (.A(\system_inst.loader.shift_reg[6] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold36 (.A(\system_inst.loader.current_state[1] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold37 (.A(\system_inst.loader.shift_reg[3] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0059_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold39 (.A(\system_inst.loader.shift_reg[1] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold40 (.A(\system_inst.neuron.v_mem[0] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold41 (.A(\system_inst.leak_rate[7] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold42 (.A(\system_inst.loader.threshold_min[7] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold43 (.A(\system_inst.leak_rate[2] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold44 (.A(\system_inst.leak_rate[6] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold45 (.A(\system_inst.neuron.v_mem[6] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold46 (.A(\system_inst.leak_rate[0] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold47 (.A(\system_inst.neuron.v_mem[5] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold48 (.A(params_ready),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0048_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold50 (.A(\system_inst.neuron.v_mem[4] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold51 (.A(\system_inst.loader.bit_count[1] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0083_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold53 (.A(\system_inst.leak_cycles[2] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0073_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold55 (.A(\system_inst.neuron.leak_counter[3] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0402_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold57 (.A(\system_inst.neuron.leak_counter[2] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0401_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold59 (.A(\system_inst.leak_cycles[1] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0072_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold61 (.A(\system_inst.neuron.v_mem[3] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold62 (.A(\system_inst.loader.shift_reg[0] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold63 (.A(\system_inst.leak_cycles[3] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold64 (.A(\system_inst.loader.weight_a[2] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold65 (.A(\system_inst.leak_rate[3] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold66 (.A(\system_inst.loader.threshold_min[2] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold67 (.A(\system_inst.loader.weight_a[0] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold68 (.A(\system_inst.loader.weight_b[1] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold69 (.A(\system_inst.loader.weight_b[2] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold70 (.A(\system_inst.loader.weight_a[1] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold71 (.A(\system_inst.loader.threshold_min[4] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold72 (.A(\system_inst.neuron.threshold[4] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold73 (.A(\system_inst.loader.weight_b[0] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold74 (.A(\system_inst.loader.threshold_min[3] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold75 (.A(\system_inst.neuron.refr_cnt[2] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0391_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold77 (.A(\system_inst.neuron.refr_cnt[0] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold78 (.A(\system_inst.neuron.threshold[5] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold79 (.A(\system_inst.neuron.threshold[1] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0047_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold81 (.A(\system_inst.neuron.threshold[0] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold82 (.A(\system_inst.neuron.threshold[7] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold83 (.A(\system_inst.loader.threshold_min[1] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold84 (.A(\system_inst.neuron.v_mem[8] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold85 (.A(\system_inst.neuron.refr_cnt[1] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold86 (.A(\system_inst.loader.threshold_min[0] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold87 (.A(\system_inst.loader.threshold_min[6] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0521_),
    .X(net218));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_fill_2 FILLER_13_56 ();
 sg13g2_fill_1 FILLER_13_58 ();
 sg13g2_decap_8 FILLER_13_85 ();
 sg13g2_decap_8 FILLER_13_92 ();
 sg13g2_decap_4 FILLER_13_99 ();
 sg13g2_fill_2 FILLER_13_103 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_4 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_233 ();
 sg13g2_decap_8 FILLER_13_240 ();
 sg13g2_decap_8 FILLER_13_247 ();
 sg13g2_decap_8 FILLER_13_254 ();
 sg13g2_decap_8 FILLER_13_261 ();
 sg13g2_decap_8 FILLER_13_268 ();
 sg13g2_decap_8 FILLER_13_275 ();
 sg13g2_decap_8 FILLER_13_282 ();
 sg13g2_decap_8 FILLER_13_289 ();
 sg13g2_decap_8 FILLER_13_296 ();
 sg13g2_decap_8 FILLER_13_303 ();
 sg13g2_decap_8 FILLER_13_310 ();
 sg13g2_decap_8 FILLER_13_317 ();
 sg13g2_decap_8 FILLER_13_324 ();
 sg13g2_decap_8 FILLER_13_331 ();
 sg13g2_decap_8 FILLER_13_338 ();
 sg13g2_decap_8 FILLER_13_345 ();
 sg13g2_decap_8 FILLER_13_352 ();
 sg13g2_decap_8 FILLER_13_359 ();
 sg13g2_decap_8 FILLER_13_366 ();
 sg13g2_decap_8 FILLER_13_373 ();
 sg13g2_decap_8 FILLER_13_380 ();
 sg13g2_decap_8 FILLER_13_387 ();
 sg13g2_decap_8 FILLER_13_394 ();
 sg13g2_decap_8 FILLER_13_401 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_fill_1 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_61 ();
 sg13g2_fill_2 FILLER_14_68 ();
 sg13g2_decap_8 FILLER_14_74 ();
 sg13g2_fill_2 FILLER_14_81 ();
 sg13g2_fill_1 FILLER_14_83 ();
 sg13g2_decap_8 FILLER_14_129 ();
 sg13g2_decap_8 FILLER_14_136 ();
 sg13g2_decap_4 FILLER_14_143 ();
 sg13g2_fill_1 FILLER_14_147 ();
 sg13g2_fill_2 FILLER_14_152 ();
 sg13g2_fill_1 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_225 ();
 sg13g2_decap_8 FILLER_14_232 ();
 sg13g2_decap_8 FILLER_14_239 ();
 sg13g2_decap_8 FILLER_14_246 ();
 sg13g2_decap_8 FILLER_14_253 ();
 sg13g2_decap_8 FILLER_14_260 ();
 sg13g2_decap_8 FILLER_14_267 ();
 sg13g2_decap_8 FILLER_14_274 ();
 sg13g2_decap_8 FILLER_14_281 ();
 sg13g2_fill_2 FILLER_14_288 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_fill_1 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_349 ();
 sg13g2_decap_8 FILLER_14_356 ();
 sg13g2_decap_8 FILLER_14_363 ();
 sg13g2_decap_8 FILLER_14_370 ();
 sg13g2_decap_8 FILLER_14_377 ();
 sg13g2_decap_8 FILLER_14_384 ();
 sg13g2_decap_8 FILLER_14_391 ();
 sg13g2_decap_8 FILLER_14_398 ();
 sg13g2_decap_4 FILLER_14_405 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_4 FILLER_15_35 ();
 sg13g2_fill_2 FILLER_15_65 ();
 sg13g2_fill_2 FILLER_15_85 ();
 sg13g2_fill_1 FILLER_15_87 ();
 sg13g2_decap_4 FILLER_15_97 ();
 sg13g2_fill_1 FILLER_15_101 ();
 sg13g2_decap_4 FILLER_15_117 ();
 sg13g2_decap_4 FILLER_15_133 ();
 sg13g2_decap_4 FILLER_15_163 ();
 sg13g2_fill_2 FILLER_15_180 ();
 sg13g2_fill_1 FILLER_15_182 ();
 sg13g2_fill_2 FILLER_15_188 ();
 sg13g2_fill_1 FILLER_15_215 ();
 sg13g2_fill_2 FILLER_15_225 ();
 sg13g2_fill_1 FILLER_15_227 ();
 sg13g2_decap_8 FILLER_15_254 ();
 sg13g2_fill_1 FILLER_15_261 ();
 sg13g2_decap_4 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_305 ();
 sg13g2_fill_1 FILLER_15_338 ();
 sg13g2_decap_8 FILLER_15_374 ();
 sg13g2_decap_8 FILLER_15_381 ();
 sg13g2_decap_8 FILLER_15_388 ();
 sg13g2_decap_8 FILLER_15_395 ();
 sg13g2_decap_8 FILLER_15_402 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_fill_2 FILLER_16_35 ();
 sg13g2_fill_1 FILLER_16_37 ();
 sg13g2_fill_2 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_4 FILLER_16_70 ();
 sg13g2_fill_2 FILLER_16_74 ();
 sg13g2_fill_2 FILLER_16_105 ();
 sg13g2_fill_1 FILLER_16_107 ();
 sg13g2_decap_4 FILLER_16_119 ();
 sg13g2_fill_1 FILLER_16_123 ();
 sg13g2_fill_1 FILLER_16_132 ();
 sg13g2_decap_8 FILLER_16_146 ();
 sg13g2_decap_8 FILLER_16_153 ();
 sg13g2_fill_2 FILLER_16_160 ();
 sg13g2_fill_2 FILLER_16_185 ();
 sg13g2_fill_1 FILLER_16_187 ();
 sg13g2_fill_2 FILLER_16_193 ();
 sg13g2_fill_1 FILLER_16_195 ();
 sg13g2_fill_1 FILLER_16_216 ();
 sg13g2_decap_8 FILLER_16_244 ();
 sg13g2_fill_1 FILLER_16_277 ();
 sg13g2_decap_8 FILLER_16_300 ();
 sg13g2_decap_4 FILLER_16_307 ();
 sg13g2_decap_4 FILLER_16_342 ();
 sg13g2_decap_8 FILLER_16_368 ();
 sg13g2_decap_8 FILLER_16_375 ();
 sg13g2_decap_8 FILLER_16_382 ();
 sg13g2_decap_8 FILLER_16_389 ();
 sg13g2_decap_8 FILLER_16_396 ();
 sg13g2_decap_4 FILLER_16_403 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_fill_2 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_20 ();
 sg13g2_decap_4 FILLER_17_27 ();
 sg13g2_decap_8 FILLER_17_54 ();
 sg13g2_fill_1 FILLER_17_61 ();
 sg13g2_fill_1 FILLER_17_67 ();
 sg13g2_decap_8 FILLER_17_75 ();
 sg13g2_decap_8 FILLER_17_82 ();
 sg13g2_decap_8 FILLER_17_101 ();
 sg13g2_fill_2 FILLER_17_118 ();
 sg13g2_decap_8 FILLER_17_124 ();
 sg13g2_decap_4 FILLER_17_131 ();
 sg13g2_fill_2 FILLER_17_135 ();
 sg13g2_decap_4 FILLER_17_145 ();
 sg13g2_fill_2 FILLER_17_149 ();
 sg13g2_decap_4 FILLER_17_177 ();
 sg13g2_decap_8 FILLER_17_191 ();
 sg13g2_fill_2 FILLER_17_207 ();
 sg13g2_fill_1 FILLER_17_209 ();
 sg13g2_decap_8 FILLER_17_219 ();
 sg13g2_fill_2 FILLER_17_230 ();
 sg13g2_decap_4 FILLER_17_237 ();
 sg13g2_fill_1 FILLER_17_241 ();
 sg13g2_fill_2 FILLER_17_260 ();
 sg13g2_fill_1 FILLER_17_267 ();
 sg13g2_fill_1 FILLER_17_282 ();
 sg13g2_fill_2 FILLER_17_315 ();
 sg13g2_fill_1 FILLER_17_333 ();
 sg13g2_fill_2 FILLER_17_339 ();
 sg13g2_decap_8 FILLER_17_361 ();
 sg13g2_decap_8 FILLER_17_368 ();
 sg13g2_decap_8 FILLER_17_375 ();
 sg13g2_decap_8 FILLER_17_382 ();
 sg13g2_decap_8 FILLER_17_389 ();
 sg13g2_decap_8 FILLER_17_396 ();
 sg13g2_decap_4 FILLER_17_403 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_4 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_4 ();
 sg13g2_fill_1 FILLER_18_31 ();
 sg13g2_decap_4 FILLER_18_70 ();
 sg13g2_fill_2 FILLER_18_74 ();
 sg13g2_fill_2 FILLER_18_81 ();
 sg13g2_decap_8 FILLER_18_96 ();
 sg13g2_fill_2 FILLER_18_103 ();
 sg13g2_fill_2 FILLER_18_115 ();
 sg13g2_fill_1 FILLER_18_117 ();
 sg13g2_decap_8 FILLER_18_153 ();
 sg13g2_decap_4 FILLER_18_160 ();
 sg13g2_fill_1 FILLER_18_164 ();
 sg13g2_decap_8 FILLER_18_183 ();
 sg13g2_fill_2 FILLER_18_190 ();
 sg13g2_fill_2 FILLER_18_218 ();
 sg13g2_fill_1 FILLER_18_251 ();
 sg13g2_decap_4 FILLER_18_291 ();
 sg13g2_fill_2 FILLER_18_295 ();
 sg13g2_fill_1 FILLER_18_309 ();
 sg13g2_decap_4 FILLER_18_341 ();
 sg13g2_fill_1 FILLER_18_345 ();
 sg13g2_decap_4 FILLER_18_355 ();
 sg13g2_decap_8 FILLER_18_390 ();
 sg13g2_decap_8 FILLER_18_397 ();
 sg13g2_decap_4 FILLER_18_404 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_fill_2 FILLER_19_14 ();
 sg13g2_fill_1 FILLER_19_16 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_4 FILLER_19_61 ();
 sg13g2_fill_2 FILLER_19_65 ();
 sg13g2_decap_4 FILLER_19_71 ();
 sg13g2_fill_2 FILLER_19_75 ();
 sg13g2_fill_2 FILLER_19_93 ();
 sg13g2_fill_1 FILLER_19_95 ();
 sg13g2_fill_1 FILLER_19_111 ();
 sg13g2_decap_8 FILLER_19_125 ();
 sg13g2_fill_2 FILLER_19_132 ();
 sg13g2_fill_1 FILLER_19_134 ();
 sg13g2_fill_1 FILLER_19_139 ();
 sg13g2_fill_1 FILLER_19_146 ();
 sg13g2_fill_1 FILLER_19_181 ();
 sg13g2_fill_2 FILLER_19_187 ();
 sg13g2_decap_4 FILLER_19_202 ();
 sg13g2_fill_2 FILLER_19_206 ();
 sg13g2_fill_1 FILLER_19_216 ();
 sg13g2_fill_1 FILLER_19_222 ();
 sg13g2_fill_2 FILLER_19_244 ();
 sg13g2_fill_1 FILLER_19_246 ();
 sg13g2_decap_4 FILLER_19_251 ();
 sg13g2_fill_1 FILLER_19_255 ();
 sg13g2_fill_2 FILLER_19_261 ();
 sg13g2_fill_1 FILLER_19_263 ();
 sg13g2_decap_8 FILLER_19_277 ();
 sg13g2_fill_1 FILLER_19_284 ();
 sg13g2_fill_1 FILLER_19_296 ();
 sg13g2_fill_1 FILLER_19_330 ();
 sg13g2_decap_4 FILLER_19_341 ();
 sg13g2_fill_2 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_391 ();
 sg13g2_decap_8 FILLER_19_398 ();
 sg13g2_decap_4 FILLER_19_405 ();
 sg13g2_decap_4 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_4 ();
 sg13g2_fill_2 FILLER_20_32 ();
 sg13g2_decap_8 FILLER_20_69 ();
 sg13g2_decap_4 FILLER_20_76 ();
 sg13g2_decap_8 FILLER_20_92 ();
 sg13g2_decap_8 FILLER_20_99 ();
 sg13g2_fill_2 FILLER_20_106 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_fill_2 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_fill_1 FILLER_20_161 ();
 sg13g2_fill_2 FILLER_20_174 ();
 sg13g2_decap_8 FILLER_20_180 ();
 sg13g2_fill_2 FILLER_20_187 ();
 sg13g2_fill_1 FILLER_20_189 ();
 sg13g2_decap_4 FILLER_20_226 ();
 sg13g2_fill_1 FILLER_20_256 ();
 sg13g2_decap_4 FILLER_20_262 ();
 sg13g2_decap_4 FILLER_20_269 ();
 sg13g2_decap_8 FILLER_20_277 ();
 sg13g2_decap_8 FILLER_20_284 ();
 sg13g2_decap_8 FILLER_20_291 ();
 sg13g2_fill_2 FILLER_20_298 ();
 sg13g2_fill_1 FILLER_20_300 ();
 sg13g2_decap_4 FILLER_20_304 ();
 sg13g2_decap_8 FILLER_20_319 ();
 sg13g2_decap_8 FILLER_20_326 ();
 sg13g2_decap_8 FILLER_20_333 ();
 sg13g2_decap_8 FILLER_20_340 ();
 sg13g2_fill_2 FILLER_20_355 ();
 sg13g2_fill_2 FILLER_20_361 ();
 sg13g2_decap_8 FILLER_20_389 ();
 sg13g2_decap_8 FILLER_20_396 ();
 sg13g2_decap_4 FILLER_20_403 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_fill_2 FILLER_21_28 ();
 sg13g2_fill_1 FILLER_21_30 ();
 sg13g2_decap_8 FILLER_21_55 ();
 sg13g2_fill_1 FILLER_21_62 ();
 sg13g2_decap_8 FILLER_21_71 ();
 sg13g2_fill_2 FILLER_21_78 ();
 sg13g2_fill_2 FILLER_21_95 ();
 sg13g2_fill_1 FILLER_21_97 ();
 sg13g2_decap_8 FILLER_21_125 ();
 sg13g2_fill_2 FILLER_21_132 ();
 sg13g2_fill_1 FILLER_21_134 ();
 sg13g2_decap_4 FILLER_21_147 ();
 sg13g2_fill_2 FILLER_21_151 ();
 sg13g2_decap_4 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_fill_1 FILLER_21_203 ();
 sg13g2_fill_2 FILLER_21_209 ();
 sg13g2_decap_4 FILLER_21_215 ();
 sg13g2_fill_1 FILLER_21_228 ();
 sg13g2_fill_2 FILLER_21_239 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_fill_1 FILLER_21_252 ();
 sg13g2_fill_2 FILLER_21_257 ();
 sg13g2_fill_1 FILLER_21_314 ();
 sg13g2_fill_2 FILLER_21_346 ();
 sg13g2_decap_4 FILLER_21_363 ();
 sg13g2_fill_2 FILLER_21_380 ();
 sg13g2_fill_1 FILLER_21_382 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_4 FILLER_22_21 ();
 sg13g2_fill_2 FILLER_22_25 ();
 sg13g2_decap_8 FILLER_22_47 ();
 sg13g2_decap_4 FILLER_22_54 ();
 sg13g2_fill_2 FILLER_22_58 ();
 sg13g2_decap_4 FILLER_22_70 ();
 sg13g2_decap_4 FILLER_22_78 ();
 sg13g2_fill_2 FILLER_22_82 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_4 FILLER_22_98 ();
 sg13g2_fill_1 FILLER_22_102 ();
 sg13g2_decap_4 FILLER_22_125 ();
 sg13g2_fill_2 FILLER_22_129 ();
 sg13g2_decap_8 FILLER_22_145 ();
 sg13g2_fill_1 FILLER_22_152 ();
 sg13g2_decap_8 FILLER_22_165 ();
 sg13g2_decap_8 FILLER_22_172 ();
 sg13g2_decap_8 FILLER_22_192 ();
 sg13g2_decap_4 FILLER_22_199 ();
 sg13g2_fill_2 FILLER_22_207 ();
 sg13g2_fill_1 FILLER_22_209 ();
 sg13g2_fill_1 FILLER_22_214 ();
 sg13g2_fill_2 FILLER_22_224 ();
 sg13g2_decap_4 FILLER_22_236 ();
 sg13g2_fill_2 FILLER_22_240 ();
 sg13g2_fill_2 FILLER_22_252 ();
 sg13g2_fill_1 FILLER_22_254 ();
 sg13g2_decap_4 FILLER_22_264 ();
 sg13g2_fill_2 FILLER_22_268 ();
 sg13g2_fill_1 FILLER_22_275 ();
 sg13g2_decap_4 FILLER_22_310 ();
 sg13g2_fill_1 FILLER_22_314 ();
 sg13g2_fill_1 FILLER_22_332 ();
 sg13g2_fill_1 FILLER_22_343 ();
 sg13g2_fill_2 FILLER_22_373 ();
 sg13g2_decap_4 FILLER_22_380 ();
 sg13g2_fill_1 FILLER_22_384 ();
 sg13g2_decap_8 FILLER_22_398 ();
 sg13g2_decap_4 FILLER_22_405 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_fill_1 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_45 ();
 sg13g2_fill_2 FILLER_23_52 ();
 sg13g2_fill_1 FILLER_23_54 ();
 sg13g2_fill_1 FILLER_23_78 ();
 sg13g2_decap_8 FILLER_23_94 ();
 sg13g2_decap_4 FILLER_23_101 ();
 sg13g2_fill_2 FILLER_23_105 ();
 sg13g2_fill_2 FILLER_23_111 ();
 sg13g2_decap_8 FILLER_23_118 ();
 sg13g2_decap_4 FILLER_23_125 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_fill_2 FILLER_23_154 ();
 sg13g2_fill_1 FILLER_23_156 ();
 sg13g2_decap_4 FILLER_23_161 ();
 sg13g2_fill_1 FILLER_23_168 ();
 sg13g2_decap_4 FILLER_23_231 ();
 sg13g2_fill_2 FILLER_23_235 ();
 sg13g2_fill_2 FILLER_23_268 ();
 sg13g2_decap_8 FILLER_23_302 ();
 sg13g2_decap_8 FILLER_23_309 ();
 sg13g2_fill_2 FILLER_23_325 ();
 sg13g2_fill_1 FILLER_23_345 ();
 sg13g2_fill_2 FILLER_23_380 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_4 FILLER_24_28 ();
 sg13g2_decap_4 FILLER_24_47 ();
 sg13g2_fill_2 FILLER_24_51 ();
 sg13g2_decap_8 FILLER_24_67 ();
 sg13g2_decap_8 FILLER_24_74 ();
 sg13g2_fill_1 FILLER_24_81 ();
 sg13g2_decap_4 FILLER_24_105 ();
 sg13g2_fill_2 FILLER_24_109 ();
 sg13g2_fill_2 FILLER_24_129 ();
 sg13g2_fill_1 FILLER_24_131 ();
 sg13g2_fill_1 FILLER_24_135 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_fill_1 FILLER_24_147 ();
 sg13g2_fill_1 FILLER_24_188 ();
 sg13g2_decap_8 FILLER_24_194 ();
 sg13g2_decap_8 FILLER_24_201 ();
 sg13g2_fill_2 FILLER_24_208 ();
 sg13g2_fill_1 FILLER_24_210 ();
 sg13g2_decap_4 FILLER_24_216 ();
 sg13g2_fill_2 FILLER_24_220 ();
 sg13g2_decap_8 FILLER_24_235 ();
 sg13g2_decap_8 FILLER_24_251 ();
 sg13g2_decap_4 FILLER_24_258 ();
 sg13g2_fill_1 FILLER_24_271 ();
 sg13g2_decap_4 FILLER_24_275 ();
 sg13g2_fill_1 FILLER_24_279 ();
 sg13g2_decap_4 FILLER_24_284 ();
 sg13g2_fill_2 FILLER_24_291 ();
 sg13g2_fill_2 FILLER_24_306 ();
 sg13g2_decap_4 FILLER_24_370 ();
 sg13g2_decap_8 FILLER_24_379 ();
 sg13g2_decap_8 FILLER_24_386 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_4 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_44 ();
 sg13g2_decap_4 FILLER_25_51 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_4 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_99 ();
 sg13g2_decap_8 FILLER_25_106 ();
 sg13g2_decap_8 FILLER_25_121 ();
 sg13g2_decap_8 FILLER_25_143 ();
 sg13g2_decap_8 FILLER_25_150 ();
 sg13g2_fill_2 FILLER_25_157 ();
 sg13g2_fill_2 FILLER_25_163 ();
 sg13g2_fill_1 FILLER_25_165 ();
 sg13g2_fill_2 FILLER_25_175 ();
 sg13g2_fill_1 FILLER_25_177 ();
 sg13g2_fill_2 FILLER_25_192 ();
 sg13g2_fill_2 FILLER_25_199 ();
 sg13g2_decap_4 FILLER_25_237 ();
 sg13g2_fill_2 FILLER_25_249 ();
 sg13g2_decap_4 FILLER_25_287 ();
 sg13g2_fill_1 FILLER_25_291 ();
 sg13g2_decap_8 FILLER_25_306 ();
 sg13g2_fill_2 FILLER_25_313 ();
 sg13g2_fill_1 FILLER_25_315 ();
 sg13g2_decap_8 FILLER_25_321 ();
 sg13g2_decap_4 FILLER_25_332 ();
 sg13g2_fill_1 FILLER_25_336 ();
 sg13g2_fill_1 FILLER_25_347 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_fill_1 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_33 ();
 sg13g2_fill_1 FILLER_26_40 ();
 sg13g2_fill_2 FILLER_26_67 ();
 sg13g2_fill_1 FILLER_26_73 ();
 sg13g2_fill_2 FILLER_26_82 ();
 sg13g2_fill_1 FILLER_26_84 ();
 sg13g2_decap_4 FILLER_26_89 ();
 sg13g2_fill_2 FILLER_26_122 ();
 sg13g2_fill_1 FILLER_26_143 ();
 sg13g2_decap_4 FILLER_26_149 ();
 sg13g2_fill_1 FILLER_26_153 ();
 sg13g2_decap_8 FILLER_26_167 ();
 sg13g2_fill_1 FILLER_26_174 ();
 sg13g2_decap_4 FILLER_26_201 ();
 sg13g2_decap_8 FILLER_26_222 ();
 sg13g2_decap_4 FILLER_26_229 ();
 sg13g2_fill_1 FILLER_26_233 ();
 sg13g2_decap_8 FILLER_26_278 ();
 sg13g2_fill_2 FILLER_26_285 ();
 sg13g2_fill_1 FILLER_26_287 ();
 sg13g2_decap_4 FILLER_26_314 ();
 sg13g2_fill_2 FILLER_26_318 ();
 sg13g2_decap_4 FILLER_26_343 ();
 sg13g2_fill_1 FILLER_26_347 ();
 sg13g2_decap_4 FILLER_26_389 ();
 sg13g2_fill_1 FILLER_26_393 ();
 sg13g2_fill_2 FILLER_26_398 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_fill_2 FILLER_27_49 ();
 sg13g2_fill_1 FILLER_27_64 ();
 sg13g2_fill_2 FILLER_27_79 ();
 sg13g2_fill_1 FILLER_27_91 ();
 sg13g2_fill_1 FILLER_27_101 ();
 sg13g2_decap_8 FILLER_27_115 ();
 sg13g2_decap_8 FILLER_27_122 ();
 sg13g2_fill_2 FILLER_27_129 ();
 sg13g2_fill_1 FILLER_27_136 ();
 sg13g2_fill_1 FILLER_27_147 ();
 sg13g2_decap_4 FILLER_27_170 ();
 sg13g2_fill_2 FILLER_27_174 ();
 sg13g2_fill_2 FILLER_27_184 ();
 sg13g2_decap_8 FILLER_27_190 ();
 sg13g2_fill_2 FILLER_27_197 ();
 sg13g2_fill_1 FILLER_27_199 ();
 sg13g2_decap_8 FILLER_27_205 ();
 sg13g2_decap_8 FILLER_27_212 ();
 sg13g2_fill_2 FILLER_27_219 ();
 sg13g2_decap_8 FILLER_27_230 ();
 sg13g2_decap_8 FILLER_27_237 ();
 sg13g2_decap_8 FILLER_27_251 ();
 sg13g2_decap_4 FILLER_27_258 ();
 sg13g2_decap_4 FILLER_27_293 ();
 sg13g2_fill_1 FILLER_27_297 ();
 sg13g2_decap_4 FILLER_27_303 ();
 sg13g2_fill_2 FILLER_27_351 ();
 sg13g2_fill_1 FILLER_27_353 ();
 sg13g2_decap_8 FILLER_27_357 ();
 sg13g2_fill_1 FILLER_27_364 ();
 sg13g2_decap_4 FILLER_27_404 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_4 FILLER_28_35 ();
 sg13g2_fill_1 FILLER_28_39 ();
 sg13g2_decap_8 FILLER_28_66 ();
 sg13g2_decap_8 FILLER_28_86 ();
 sg13g2_decap_4 FILLER_28_93 ();
 sg13g2_fill_1 FILLER_28_97 ();
 sg13g2_decap_4 FILLER_28_102 ();
 sg13g2_fill_1 FILLER_28_106 ();
 sg13g2_decap_8 FILLER_28_124 ();
 sg13g2_fill_1 FILLER_28_131 ();
 sg13g2_fill_1 FILLER_28_136 ();
 sg13g2_decap_8 FILLER_28_141 ();
 sg13g2_decap_4 FILLER_28_148 ();
 sg13g2_fill_2 FILLER_28_152 ();
 sg13g2_decap_8 FILLER_28_159 ();
 sg13g2_fill_2 FILLER_28_166 ();
 sg13g2_fill_2 FILLER_28_191 ();
 sg13g2_fill_2 FILLER_28_237 ();
 sg13g2_fill_1 FILLER_28_239 ();
 sg13g2_decap_8 FILLER_28_252 ();
 sg13g2_decap_4 FILLER_28_259 ();
 sg13g2_decap_4 FILLER_28_268 ();
 sg13g2_fill_1 FILLER_28_272 ();
 sg13g2_fill_2 FILLER_28_280 ();
 sg13g2_decap_4 FILLER_28_317 ();
 sg13g2_decap_8 FILLER_28_326 ();
 sg13g2_fill_2 FILLER_28_333 ();
 sg13g2_fill_1 FILLER_28_335 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_fill_2 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_55 ();
 sg13g2_decap_8 FILLER_29_62 ();
 sg13g2_fill_2 FILLER_29_69 ();
 sg13g2_fill_1 FILLER_29_71 ();
 sg13g2_fill_2 FILLER_29_130 ();
 sg13g2_fill_1 FILLER_29_132 ();
 sg13g2_decap_4 FILLER_29_155 ();
 sg13g2_fill_2 FILLER_29_159 ();
 sg13g2_decap_8 FILLER_29_164 ();
 sg13g2_decap_8 FILLER_29_192 ();
 sg13g2_decap_8 FILLER_29_208 ();
 sg13g2_decap_4 FILLER_29_215 ();
 sg13g2_fill_2 FILLER_29_219 ();
 sg13g2_decap_8 FILLER_29_229 ();
 sg13g2_fill_2 FILLER_29_236 ();
 sg13g2_fill_2 FILLER_29_251 ();
 sg13g2_fill_1 FILLER_29_265 ();
 sg13g2_decap_4 FILLER_29_280 ();
 sg13g2_fill_2 FILLER_29_284 ();
 sg13g2_fill_2 FILLER_29_291 ();
 sg13g2_fill_1 FILLER_29_293 ();
 sg13g2_fill_2 FILLER_29_312 ();
 sg13g2_fill_2 FILLER_29_345 ();
 sg13g2_decap_8 FILLER_29_396 ();
 sg13g2_decap_4 FILLER_29_403 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_4 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_85 ();
 sg13g2_fill_2 FILLER_30_92 ();
 sg13g2_decap_4 FILLER_30_98 ();
 sg13g2_fill_2 FILLER_30_102 ();
 sg13g2_fill_2 FILLER_30_108 ();
 sg13g2_fill_1 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_125 ();
 sg13g2_decap_8 FILLER_30_132 ();
 sg13g2_decap_8 FILLER_30_139 ();
 sg13g2_decap_4 FILLER_30_160 ();
 sg13g2_fill_1 FILLER_30_164 ();
 sg13g2_fill_1 FILLER_30_192 ();
 sg13g2_decap_8 FILLER_30_198 ();
 sg13g2_decap_8 FILLER_30_205 ();
 sg13g2_fill_2 FILLER_30_216 ();
 sg13g2_fill_1 FILLER_30_218 ();
 sg13g2_fill_1 FILLER_30_224 ();
 sg13g2_decap_4 FILLER_30_234 ();
 sg13g2_decap_8 FILLER_30_247 ();
 sg13g2_fill_2 FILLER_30_254 ();
 sg13g2_fill_1 FILLER_30_256 ();
 sg13g2_decap_8 FILLER_30_273 ();
 sg13g2_decap_8 FILLER_30_280 ();
 sg13g2_decap_4 FILLER_30_287 ();
 sg13g2_decap_8 FILLER_30_319 ();
 sg13g2_fill_1 FILLER_30_347 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_fill_1 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_61 ();
 sg13g2_decap_4 FILLER_31_68 ();
 sg13g2_fill_2 FILLER_31_72 ();
 sg13g2_fill_1 FILLER_31_86 ();
 sg13g2_fill_1 FILLER_31_97 ();
 sg13g2_fill_1 FILLER_31_125 ();
 sg13g2_decap_8 FILLER_31_131 ();
 sg13g2_fill_2 FILLER_31_138 ();
 sg13g2_fill_2 FILLER_31_148 ();
 sg13g2_fill_1 FILLER_31_150 ();
 sg13g2_fill_2 FILLER_31_159 ();
 sg13g2_decap_4 FILLER_31_201 ();
 sg13g2_decap_8 FILLER_31_219 ();
 sg13g2_decap_4 FILLER_31_226 ();
 sg13g2_fill_2 FILLER_31_230 ();
 sg13g2_decap_4 FILLER_31_240 ();
 sg13g2_decap_8 FILLER_31_255 ();
 sg13g2_decap_8 FILLER_31_262 ();
 sg13g2_decap_8 FILLER_31_269 ();
 sg13g2_decap_8 FILLER_31_276 ();
 sg13g2_decap_8 FILLER_31_283 ();
 sg13g2_decap_8 FILLER_31_316 ();
 sg13g2_fill_2 FILLER_31_357 ();
 sg13g2_fill_1 FILLER_31_359 ();
 sg13g2_fill_2 FILLER_31_365 ();
 sg13g2_fill_2 FILLER_31_391 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_4 FILLER_32_84 ();
 sg13g2_decap_4 FILLER_32_114 ();
 sg13g2_fill_2 FILLER_32_118 ();
 sg13g2_decap_8 FILLER_32_125 ();
 sg13g2_decap_8 FILLER_32_139 ();
 sg13g2_fill_1 FILLER_32_146 ();
 sg13g2_decap_8 FILLER_32_151 ();
 sg13g2_fill_1 FILLER_32_158 ();
 sg13g2_decap_4 FILLER_32_164 ();
 sg13g2_decap_8 FILLER_32_198 ();
 sg13g2_fill_2 FILLER_32_205 ();
 sg13g2_fill_1 FILLER_32_207 ();
 sg13g2_fill_2 FILLER_32_236 ();
 sg13g2_fill_1 FILLER_32_238 ();
 sg13g2_decap_8 FILLER_32_246 ();
 sg13g2_fill_2 FILLER_32_253 ();
 sg13g2_decap_4 FILLER_32_272 ();
 sg13g2_decap_4 FILLER_32_296 ();
 sg13g2_fill_1 FILLER_32_300 ();
 sg13g2_decap_4 FILLER_32_314 ();
 sg13g2_fill_2 FILLER_32_318 ();
 sg13g2_decap_8 FILLER_32_324 ();
 sg13g2_decap_8 FILLER_32_331 ();
 sg13g2_fill_1 FILLER_32_351 ();
 sg13g2_fill_1 FILLER_32_364 ();
 sg13g2_fill_1 FILLER_32_369 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_4 FILLER_33_96 ();
 sg13g2_decap_4 FILLER_33_104 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_4 FILLER_33_131 ();
 sg13g2_fill_1 FILLER_33_135 ();
 sg13g2_decap_8 FILLER_33_172 ();
 sg13g2_fill_2 FILLER_33_183 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_decap_4 FILLER_33_203 ();
 sg13g2_fill_1 FILLER_33_207 ();
 sg13g2_decap_8 FILLER_33_242 ();
 sg13g2_decap_4 FILLER_33_249 ();
 sg13g2_fill_2 FILLER_33_275 ();
 sg13g2_decap_4 FILLER_33_294 ();
 sg13g2_fill_1 FILLER_33_298 ();
 sg13g2_decap_8 FILLER_33_303 ();
 sg13g2_decap_4 FILLER_33_310 ();
 sg13g2_decap_4 FILLER_33_336 ();
 sg13g2_fill_1 FILLER_33_340 ();
 sg13g2_decap_8 FILLER_33_353 ();
 sg13g2_fill_2 FILLER_33_360 ();
 sg13g2_fill_1 FILLER_33_371 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_4 FILLER_34_63 ();
 sg13g2_fill_1 FILLER_34_67 ();
 sg13g2_fill_2 FILLER_34_94 ();
 sg13g2_fill_1 FILLER_34_96 ();
 sg13g2_decap_8 FILLER_34_137 ();
 sg13g2_fill_1 FILLER_34_144 ();
 sg13g2_decap_8 FILLER_34_153 ();
 sg13g2_decap_4 FILLER_34_160 ();
 sg13g2_fill_2 FILLER_34_186 ();
 sg13g2_fill_1 FILLER_34_188 ();
 sg13g2_fill_2 FILLER_34_205 ();
 sg13g2_fill_1 FILLER_34_207 ();
 sg13g2_fill_2 FILLER_34_221 ();
 sg13g2_fill_1 FILLER_34_223 ();
 sg13g2_fill_2 FILLER_34_229 ();
 sg13g2_fill_1 FILLER_34_231 ();
 sg13g2_fill_2 FILLER_34_237 ();
 sg13g2_decap_8 FILLER_34_247 ();
 sg13g2_fill_2 FILLER_34_254 ();
 sg13g2_decap_8 FILLER_34_272 ();
 sg13g2_decap_4 FILLER_34_279 ();
 sg13g2_decap_4 FILLER_34_287 ();
 sg13g2_fill_1 FILLER_34_291 ();
 sg13g2_decap_8 FILLER_34_306 ();
 sg13g2_decap_4 FILLER_34_313 ();
 sg13g2_fill_2 FILLER_34_317 ();
 sg13g2_fill_1 FILLER_34_331 ();
 sg13g2_fill_2 FILLER_34_336 ();
 sg13g2_decap_8 FILLER_34_355 ();
 sg13g2_fill_2 FILLER_34_362 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_fill_2 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_83 ();
 sg13g2_decap_8 FILLER_35_90 ();
 sg13g2_decap_8 FILLER_35_97 ();
 sg13g2_decap_4 FILLER_35_104 ();
 sg13g2_decap_4 FILLER_35_116 ();
 sg13g2_fill_1 FILLER_35_145 ();
 sg13g2_fill_2 FILLER_35_159 ();
 sg13g2_fill_1 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_4 FILLER_35_189 ();
 sg13g2_fill_2 FILLER_35_193 ();
 sg13g2_fill_1 FILLER_35_221 ();
 sg13g2_fill_2 FILLER_35_230 ();
 sg13g2_fill_1 FILLER_35_232 ();
 sg13g2_decap_8 FILLER_35_253 ();
 sg13g2_fill_1 FILLER_35_260 ();
 sg13g2_decap_4 FILLER_35_278 ();
 sg13g2_fill_2 FILLER_35_282 ();
 sg13g2_decap_8 FILLER_35_305 ();
 sg13g2_decap_4 FILLER_35_312 ();
 sg13g2_fill_1 FILLER_35_316 ();
 sg13g2_decap_8 FILLER_35_333 ();
 sg13g2_decap_4 FILLER_35_340 ();
 sg13g2_fill_2 FILLER_35_360 ();
 sg13g2_fill_2 FILLER_35_366 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_4 FILLER_36_98 ();
 sg13g2_decap_4 FILLER_36_128 ();
 sg13g2_fill_2 FILLER_36_132 ();
 sg13g2_decap_8 FILLER_36_149 ();
 sg13g2_decap_8 FILLER_36_156 ();
 sg13g2_decap_4 FILLER_36_163 ();
 sg13g2_fill_1 FILLER_36_167 ();
 sg13g2_decap_8 FILLER_36_181 ();
 sg13g2_decap_8 FILLER_36_201 ();
 sg13g2_fill_2 FILLER_36_217 ();
 sg13g2_decap_8 FILLER_36_235 ();
 sg13g2_fill_2 FILLER_36_242 ();
 sg13g2_decap_8 FILLER_36_249 ();
 sg13g2_decap_8 FILLER_36_256 ();
 sg13g2_decap_4 FILLER_36_263 ();
 sg13g2_fill_1 FILLER_36_267 ();
 sg13g2_decap_4 FILLER_36_280 ();
 sg13g2_fill_1 FILLER_36_284 ();
 sg13g2_decap_8 FILLER_36_305 ();
 sg13g2_decap_8 FILLER_36_312 ();
 sg13g2_fill_1 FILLER_36_319 ();
 sg13g2_decap_4 FILLER_36_336 ();
 sg13g2_fill_1 FILLER_36_340 ();
 sg13g2_fill_2 FILLER_36_349 ();
 sg13g2_fill_1 FILLER_36_351 ();
 sg13g2_fill_1 FILLER_36_365 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_4 FILLER_37_126 ();
 sg13g2_fill_1 FILLER_37_130 ();
 sg13g2_fill_1 FILLER_37_150 ();
 sg13g2_fill_1 FILLER_37_159 ();
 sg13g2_fill_2 FILLER_37_181 ();
 sg13g2_fill_2 FILLER_37_214 ();
 sg13g2_fill_1 FILLER_37_216 ();
 sg13g2_fill_1 FILLER_37_238 ();
 sg13g2_fill_2 FILLER_37_260 ();
 sg13g2_fill_1 FILLER_37_262 ();
 sg13g2_decap_8 FILLER_37_276 ();
 sg13g2_decap_4 FILLER_37_307 ();
 sg13g2_fill_1 FILLER_37_311 ();
 sg13g2_fill_2 FILLER_37_333 ();
 sg13g2_fill_2 FILLER_37_385 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_fill_2 FILLER_38_132 ();
 sg13g2_fill_2 FILLER_38_142 ();
 sg13g2_fill_1 FILLER_38_151 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_fill_1 FILLER_38_164 ();
 sg13g2_decap_8 FILLER_38_176 ();
 sg13g2_decap_4 FILLER_38_183 ();
 sg13g2_fill_1 FILLER_38_187 ();
 sg13g2_fill_2 FILLER_38_196 ();
 sg13g2_fill_1 FILLER_38_198 ();
 sg13g2_decap_8 FILLER_38_203 ();
 sg13g2_decap_8 FILLER_38_210 ();
 sg13g2_decap_8 FILLER_38_217 ();
 sg13g2_decap_8 FILLER_38_232 ();
 sg13g2_decap_8 FILLER_38_239 ();
 sg13g2_decap_8 FILLER_38_246 ();
 sg13g2_decap_8 FILLER_38_253 ();
 sg13g2_fill_2 FILLER_38_260 ();
 sg13g2_decap_8 FILLER_38_278 ();
 sg13g2_fill_1 FILLER_38_303 ();
 sg13g2_fill_2 FILLER_38_309 ();
 sg13g2_fill_1 FILLER_38_311 ();
 sg13g2_fill_2 FILLER_38_316 ();
 sg13g2_fill_1 FILLER_38_335 ();
 sg13g2_fill_2 FILLER_38_341 ();
 sg13g2_fill_1 FILLER_38_343 ();
 sg13g2_fill_2 FILLER_38_349 ();
 sg13g2_fill_1 FILLER_38_360 ();
 sg13g2_fill_2 FILLER_38_370 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net94;
 assign uio_oe[1] = net11;
 assign uio_oe[2] = net12;
 assign uio_oe[3] = net13;
 assign uio_oe[4] = net14;
 assign uio_oe[5] = net15;
 assign uio_oe[6] = net16;
 assign uio_oe[7] = net17;
 assign uio_out[1] = net18;
 assign uio_out[2] = net19;
 assign uio_out[3] = net20;
 assign uio_out[4] = net21;
 assign uio_out[5] = net22;
 assign uio_out[6] = net23;
 assign uio_out[7] = net24;
endmodule
