module tt_um_dpi_adexp (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire clknet_leaf_0_clk;
 wire \core.C_q[10] ;
 wire \core.C_q[11] ;
 wire \core.C_q[4] ;
 wire \core.C_q[5] ;
 wire \core.C_q[6] ;
 wire \core.C_q[7] ;
 wire \core.C_q[8] ;
 wire \core.C_q[9] ;
 wire \core.TauW_q[10] ;
 wire \core.TauW_q[11] ;
 wire \core.TauW_q[4] ;
 wire \core.TauW_q[5] ;
 wire \core.TauW_q[6] ;
 wire \core.TauW_q[7] ;
 wire \core.TauW_q[8] ;
 wire \core.TauW_q[9] ;
 wire \core.VT_q[10] ;
 wire \core.VT_q[11] ;
 wire \core.VT_q[4] ;
 wire \core.VT_q[5] ;
 wire \core.VT_q[6] ;
 wire \core.VT_q[7] ;
 wire \core.VT_q[8] ;
 wire \core.VT_q[9] ;
 wire \core.V[0] ;
 wire \core.V[10] ;
 wire \core.V[11] ;
 wire \core.V[12] ;
 wire \core.V[13] ;
 wire \core.V[14] ;
 wire \core.V[15] ;
 wire \core.V[1] ;
 wire \core.V[2] ;
 wire \core.V[3] ;
 wire \core.V[4] ;
 wire \core.V[5] ;
 wire \core.V[6] ;
 wire \core.V[7] ;
 wire \core.V[8] ;
 wire \core.V[9] ;
 wire \core.Vreset_q[10] ;
 wire \core.Vreset_q[11] ;
 wire \core.Vreset_q[4] ;
 wire \core.Vreset_q[5] ;
 wire \core.Vreset_q[6] ;
 wire \core.Vreset_q[7] ;
 wire \core.Vreset_q[8] ;
 wire \core.Vreset_q[9] ;
 wire \core.a_q[10] ;
 wire \core.a_q[11] ;
 wire \core.a_q[4] ;
 wire \core.a_q[5] ;
 wire \core.a_q[6] ;
 wire \core.a_q[7] ;
 wire \core.a_q[8] ;
 wire \core.a_q[9] ;
 wire \core.b_q[10] ;
 wire \core.b_q[11] ;
 wire \core.b_q[4] ;
 wire \core.b_q[5] ;
 wire \core.b_q[6] ;
 wire \core.b_q[7] ;
 wire \core.b_q[8] ;
 wire \core.b_q[9] ;
 wire \core.byte_acc[0] ;
 wire \core.byte_acc[1] ;
 wire \core.byte_acc[2] ;
 wire \core.byte_acc[3] ;
 wire \core.byte_acc[4] ;
 wire \core.byte_acc[5] ;
 wire \core.byte_acc[6] ;
 wire \core.byte_acc[7] ;
 wire \core.dV[0] ;
 wire \core.dV[10] ;
 wire \core.dV[11] ;
 wire \core.dV[12] ;
 wire \core.dV[13] ;
 wire \core.dV[14] ;
 wire \core.dV[15] ;
 wire \core.dV[1] ;
 wire \core.dV[2] ;
 wire \core.dV[3] ;
 wire \core.dV[4] ;
 wire \core.dV[5] ;
 wire \core.dV[6] ;
 wire \core.dV[7] ;
 wire \core.dV[8] ;
 wire \core.dV[9] ;
 wire \core.drive[0] ;
 wire \core.drive[1] ;
 wire \core.drive[2] ;
 wire \core.drive[3] ;
 wire \core.dw[0] ;
 wire \core.dw[10] ;
 wire \core.dw[11] ;
 wire \core.dw[12] ;
 wire \core.dw[13] ;
 wire \core.dw[14] ;
 wire \core.dw[15] ;
 wire \core.dw[1] ;
 wire \core.dw[2] ;
 wire \core.dw[3] ;
 wire \core.dw[4] ;
 wire \core.dw[5] ;
 wire \core.dw[6] ;
 wire \core.dw[7] ;
 wire \core.dw[8] ;
 wire \core.dw[9] ;
 wire \core.leak[10] ;
 wire \core.leak[1] ;
 wire \core.leak[2] ;
 wire \core.load_prev ;
 wire \core.lstate[0] ;
 wire \core.lstate[1] ;
 wire \core.lstate[2] ;
 wire \core.nibble_cnt ;
 wire \core.p_C[0] ;
 wire \core.p_C[1] ;
 wire \core.p_C[2] ;
 wire \core.p_C[3] ;
 wire \core.p_C[4] ;
 wire \core.p_C[5] ;
 wire \core.p_C[6] ;
 wire \core.p_C[7] ;
 wire \core.p_TauW[0] ;
 wire \core.p_TauW[1] ;
 wire \core.p_TauW[2] ;
 wire \core.p_TauW[3] ;
 wire \core.p_TauW[4] ;
 wire \core.p_TauW[5] ;
 wire \core.p_TauW[6] ;
 wire \core.p_TauW[7] ;
 wire \core.p_VT[0] ;
 wire \core.p_VT[1] ;
 wire \core.p_VT[2] ;
 wire \core.p_VT[3] ;
 wire \core.p_VT[4] ;
 wire \core.p_VT[5] ;
 wire \core.p_VT[6] ;
 wire \core.p_VT[7] ;
 wire \core.p_Vreset[0] ;
 wire \core.p_Vreset[1] ;
 wire \core.p_Vreset[2] ;
 wire \core.p_Vreset[3] ;
 wire \core.p_Vreset[4] ;
 wire \core.p_Vreset[5] ;
 wire \core.p_Vreset[6] ;
 wire \core.p_Vreset[7] ;
 wire \core.p_a[0] ;
 wire \core.p_a[1] ;
 wire \core.p_a[2] ;
 wire \core.p_a[3] ;
 wire \core.p_a[4] ;
 wire \core.p_a[5] ;
 wire \core.p_a[6] ;
 wire \core.p_a[7] ;
 wire \core.p_b[0] ;
 wire \core.p_b[1] ;
 wire \core.p_b[2] ;
 wire \core.p_b[3] ;
 wire \core.p_b[4] ;
 wire \core.p_b[5] ;
 wire \core.p_b[6] ;
 wire \core.p_b[7] ;
 wire \core.param_idx[0] ;
 wire \core.param_idx[1] ;
 wire \core.param_idx[2] ;
 wire \core.param_idx[3] ;
 wire \core.params_ready ;
 wire \core.s_C[0] ;
 wire \core.s_C[1] ;
 wire \core.s_C[2] ;
 wire \core.s_C[3] ;
 wire \core.s_C[4] ;
 wire \core.s_C[5] ;
 wire \core.s_C[6] ;
 wire \core.s_C[7] ;
 wire \core.s_TauW[0] ;
 wire \core.s_TauW[1] ;
 wire \core.s_TauW[2] ;
 wire \core.s_TauW[3] ;
 wire \core.s_TauW[4] ;
 wire \core.s_TauW[5] ;
 wire \core.s_TauW[6] ;
 wire \core.s_TauW[7] ;
 wire \core.s_VT[0] ;
 wire \core.s_VT[1] ;
 wire \core.s_VT[2] ;
 wire \core.s_VT[3] ;
 wire \core.s_VT[4] ;
 wire \core.s_VT[5] ;
 wire \core.s_VT[6] ;
 wire \core.s_VT[7] ;
 wire \core.s_Vreset[0] ;
 wire \core.s_Vreset[1] ;
 wire \core.s_Vreset[2] ;
 wire \core.s_Vreset[3] ;
 wire \core.s_Vreset[4] ;
 wire \core.s_Vreset[5] ;
 wire \core.s_Vreset[6] ;
 wire \core.s_Vreset[7] ;
 wire \core.s_a[0] ;
 wire \core.s_a[1] ;
 wire \core.s_a[2] ;
 wire \core.s_a[3] ;
 wire \core.s_a[4] ;
 wire \core.s_a[5] ;
 wire \core.s_a[6] ;
 wire \core.s_a[7] ;
 wire \core.s_b[0] ;
 wire \core.s_b[1] ;
 wire \core.s_b[2] ;
 wire \core.s_b[3] ;
 wire \core.s_b[4] ;
 wire \core.s_b[5] ;
 wire \core.s_b[6] ;
 wire \core.s_b[7] ;
 wire \core.spike_reg ;
 wire \core.vm8_reg[2] ;
 wire \core.vm8_reg[3] ;
 wire \core.vm8_reg[7] ;
 wire \core.w8_reg[2] ;
 wire \core.w8_reg[3] ;
 wire \core.w8_reg[7] ;
 wire \core.w[0] ;
 wire \core.w[10] ;
 wire \core.w[11] ;
 wire \core.w[12] ;
 wire \core.w[13] ;
 wire \core.w[14] ;
 wire \core.w[15] ;
 wire \core.w[1] ;
 wire \core.w[2] ;
 wire \core.w[3] ;
 wire \core.w[4] ;
 wire \core.w[5] ;
 wire \core.w[6] ;
 wire \core.w[7] ;
 wire \core.w[8] ;
 wire \core.w[9] ;
 wire \core.watchdog_cnt[0] ;
 wire \core.watchdog_cnt[10] ;
 wire \core.watchdog_cnt[11] ;
 wire \core.watchdog_cnt[12] ;
 wire \core.watchdog_cnt[13] ;
 wire \core.watchdog_cnt[14] ;
 wire \core.watchdog_cnt[15] ;
 wire \core.watchdog_cnt[1] ;
 wire \core.watchdog_cnt[2] ;
 wire \core.watchdog_cnt[3] ;
 wire \core.watchdog_cnt[4] ;
 wire \core.watchdog_cnt[5] ;
 wire \core.watchdog_cnt[6] ;
 wire \core.watchdog_cnt[7] ;
 wire \core.watchdog_cnt[8] ;
 wire \core.watchdog_cnt[9] ;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_35_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;

 sg13g2_inv_4 _2736_ (.A(net562),
    .Y(_1851_));
 sg13g2_inv_1 _2737_ (.Y(_1852_),
    .A(net365));
 sg13g2_inv_2 _2738_ (.Y(_1853_),
    .A(net557));
 sg13g2_inv_1 _2739_ (.Y(_1854_),
    .A(net371));
 sg13g2_inv_2 _2740_ (.Y(_1855_),
    .A(net577));
 sg13g2_inv_4 _2741_ (.A(net545),
    .Y(_1856_));
 sg13g2_inv_4 _2742_ (.A(net575),
    .Y(_1857_));
 sg13g2_inv_4 _2743_ (.A(net570),
    .Y(_1858_));
 sg13g2_inv_1 _2744_ (.Y(_1859_),
    .A(net378));
 sg13g2_inv_4 _2745_ (.A(net568),
    .Y(_1860_));
 sg13g2_inv_4 _2746_ (.A(net548),
    .Y(_1861_));
 sg13g2_inv_1 _2747_ (.Y(_1862_),
    .A(net392));
 sg13g2_inv_1 _2748_ (.Y(_1863_),
    .A(net390));
 sg13g2_inv_1 _2749_ (.Y(_1864_),
    .A(net376));
 sg13g2_inv_1 _2750_ (.Y(_1865_),
    .A(net496));
 sg13g2_inv_1 _2751_ (.Y(_1866_),
    .A(net425));
 sg13g2_inv_1 _2752_ (.Y(_1867_),
    .A(net363));
 sg13g2_inv_1 _2753_ (.Y(_1868_),
    .A(net403));
 sg13g2_inv_1 _2754_ (.Y(_1869_),
    .A(net352));
 sg13g2_inv_1 _2755_ (.Y(_1870_),
    .A(net355));
 sg13g2_inv_1 _2756_ (.Y(_1871_),
    .A(net380));
 sg13g2_inv_1 _2757_ (.Y(_1872_),
    .A(net353));
 sg13g2_inv_1 _2758_ (.Y(_1873_),
    .A(net367));
 sg13g2_inv_1 _2759_ (.Y(_1874_),
    .A(net357));
 sg13g2_inv_1 _2760_ (.Y(_1875_),
    .A(net386));
 sg13g2_inv_1 _2761_ (.Y(_1876_),
    .A(net398));
 sg13g2_inv_1 _2762_ (.Y(_1877_),
    .A(net396));
 sg13g2_inv_1 _2763_ (.Y(_1878_),
    .A(net415));
 sg13g2_inv_1 _2764_ (.Y(_1879_),
    .A(net373));
 sg13g2_inv_1 _2765_ (.Y(_1880_),
    .A(net427));
 sg13g2_inv_1 _2766_ (.Y(_1881_),
    .A(net434));
 sg13g2_inv_1 _2767_ (.Y(_1882_),
    .A(net445));
 sg13g2_inv_1 _2768_ (.Y(_1883_),
    .A(net535));
 sg13g2_inv_1 _2769_ (.Y(_1884_),
    .A(net456));
 sg13g2_inv_1 _2770_ (.Y(_1885_),
    .A(net484));
 sg13g2_inv_1 _2771_ (.Y(_1886_),
    .A(net423));
 sg13g2_inv_1 _2772_ (.Y(_1887_),
    .A(net451));
 sg13g2_inv_1 _2773_ (.Y(_1888_),
    .A(net409));
 sg13g2_inv_1 _2774_ (.Y(_1889_),
    .A(net599));
 sg13g2_inv_1 _2775_ (.Y(_1890_),
    .A(net429));
 sg13g2_inv_1 _2776_ (.Y(_1891_),
    .A(net448));
 sg13g2_inv_1 _2777_ (.Y(_1892_),
    .A(net529));
 sg13g2_inv_1 _2778_ (.Y(_1893_),
    .A(net349));
 sg13g2_inv_1 _2779_ (.Y(_1894_),
    .A(net384));
 sg13g2_inv_1 _2780_ (.Y(_1895_),
    .A(net361));
 sg13g2_inv_1 _2781_ (.Y(_1896_),
    .A(net359));
 sg13g2_inv_1 _2782_ (.Y(_1897_),
    .A(net419));
 sg13g2_inv_1 _2783_ (.Y(_1898_),
    .A(net404));
 sg13g2_inv_1 _2784_ (.Y(_1899_),
    .A(net481));
 sg13g2_inv_1 _2785_ (.Y(_1900_),
    .A(net537));
 sg13g2_inv_1 _2786_ (.Y(_1901_),
    .A(net442));
 sg13g2_inv_1 _2787_ (.Y(_1902_),
    .A(net432));
 sg13g2_inv_1 _2788_ (.Y(_1903_),
    .A(net470));
 sg13g2_inv_1 _2789_ (.Y(_1904_),
    .A(net501));
 sg13g2_inv_1 _2790_ (.Y(_1905_),
    .A(net487));
 sg13g2_inv_1 _2791_ (.Y(_1906_),
    .A(net388));
 sg13g2_inv_1 _2792_ (.Y(_1907_),
    .A(net351));
 sg13g2_inv_1 _2793_ (.Y(_1908_),
    .A(\core.p_a[6] ));
 sg13g2_inv_1 _2794_ (.Y(_1909_),
    .A(net837));
 sg13g2_inv_1 _2795_ (.Y(_1910_),
    .A(net828));
 sg13g2_inv_1 _2796_ (.Y(_1911_),
    .A(net508));
 sg13g2_inv_1 _2797_ (.Y(_1912_),
    .A(net465));
 sg13g2_inv_1 _2798_ (.Y(_1913_),
    .A(net394));
 sg13g2_inv_1 _2799_ (.Y(_1914_),
    .A(net611));
 sg13g2_inv_1 _2800_ (.Y(_1915_),
    .A(net463));
 sg13g2_inv_1 _2801_ (.Y(_1916_),
    .A(net436));
 sg13g2_inv_1 _2802_ (.Y(_1917_),
    .A(net369));
 sg13g2_inv_1 _2803_ (.Y(_1918_),
    .A(net584));
 sg13g2_inv_1 _2804_ (.Y(_1919_),
    .A(net878));
 sg13g2_inv_1 _2805_ (.Y(_1920_),
    .A(\core.w[2] ));
 sg13g2_inv_2 _2806_ (.Y(_1921_),
    .A(net2));
 sg13g2_inv_1 _2807_ (.Y(_1922_),
    .A(\core.V[9] ));
 sg13g2_inv_1 _2808_ (.Y(_1923_),
    .A(\core.V[8] ));
 sg13g2_inv_1 _2809_ (.Y(_1924_),
    .A(net719));
 sg13g2_inv_2 _2810_ (.Y(_1925_),
    .A(\core.TauW_q[11] ));
 sg13g2_inv_4 _2811_ (.A(\core.TauW_q[10] ),
    .Y(_1926_));
 sg13g2_inv_4 _2812_ (.A(\core.TauW_q[9] ),
    .Y(_1927_));
 sg13g2_inv_2 _2813_ (.Y(_1928_),
    .A(net731));
 sg13g2_inv_1 _2814_ (.Y(_1929_),
    .A(net732));
 sg13g2_inv_1 _2815_ (.Y(_1930_),
    .A(\core.TauW_q[5] ));
 sg13g2_inv_1 _2816_ (.Y(_1931_),
    .A(net737));
 sg13g2_inv_1 _2817_ (.Y(_1932_),
    .A(net747));
 sg13g2_inv_1 _2818_ (.Y(_1933_),
    .A(net573));
 sg13g2_inv_1 _2819_ (.Y(_1934_),
    .A(net597));
 sg13g2_inv_1 _2820_ (.Y(_1935_),
    .A(\core.Vreset_q[11] ));
 sg13g2_inv_1 _2821_ (.Y(_1936_),
    .A(net512));
 sg13g2_inv_1 _2822_ (.Y(_1937_),
    .A(\core.Vreset_q[8] ));
 sg13g2_inv_1 _2823_ (.Y(_1938_),
    .A(net533));
 sg13g2_inv_1 _2824_ (.Y(_1939_),
    .A(\core.Vreset_q[6] ));
 sg13g2_inv_1 _2825_ (.Y(_1940_),
    .A(net490));
 sg13g2_inv_1 _2826_ (.Y(_1941_),
    .A(net492));
 sg13g2_inv_1 _2827_ (.Y(_1942_),
    .A(\core.VT_q[11] ));
 sg13g2_inv_2 _2828_ (.Y(_1943_),
    .A(net482));
 sg13g2_inv_1 _2829_ (.Y(_1944_),
    .A(\core.VT_q[8] ));
 sg13g2_inv_1 _2830_ (.Y(_1945_),
    .A(net531));
 sg13g2_inv_1 _2831_ (.Y(_1946_),
    .A(net494));
 sg13g2_inv_1 _2832_ (.Y(_1947_),
    .A(net515));
 sg13g2_inv_1 _2833_ (.Y(_1948_),
    .A(\core.VT_q[4] ));
 sg13g2_inv_2 _2834_ (.Y(_1949_),
    .A(net826));
 sg13g2_inv_2 _2835_ (.Y(_1950_),
    .A(net341));
 sg13g2_inv_2 _2836_ (.Y(_1951_),
    .A(\core.C_q[9] ));
 sg13g2_inv_2 _2837_ (.Y(_1952_),
    .A(\core.C_q[8] ));
 sg13g2_inv_4 _2838_ (.A(\core.C_q[7] ),
    .Y(_1953_));
 sg13g2_inv_2 _2839_ (.Y(_1954_),
    .A(\core.C_q[6] ));
 sg13g2_inv_2 _2840_ (.Y(_1955_),
    .A(net758));
 sg13g2_inv_1 _2841_ (.Y(_1956_),
    .A(\core.w[7] ));
 sg13g2_inv_1 _2842_ (.Y(_1957_),
    .A(net850));
 sg13g2_inv_4 _2843_ (.A(net810),
    .Y(_1958_));
 sg13g2_inv_1 _2844_ (.Y(_1959_),
    .A(\core.watchdog_cnt[14] ));
 sg13g2_inv_1 _2845_ (.Y(_1960_),
    .A(net477));
 sg13g2_inv_1 _2846_ (.Y(_1961_),
    .A(net853));
 sg13g2_inv_2 _2847_ (.Y(_1962_),
    .A(_0025_));
 sg13g2_inv_1 _2848_ (.Y(_1963_),
    .A(net757));
 sg13g2_inv_1 _2849_ (.Y(_1964_),
    .A(net753));
 sg13g2_inv_2 _2850_ (.Y(_1965_),
    .A(net752));
 sg13g2_inv_2 _2851_ (.Y(_1966_),
    .A(_0022_));
 sg13g2_inv_1 _2852_ (.Y(_1967_),
    .A(_0021_));
 sg13g2_inv_2 _2853_ (.Y(_1968_),
    .A(_0000_));
 sg13g2_inv_4 _2854_ (.A(net735),
    .Y(_1969_));
 sg13g2_inv_2 _2855_ (.Y(_1970_),
    .A(net733));
 sg13g2_inv_2 _2856_ (.Y(_1971_),
    .A(_0003_));
 sg13g2_inv_2 _2857_ (.Y(_1972_),
    .A(_0004_));
 sg13g2_inv_2 _2858_ (.Y(_1973_),
    .A(_0005_));
 sg13g2_inv_1 _2859_ (.Y(_1974_),
    .A(net558));
 sg13g2_inv_1 _2860_ (.Y(_1975_),
    .A(net606));
 sg13g2_inv_1 _2861_ (.Y(_1976_),
    .A(\core.dw[3] ));
 sg13g2_inv_1 _2862_ (.Y(_1977_),
    .A(net823));
 sg13g2_inv_1 _2863_ (.Y(_1978_),
    .A(_0035_));
 sg13g2_inv_1 _2864_ (.Y(_1979_),
    .A(net553));
 sg13g2_inv_1 _2865_ (.Y(_1980_),
    .A(net417));
 sg13g2_inv_1 _2866_ (.Y(_1981_),
    .A(net485));
 sg13g2_mux2_2 _2867_ (.A0(\core.vm8_reg[2] ),
    .A1(\core.w8_reg[2] ),
    .S(net1),
    .X(uo_out[1]));
 sg13g2_nor2_1 _2868_ (.A(net1),
    .B(\core.vm8_reg[3] ),
    .Y(_1982_));
 sg13g2_a21oi_2 _2869_ (.B1(_1982_),
    .Y(uo_out[5]),
    .A2(_1981_),
    .A1(net1));
 sg13g2_mux2_2 _2870_ (.A0(\core.vm8_reg[7] ),
    .A1(\core.w8_reg[7] ),
    .S(net1),
    .X(uo_out[6]));
 sg13g2_or4_1 _2871_ (.A(\core.w[1] ),
    .B(net708),
    .C(\core.w[13] ),
    .D(\core.w[12] ),
    .X(_1983_));
 sg13g2_nor3_2 _2872_ (.A(\core.w[3] ),
    .B(\core.w[2] ),
    .C(_1983_),
    .Y(_1984_));
 sg13g2_nor4_1 _2873_ (.A(\core.w[11] ),
    .B(\core.w[10] ),
    .C(\core.w[9] ),
    .D(\core.w[8] ),
    .Y(_1985_));
 sg13g2_nor4_1 _2874_ (.A(\core.w[7] ),
    .B(\core.w[6] ),
    .C(\core.w[5] ),
    .D(\core.w[4] ),
    .Y(_1986_));
 sg13g2_nand3_1 _2875_ (.B(_1985_),
    .C(_1986_),
    .A(_1984_),
    .Y(_1987_));
 sg13g2_nand3b_1 _2876_ (.B(\core.w[14] ),
    .C(_1987_),
    .Y(_1988_),
    .A_N(\core.w[15] ));
 sg13g2_nand2b_1 _2877_ (.Y(_1989_),
    .B(net820),
    .A_N(net763));
 sg13g2_and2_2 _2878_ (.A(_1988_),
    .B(_1989_),
    .X(_1990_));
 sg13g2_nand2_2 _2879_ (.Y(_1991_),
    .A(net783),
    .B(_1990_));
 sg13g2_nand4_1 _2880_ (.B(\core.V[13] ),
    .C(\core.V[12] ),
    .A(\core.V[14] ),
    .Y(_1992_),
    .D(\core.V[11] ));
 sg13g2_and2_1 _2881_ (.A(\core.VT_q[11] ),
    .B(_1992_),
    .X(_1993_));
 sg13g2_nor2_1 _2882_ (.A(_1922_),
    .B(\core.VT_q[9] ),
    .Y(_1994_));
 sg13g2_nand2b_1 _2883_ (.Y(_1995_),
    .B(\core.VT_q[6] ),
    .A_N(net712));
 sg13g2_o21ai_1 _2884_ (.B1(_1995_),
    .Y(_1996_),
    .A1(net308),
    .A2(_1945_));
 sg13g2_nor4_2 _2885_ (.A(net328),
    .B(net722),
    .C(net725),
    .Y(_1997_),
    .D(net726));
 sg13g2_nor2_1 _2886_ (.A(net313),
    .B(_1948_),
    .Y(_1998_));
 sg13g2_nand2b_1 _2887_ (.Y(_1999_),
    .B(\core.VT_q[5] ),
    .A_N(net314));
 sg13g2_a22oi_1 _2888_ (.Y(_2000_),
    .B1(_1948_),
    .B2(net313),
    .A2(_1947_),
    .A1(net314));
 sg13g2_o21ai_1 _2889_ (.B1(_2000_),
    .Y(_2001_),
    .A1(_1997_),
    .A2(_1998_));
 sg13g2_a22oi_1 _2890_ (.Y(_2002_),
    .B1(_1999_),
    .B2(_2001_),
    .A2(_1946_),
    .A1(net712));
 sg13g2_a22oi_1 _2891_ (.Y(_2003_),
    .B1(_1945_),
    .B2(net308),
    .A2(_1944_),
    .A1(\core.V[8] ));
 sg13g2_o21ai_1 _2892_ (.B1(_2003_),
    .Y(_2004_),
    .A1(_1996_),
    .A2(_2002_));
 sg13g2_a22oi_1 _2893_ (.Y(_2005_),
    .B1(\core.VT_q[8] ),
    .B2(_1923_),
    .A2(\core.VT_q[9] ),
    .A1(_1922_));
 sg13g2_a21o_1 _2894_ (.A2(_2005_),
    .A1(_2004_),
    .B1(_1994_),
    .X(_2006_));
 sg13g2_o21ai_1 _2895_ (.B1(_2006_),
    .Y(_2007_),
    .A1(\core.V[10] ),
    .A2(_1943_));
 sg13g2_or2_1 _2896_ (.X(_2008_),
    .B(\core.V[11] ),
    .A(\core.V[14] ));
 sg13g2_a22oi_1 _2897_ (.Y(_2009_),
    .B1(_2008_),
    .B2(_1942_),
    .A2(_1943_),
    .A1(\core.V[10] ));
 sg13g2_a221oi_1 _2898_ (.B2(_2009_),
    .C1(_1993_),
    .B1(_2007_),
    .A1(\core.V[15] ),
    .Y(_2010_),
    .A2(_1942_));
 sg13g2_nor2_1 _2899_ (.A(\core.V[13] ),
    .B(\core.V[12] ),
    .Y(_2011_));
 sg13g2_a21oi_1 _2900_ (.A1(_1942_),
    .A2(_2011_),
    .Y(_2012_),
    .B1(\core.V[15] ));
 sg13g2_nor2_2 _2901_ (.A(_2010_),
    .B(_2012_),
    .Y(_2013_));
 sg13g2_inv_1 _2902_ (.Y(_2014_),
    .A(net636));
 sg13g2_nand2_1 _2903_ (.Y(_2015_),
    .A(\core.b_q[4] ),
    .B(\core.w[4] ));
 sg13g2_nor2_1 _2904_ (.A(\core.b_q[4] ),
    .B(\core.w[4] ),
    .Y(_2016_));
 sg13g2_nor2_1 _2905_ (.A(net635),
    .B(_2016_),
    .Y(_2017_));
 sg13g2_xnor2_1 _2906_ (.Y(_2018_),
    .A(\core.w[2] ),
    .B(\core.dw[2] ));
 sg13g2_nand2_1 _2907_ (.Y(_2019_),
    .A(net708),
    .B(net472));
 sg13g2_xnor2_1 _2908_ (.Y(_2020_),
    .A(\core.w[1] ),
    .B(net498));
 sg13g2_nor2_1 _2909_ (.A(_2019_),
    .B(_2020_),
    .Y(_2021_));
 sg13g2_a21oi_1 _2910_ (.A1(\core.w[1] ),
    .A2(\core.dw[1] ),
    .Y(_2022_),
    .B1(_2021_));
 sg13g2_nor2_1 _2911_ (.A(_2018_),
    .B(_2022_),
    .Y(_2023_));
 sg13g2_a21oi_2 _2912_ (.B1(_2023_),
    .Y(_2024_),
    .A2(\core.dw[2] ),
    .A1(\core.w[2] ));
 sg13g2_xor2_1 _2913_ (.B(\core.dw[3] ),
    .A(\core.w[3] ),
    .X(_2025_));
 sg13g2_nand2b_1 _2914_ (.Y(_2026_),
    .B(_2025_),
    .A_N(_2024_));
 sg13g2_o21ai_1 _2915_ (.B1(_2026_),
    .Y(_2027_),
    .A1(_1919_),
    .A2(_1976_));
 sg13g2_and2_1 _2916_ (.A(\core.w[4] ),
    .B(\core.dw[4] ),
    .X(_2028_));
 sg13g2_xor2_1 _2917_ (.B(\core.dw[4] ),
    .A(\core.w[4] ),
    .X(_2029_));
 sg13g2_xor2_1 _2918_ (.B(_2029_),
    .A(_2027_),
    .X(_2030_));
 sg13g2_a22oi_1 _2919_ (.Y(_2031_),
    .B1(_2030_),
    .B2(net635),
    .A2(_2017_),
    .A1(_2015_));
 sg13g2_nor2_1 _2920_ (.A(net638),
    .B(_2031_),
    .Y(_2032_));
 sg13g2_a21oi_1 _2921_ (.A1(net782),
    .A2(net834),
    .Y(_2033_),
    .B1(_2032_));
 sg13g2_nor2_1 _2922_ (.A(net776),
    .B(_2033_),
    .Y(_0036_));
 sg13g2_nand2_1 _2923_ (.Y(_2034_),
    .A(\core.b_q[5] ),
    .B(\core.w[5] ));
 sg13g2_xnor2_1 _2924_ (.Y(_2035_),
    .A(\core.b_q[5] ),
    .B(\core.w[5] ));
 sg13g2_xnor2_1 _2925_ (.Y(_2036_),
    .A(_2015_),
    .B(_2035_));
 sg13g2_nand2_1 _2926_ (.Y(_2037_),
    .A(_2014_),
    .B(_2036_));
 sg13g2_a21oi_1 _2927_ (.A1(_2027_),
    .A2(_2029_),
    .Y(_2038_),
    .B1(_2028_));
 sg13g2_nand2_1 _2928_ (.Y(_2039_),
    .A(\core.w[5] ),
    .B(\core.dw[5] ));
 sg13g2_xnor2_1 _2929_ (.Y(_2040_),
    .A(\core.w[5] ),
    .B(\core.dw[5] ));
 sg13g2_xnor2_1 _2930_ (.Y(_2041_),
    .A(_2038_),
    .B(_2040_));
 sg13g2_a21oi_1 _2931_ (.A1(net634),
    .A2(_2041_),
    .Y(_2042_),
    .B1(net637));
 sg13g2_a22oi_1 _2932_ (.Y(_2043_),
    .B1(_2037_),
    .B2(_2042_),
    .A2(net849),
    .A1(net781));
 sg13g2_nor2_1 _2933_ (.A(net775),
    .B(_2043_),
    .Y(_0037_));
 sg13g2_nand2_1 _2934_ (.Y(_2044_),
    .A(net781),
    .B(net877));
 sg13g2_xnor2_1 _2935_ (.Y(_2045_),
    .A(\core.w[6] ),
    .B(\core.dw[6] ));
 sg13g2_nand2_1 _2936_ (.Y(_2046_),
    .A(_2038_),
    .B(_2039_));
 sg13g2_o21ai_1 _2937_ (.B1(_2046_),
    .Y(_2047_),
    .A1(\core.w[5] ),
    .A2(\core.dw[5] ));
 sg13g2_nor2_1 _2938_ (.A(_2045_),
    .B(_2047_),
    .Y(_2048_));
 sg13g2_xor2_1 _2939_ (.B(_2047_),
    .A(_2045_),
    .X(_2049_));
 sg13g2_o21ai_1 _2940_ (.B1(_2034_),
    .Y(_2050_),
    .A1(_2015_),
    .A2(_2035_));
 sg13g2_and2_1 _2941_ (.A(\core.b_q[6] ),
    .B(\core.w[6] ),
    .X(_2051_));
 sg13g2_xor2_1 _2942_ (.B(\core.w[6] ),
    .A(\core.b_q[6] ),
    .X(_2052_));
 sg13g2_xnor2_1 _2943_ (.Y(_2053_),
    .A(_2050_),
    .B(_2052_));
 sg13g2_nor2_1 _2944_ (.A(net635),
    .B(_2053_),
    .Y(_2054_));
 sg13g2_a21oi_1 _2945_ (.A1(net634),
    .A2(_2049_),
    .Y(_2055_),
    .B1(_2054_));
 sg13g2_o21ai_1 _2946_ (.B1(_2044_),
    .Y(_2056_),
    .A1(net637),
    .A2(_2055_));
 sg13g2_and2_1 _2947_ (.A(net810),
    .B(_2056_),
    .X(_0038_));
 sg13g2_nand2_1 _2948_ (.Y(_2057_),
    .A(net781),
    .B(net881));
 sg13g2_a21oi_1 _2949_ (.A1(_2050_),
    .A2(_2052_),
    .Y(_2058_),
    .B1(_2051_));
 sg13g2_xor2_1 _2950_ (.B(\core.w[7] ),
    .A(\core.b_q[7] ),
    .X(_2059_));
 sg13g2_nand2b_1 _2951_ (.Y(_2060_),
    .B(_2059_),
    .A_N(_2058_));
 sg13g2_xnor2_1 _2952_ (.Y(_2061_),
    .A(_2058_),
    .B(_2059_));
 sg13g2_a21oi_1 _2953_ (.A1(\core.w[6] ),
    .A2(\core.dw[6] ),
    .Y(_2062_),
    .B1(_2048_));
 sg13g2_xnor2_1 _2954_ (.Y(_2063_),
    .A(\core.w[7] ),
    .B(\core.dw[7] ));
 sg13g2_nand2_1 _2955_ (.Y(_2064_),
    .A(_2062_),
    .B(_2063_));
 sg13g2_nor2_1 _2956_ (.A(_2062_),
    .B(_2063_),
    .Y(_2065_));
 sg13g2_nor2_1 _2957_ (.A(net631),
    .B(_2065_),
    .Y(_2066_));
 sg13g2_a22oi_1 _2958_ (.Y(_2067_),
    .B1(_2064_),
    .B2(_2066_),
    .A2(_2061_),
    .A1(net631));
 sg13g2_o21ai_1 _2959_ (.B1(_2057_),
    .Y(_2068_),
    .A1(net638),
    .A2(_2067_));
 sg13g2_and2_1 _2960_ (.A(net810),
    .B(_2068_),
    .X(_0039_));
 sg13g2_nand2_1 _2961_ (.Y(_2069_),
    .A(net781),
    .B(net842));
 sg13g2_a21oi_1 _2962_ (.A1(\core.w[7] ),
    .A2(\core.dw[7] ),
    .Y(_2070_),
    .B1(_2065_));
 sg13g2_nand2_1 _2963_ (.Y(_2071_),
    .A(\core.w[8] ),
    .B(\core.dw[8] ));
 sg13g2_xnor2_1 _2964_ (.Y(_2072_),
    .A(\core.w[8] ),
    .B(\core.dw[8] ));
 sg13g2_xnor2_1 _2965_ (.Y(_2073_),
    .A(_2070_),
    .B(_2072_));
 sg13g2_o21ai_1 _2966_ (.B1(_2060_),
    .Y(_2074_),
    .A1(_1934_),
    .A2(_1956_));
 sg13g2_and2_1 _2967_ (.A(\core.b_q[8] ),
    .B(\core.w[8] ),
    .X(_2075_));
 sg13g2_xor2_1 _2968_ (.B(\core.w[8] ),
    .A(\core.b_q[8] ),
    .X(_2076_));
 sg13g2_xor2_1 _2969_ (.B(_2076_),
    .A(_2074_),
    .X(_2077_));
 sg13g2_a21oi_1 _2970_ (.A1(net635),
    .A2(_2073_),
    .Y(_2078_),
    .B1(net638));
 sg13g2_o21ai_1 _2971_ (.B1(_2078_),
    .Y(_2079_),
    .A1(net635),
    .A2(_2077_));
 sg13g2_a21oi_1 _2972_ (.A1(_2069_),
    .A2(_2079_),
    .Y(_0040_),
    .B1(net775));
 sg13g2_nand2_1 _2973_ (.Y(_2080_),
    .A(net781),
    .B(\core.w[9] ));
 sg13g2_o21ai_1 _2974_ (.B1(_2071_),
    .Y(_2081_),
    .A1(_2070_),
    .A2(_2072_));
 sg13g2_nor2_1 _2975_ (.A(\core.w[9] ),
    .B(\core.dw[9] ),
    .Y(_2082_));
 sg13g2_xnor2_1 _2976_ (.Y(_2083_),
    .A(\core.w[9] ),
    .B(\core.dw[9] ));
 sg13g2_o21ai_1 _2977_ (.B1(net634),
    .Y(_2084_),
    .A1(_2081_),
    .A2(_2083_));
 sg13g2_a21o_1 _2978_ (.A2(_2083_),
    .A1(_2081_),
    .B1(_2084_),
    .X(_2085_));
 sg13g2_nor2_2 _2979_ (.A(_1991_),
    .B(net630),
    .Y(_2086_));
 sg13g2_a21o_1 _2980_ (.A2(_2076_),
    .A1(_2074_),
    .B1(_2075_),
    .X(_2087_));
 sg13g2_xnor2_1 _2981_ (.Y(_2088_),
    .A(\core.b_q[9] ),
    .B(\core.w[9] ));
 sg13g2_xnor2_1 _2982_ (.Y(_2089_),
    .A(_2087_),
    .B(_2088_));
 sg13g2_o21ai_1 _2983_ (.B1(_2085_),
    .Y(_2090_),
    .A1(net634),
    .A2(_2089_));
 sg13g2_o21ai_1 _2984_ (.B1(_2080_),
    .Y(_2091_),
    .A1(net637),
    .A2(_2090_));
 sg13g2_and2_1 _2985_ (.A(net810),
    .B(_2091_),
    .X(_0041_));
 sg13g2_nand2_1 _2986_ (.Y(_2092_),
    .A(net781),
    .B(net833));
 sg13g2_xnor2_1 _2987_ (.Y(_2093_),
    .A(\core.w[10] ),
    .B(\core.dw[10] ));
 sg13g2_a21oi_1 _2988_ (.A1(\core.w[9] ),
    .A2(\core.dw[9] ),
    .Y(_2094_),
    .B1(_2081_));
 sg13g2_nor2_1 _2989_ (.A(_2082_),
    .B(_2094_),
    .Y(_2095_));
 sg13g2_nor3_1 _2990_ (.A(_2082_),
    .B(_2093_),
    .C(_2094_),
    .Y(_2096_));
 sg13g2_nand2_1 _2991_ (.Y(_2097_),
    .A(\core.b_q[10] ),
    .B(\core.w[10] ));
 sg13g2_xnor2_1 _2992_ (.Y(_2098_),
    .A(\core.b_q[10] ),
    .B(\core.w[10] ));
 sg13g2_a21o_1 _2993_ (.A2(\core.w[9] ),
    .A1(\core.b_q[9] ),
    .B1(_2087_),
    .X(_2099_));
 sg13g2_o21ai_1 _2994_ (.B1(_2099_),
    .Y(_2100_),
    .A1(\core.b_q[9] ),
    .A2(\core.w[9] ));
 sg13g2_xor2_1 _2995_ (.B(_2100_),
    .A(_2098_),
    .X(_2101_));
 sg13g2_xor2_1 _2996_ (.B(_2095_),
    .A(_2093_),
    .X(_2102_));
 sg13g2_a21oi_1 _2997_ (.A1(net634),
    .A2(_2102_),
    .Y(_2103_),
    .B1(net637));
 sg13g2_o21ai_1 _2998_ (.B1(_2103_),
    .Y(_2104_),
    .A1(net634),
    .A2(_2101_));
 sg13g2_a21oi_1 _2999_ (.A1(_2092_),
    .A2(_2104_),
    .Y(_0042_),
    .B1(net775));
 sg13g2_a21o_1 _3000_ (.A2(\core.dw[10] ),
    .A1(\core.w[10] ),
    .B1(_2096_),
    .X(_2105_));
 sg13g2_nor2_1 _3001_ (.A(\core.w[11] ),
    .B(\core.dw[11] ),
    .Y(_2106_));
 sg13g2_and2_1 _3002_ (.A(\core.w[11] ),
    .B(\core.dw[11] ),
    .X(_2107_));
 sg13g2_nor2_1 _3003_ (.A(_2106_),
    .B(_2107_),
    .Y(_2108_));
 sg13g2_o21ai_1 _3004_ (.B1(net634),
    .Y(_2109_),
    .A1(_2105_),
    .A2(_2108_));
 sg13g2_a21oi_1 _3005_ (.A1(_2105_),
    .A2(_2108_),
    .Y(_2110_),
    .B1(_2109_));
 sg13g2_o21ai_1 _3006_ (.B1(_2097_),
    .Y(_2111_),
    .A1(_2098_),
    .A2(_2100_));
 sg13g2_xor2_1 _3007_ (.B(\core.w[11] ),
    .A(\core.b_q[11] ),
    .X(_2112_));
 sg13g2_and2_1 _3008_ (.A(_2111_),
    .B(_2112_),
    .X(_2113_));
 sg13g2_o21ai_1 _3009_ (.B1(net631),
    .Y(_2114_),
    .A1(_2111_),
    .A2(_2112_));
 sg13g2_nor2_1 _3010_ (.A(_2113_),
    .B(_2114_),
    .Y(_2115_));
 sg13g2_nor2_1 _3011_ (.A(_2110_),
    .B(_2115_),
    .Y(_2116_));
 sg13g2_nor2_1 _3012_ (.A(net637),
    .B(_2116_),
    .Y(_2117_));
 sg13g2_a21oi_1 _3013_ (.A1(net781),
    .A2(net836),
    .Y(_2118_),
    .B1(_2117_));
 sg13g2_nor2_1 _3014_ (.A(net776),
    .B(_2118_),
    .Y(_0043_));
 sg13g2_nand2_1 _3015_ (.Y(_2119_),
    .A(net781),
    .B(net883));
 sg13g2_a21oi_1 _3016_ (.A1(\core.b_q[11] ),
    .A2(\core.w[11] ),
    .Y(_2120_),
    .B1(_2113_));
 sg13g2_nor2b_1 _3017_ (.A(_2120_),
    .B_N(\core.w[12] ),
    .Y(_2121_));
 sg13g2_xnor2_1 _3018_ (.Y(_2122_),
    .A(\core.w[12] ),
    .B(\core.dw[12] ));
 sg13g2_nor2_1 _3019_ (.A(_2105_),
    .B(_2107_),
    .Y(_2123_));
 sg13g2_nor3_1 _3020_ (.A(_2106_),
    .B(_2122_),
    .C(_2123_),
    .Y(_2124_));
 sg13g2_o21ai_1 _3021_ (.B1(_2122_),
    .Y(_2125_),
    .A1(_2106_),
    .A2(_2123_));
 sg13g2_xnor2_1 _3022_ (.Y(_2126_),
    .A(\core.w[12] ),
    .B(_2120_));
 sg13g2_nand2b_1 _3023_ (.Y(_2127_),
    .B(_2125_),
    .A_N(_2124_));
 sg13g2_a21oi_1 _3024_ (.A1(net634),
    .A2(_2127_),
    .Y(_2128_),
    .B1(net637));
 sg13g2_o21ai_1 _3025_ (.B1(_2128_),
    .Y(_2129_),
    .A1(net635),
    .A2(_2126_));
 sg13g2_a21oi_1 _3026_ (.A1(_2119_),
    .A2(_2129_),
    .Y(_0044_),
    .B1(net776));
 sg13g2_nand2_1 _3027_ (.Y(_2130_),
    .A(net782),
    .B(net880));
 sg13g2_a21oi_1 _3028_ (.A1(\core.w[12] ),
    .A2(\core.dw[12] ),
    .Y(_2131_),
    .B1(_2124_));
 sg13g2_nor2_1 _3029_ (.A(\core.w[13] ),
    .B(\core.dw[13] ),
    .Y(_2132_));
 sg13g2_xor2_1 _3030_ (.B(\core.dw[13] ),
    .A(\core.w[13] ),
    .X(_2133_));
 sg13g2_xnor2_1 _3031_ (.Y(_2134_),
    .A(_2131_),
    .B(_2133_));
 sg13g2_and2_1 _3032_ (.A(\core.w[13] ),
    .B(_2121_),
    .X(_2135_));
 sg13g2_xnor2_1 _3033_ (.Y(_2136_),
    .A(\core.w[13] ),
    .B(_2121_));
 sg13g2_a21oi_1 _3034_ (.A1(net631),
    .A2(_2136_),
    .Y(_2137_),
    .B1(net637));
 sg13g2_o21ai_1 _3035_ (.B1(_2137_),
    .Y(_2138_),
    .A1(net631),
    .A2(_2134_));
 sg13g2_a21oi_1 _3036_ (.A1(_2130_),
    .A2(_2138_),
    .Y(_0045_),
    .B1(net775));
 sg13g2_nor2_2 _3037_ (.A(net779),
    .B(net772),
    .Y(_2139_));
 sg13g2_nand2_1 _3038_ (.Y(_2140_),
    .A(net783),
    .B(net793));
 sg13g2_o21ai_1 _3039_ (.B1(net809),
    .Y(_2141_),
    .A1(net783),
    .A2(net763));
 sg13g2_xnor2_1 _3040_ (.Y(_2142_),
    .A(net763),
    .B(\core.dw[14] ));
 sg13g2_a221oi_1 _3041_ (.B2(\core.w[13] ),
    .C1(_2124_),
    .B1(\core.dw[13] ),
    .A1(\core.w[12] ),
    .Y(_2143_),
    .A2(\core.dw[12] ));
 sg13g2_o21ai_1 _3042_ (.B1(_2142_),
    .Y(_2144_),
    .A1(_2132_),
    .A2(_2143_));
 sg13g2_nor3_1 _3043_ (.A(_2132_),
    .B(_2142_),
    .C(_2143_),
    .Y(_2145_));
 sg13g2_nor2_1 _3044_ (.A(net631),
    .B(_2145_),
    .Y(_2146_));
 sg13g2_xor2_1 _3045_ (.B(_2135_),
    .A(net763),
    .X(_2147_));
 sg13g2_a221oi_1 _3046_ (.B2(net631),
    .C1(net637),
    .B1(_2147_),
    .A1(_2144_),
    .Y(_2148_),
    .A2(_2146_));
 sg13g2_nor2_1 _3047_ (.A(_2141_),
    .B(_2148_),
    .Y(_0046_));
 sg13g2_nand2_1 _3048_ (.Y(_2149_),
    .A(net820),
    .B(net809));
 sg13g2_a21oi_1 _3049_ (.A1(net763),
    .A2(\core.dw[14] ),
    .Y(_2150_),
    .B1(_2145_));
 sg13g2_xnor2_1 _3050_ (.Y(_2151_),
    .A(\core.w[15] ),
    .B(\core.dw[15] ));
 sg13g2_xnor2_1 _3051_ (.Y(_2152_),
    .A(_2150_),
    .B(_2151_));
 sg13g2_nand3_1 _3052_ (.B(_0035_),
    .C(_2135_),
    .A(net763),
    .Y(_2153_));
 sg13g2_a21oi_1 _3053_ (.A1(net763),
    .A2(_2135_),
    .Y(_2154_),
    .B1(_0035_));
 sg13g2_nor2_1 _3054_ (.A(net636),
    .B(_2154_),
    .Y(_2155_));
 sg13g2_a22oi_1 _3055_ (.Y(_2156_),
    .B1(_2153_),
    .B2(_2155_),
    .A2(_2152_),
    .A1(net636));
 sg13g2_a21oi_1 _3056_ (.A1(_1988_),
    .A2(_2156_),
    .Y(_2157_),
    .B1(net782));
 sg13g2_a22oi_1 _3057_ (.Y(_0047_),
    .B1(_2157_),
    .B2(net821),
    .A2(_2149_),
    .A1(net769));
 sg13g2_and2_1 _3058_ (.A(net3),
    .B(net808),
    .X(_0048_));
 sg13g2_nor2b_2 _3059_ (.A(\core.lstate[0] ),
    .B_N(_0016_),
    .Y(_2158_));
 sg13g2_nor2b_1 _3060_ (.A(\core.lstate[1] ),
    .B_N(_2158_),
    .Y(_2159_));
 sg13g2_nand2b_2 _3061_ (.Y(_2160_),
    .B(_2158_),
    .A_N(net707));
 sg13g2_nor2b_2 _3062_ (.A(\core.load_prev ),
    .B_N(net3),
    .Y(_2161_));
 sg13g2_inv_1 _3063_ (.Y(_2162_),
    .A(_2161_));
 sg13g2_nand2_1 _3064_ (.Y(_2163_),
    .A(net4),
    .B(_2161_));
 sg13g2_inv_1 _3065_ (.Y(_2164_),
    .A(_2163_));
 sg13g2_nand2_1 _3066_ (.Y(_2165_),
    .A(\core.lstate[0] ),
    .B(_0016_));
 sg13g2_nor2_1 _3067_ (.A(net707),
    .B(_2165_),
    .Y(_2166_));
 sg13g2_a22oi_1 _3068_ (.Y(_2167_),
    .B1(net677),
    .B2(_2161_),
    .A2(_2164_),
    .A1(net680));
 sg13g2_and3_1 _3069_ (.X(_2168_),
    .A(_0017_),
    .B(_2161_),
    .C(net678));
 sg13g2_nor2_2 _3070_ (.A(_2167_),
    .B(_2168_),
    .Y(_2169_));
 sg13g2_or2_1 _3071_ (.X(_2170_),
    .B(_2168_),
    .A(_2167_));
 sg13g2_a21oi_1 _3072_ (.A1(net5),
    .A2(net678),
    .Y(_2171_),
    .B1(_2170_));
 sg13g2_o21ai_1 _3073_ (.B1(net802),
    .Y(_2172_),
    .A1(net548),
    .A2(_2169_));
 sg13g2_nor2_1 _3074_ (.A(_2171_),
    .B(_2172_),
    .Y(_0049_));
 sg13g2_a21oi_1 _3075_ (.A1(net6),
    .A2(net678),
    .Y(_2173_),
    .B1(_2170_));
 sg13g2_o21ai_1 _3076_ (.B1(net802),
    .Y(_2174_),
    .A1(net568),
    .A2(_2169_));
 sg13g2_nor2_1 _3077_ (.A(_2173_),
    .B(_2174_),
    .Y(_0050_));
 sg13g2_a21oi_1 _3078_ (.A1(net7),
    .A2(net678),
    .Y(_2175_),
    .B1(_2170_));
 sg13g2_o21ai_1 _3079_ (.B1(net804),
    .Y(_2176_),
    .A1(net570),
    .A2(_2169_));
 sg13g2_nor2_1 _3080_ (.A(_2175_),
    .B(_2176_),
    .Y(_0051_));
 sg13g2_a21oi_1 _3081_ (.A1(net8),
    .A2(net678),
    .Y(_2177_),
    .B1(_2170_));
 sg13g2_o21ai_1 _3082_ (.B1(net802),
    .Y(_2178_),
    .A1(net575),
    .A2(_2169_));
 sg13g2_nor2_1 _3083_ (.A(_2177_),
    .B(_2178_),
    .Y(_0052_));
 sg13g2_mux2_1 _3084_ (.A0(net708),
    .A1(net603),
    .S(net764),
    .X(_0053_));
 sg13g2_nand2b_1 _3085_ (.Y(_2179_),
    .B(\core.leak[1] ),
    .A_N(\core.w[1] ));
 sg13g2_xor2_1 _3086_ (.B(\core.leak[1] ),
    .A(\core.w[1] ),
    .X(_2180_));
 sg13g2_xnor2_1 _3087_ (.Y(_2181_),
    .A(net708),
    .B(_2180_));
 sg13g2_nand2_1 _3088_ (.Y(_2182_),
    .A(net489),
    .B(net764));
 sg13g2_o21ai_1 _3089_ (.B1(_2182_),
    .Y(_0054_),
    .A1(net764),
    .A2(_2181_));
 sg13g2_nor2_1 _3090_ (.A(net458),
    .B(net681),
    .Y(_2183_));
 sg13g2_o21ai_1 _3091_ (.B1(_2179_),
    .Y(_2184_),
    .A1(\core.w[0] ),
    .A2(_2180_));
 sg13g2_nor2b_1 _3092_ (.A(\core.w[2] ),
    .B_N(\core.leak[2] ),
    .Y(_2185_));
 sg13g2_xnor2_1 _3093_ (.Y(_2186_),
    .A(\core.w[2] ),
    .B(\core.leak[2] ));
 sg13g2_xnor2_1 _3094_ (.Y(_2187_),
    .A(_2184_),
    .B(_2186_));
 sg13g2_a21oi_1 _3095_ (.A1(net681),
    .A2(_2187_),
    .Y(_0055_),
    .B1(_2183_));
 sg13g2_a21oi_1 _3096_ (.A1(_2184_),
    .A2(_2186_),
    .Y(_2188_),
    .B1(_2185_));
 sg13g2_xor2_1 _3097_ (.B(\core.leak[10] ),
    .A(\core.w[3] ),
    .X(_2189_));
 sg13g2_o21ai_1 _3098_ (.B1(net681),
    .Y(_2190_),
    .A1(_2188_),
    .A2(_2189_));
 sg13g2_a21oi_1 _3099_ (.A1(_2188_),
    .A2(_2189_),
    .Y(_2191_),
    .B1(_2190_));
 sg13g2_a21o_1 _3100_ (.A2(net764),
    .A1(net860),
    .B1(_2191_),
    .X(_0056_));
 sg13g2_mux2_1 _3101_ (.A0(net440),
    .A1(net763),
    .S(net807),
    .X(_0057_));
 sg13g2_o21ai_1 _3102_ (.B1(_2149_),
    .Y(_0058_),
    .A1(net807),
    .A2(_1981_));
 sg13g2_nor2_1 _3103_ (.A(net807),
    .B(net411),
    .Y(_2192_));
 sg13g2_a21oi_1 _3104_ (.A1(net807),
    .A2(_1978_),
    .Y(_0059_),
    .B1(_2192_));
 sg13g2_mux2_1 _3105_ (.A0(net421),
    .A1(\core.V[14] ),
    .S(net809),
    .X(_0060_));
 sg13g2_nor2_2 _3106_ (.A(\core.V[15] ),
    .B(net771),
    .Y(_2193_));
 sg13g2_a21oi_1 _3107_ (.A1(net775),
    .A2(_1980_),
    .Y(_0061_),
    .B1(_2193_));
 sg13g2_mux2_1 _3108_ (.A0(net382),
    .A1(_0034_),
    .S(net802),
    .X(_0062_));
 sg13g2_nand2_2 _3109_ (.Y(_2194_),
    .A(_1925_),
    .B(_1926_));
 sg13g2_or3_2 _3110_ (.A(\core.TauW_q[9] ),
    .B(net730),
    .C(_2194_),
    .X(_2195_));
 sg13g2_nand2_2 _3111_ (.Y(_2196_),
    .A(net727),
    .B(net738));
 sg13g2_and2_1 _3112_ (.A(net718),
    .B(net741),
    .X(_2197_));
 sg13g2_nand2_2 _3113_ (.Y(_2198_),
    .A(net723),
    .B(net740));
 sg13g2_nand2_2 _3114_ (.Y(_2199_),
    .A(net721),
    .B(net739));
 sg13g2_and4_1 _3115_ (.A(net721),
    .B(net724),
    .C(net739),
    .D(net740),
    .X(_2200_));
 sg13g2_a22oi_1 _3116_ (.Y(_2201_),
    .B1(net740),
    .B2(net720),
    .A2(net739),
    .A1(net724));
 sg13g2_nor2_2 _3117_ (.A(_2201_),
    .B(_2200_),
    .Y(_2202_));
 sg13g2_xor2_1 _3118_ (.B(_2197_),
    .A(_2202_),
    .X(_2203_));
 sg13g2_nand2b_1 _3119_ (.Y(_2204_),
    .B(_2203_),
    .A_N(_2196_));
 sg13g2_nand2_1 _3120_ (.Y(_2205_),
    .A(net725),
    .B(\core.a_q[11] ));
 sg13g2_nor2_2 _3121_ (.A(_2196_),
    .B(_2205_),
    .Y(_2206_));
 sg13g2_a22oi_1 _3122_ (.Y(_2207_),
    .B1(net738),
    .B2(net725),
    .A2(net312),
    .A1(net727));
 sg13g2_nor2_1 _3123_ (.A(_2206_),
    .B(_2207_),
    .Y(_2208_));
 sg13g2_nand2_1 _3124_ (.Y(_2209_),
    .A(net715),
    .B(net741));
 sg13g2_nand2_1 _3125_ (.Y(_2210_),
    .A(net719),
    .B(\core.a_q[9] ));
 sg13g2_nand2_2 _3126_ (.Y(_2211_),
    .A(net718),
    .B(net740));
 sg13g2_or2_1 _3127_ (.X(_2212_),
    .B(_2211_),
    .A(_2199_));
 sg13g2_xnor2_1 _3128_ (.Y(_2213_),
    .A(_2211_),
    .B(_2199_));
 sg13g2_xor2_1 _3129_ (.B(_2209_),
    .A(_2213_),
    .X(_2214_));
 sg13g2_nand2_1 _3130_ (.Y(_2215_),
    .A(_2208_),
    .B(net294));
 sg13g2_xnor2_1 _3131_ (.Y(_2216_),
    .A(_2208_),
    .B(_2214_));
 sg13g2_nor2_1 _3132_ (.A(net299),
    .B(net306),
    .Y(_2217_));
 sg13g2_xor2_1 _3133_ (.B(_2204_),
    .A(_2216_),
    .X(_2218_));
 sg13g2_nand2_2 _3134_ (.Y(_2219_),
    .A(net713),
    .B(net743));
 sg13g2_nand2_2 _3135_ (.Y(_2220_),
    .A(net742),
    .B(net715));
 sg13g2_nand2_2 _3136_ (.Y(_2221_),
    .A(net713),
    .B(net746));
 sg13g2_nand2_1 _3137_ (.Y(_2222_),
    .A(net711),
    .B(net748));
 sg13g2_xor2_1 _3138_ (.B(_2220_),
    .A(_2221_),
    .X(_2223_));
 sg13g2_nand2b_1 _3139_ (.Y(_2224_),
    .B(_2223_),
    .A_N(_2222_));
 sg13g2_o21ai_1 _3140_ (.B1(_2224_),
    .Y(_2225_),
    .A1(net321),
    .A2(_2221_));
 sg13g2_a21oi_2 _3141_ (.B1(_2200_),
    .Y(_2226_),
    .A2(_2202_),
    .A1(_2197_));
 sg13g2_nand2_1 _3142_ (.Y(_2227_),
    .A(net710),
    .B(net748));
 sg13g2_nand2_2 _3143_ (.Y(_2228_),
    .A(net711),
    .B(net744));
 sg13g2_nand2_2 _3144_ (.Y(_2229_),
    .A(net711),
    .B(net746));
 sg13g2_or2_1 _3145_ (.X(_2230_),
    .B(_2228_),
    .A(_2221_));
 sg13g2_xnor2_1 _3146_ (.Y(_2231_),
    .A(_2229_),
    .B(_2219_));
 sg13g2_xor2_1 _3147_ (.B(_2227_),
    .A(_2231_),
    .X(_2232_));
 sg13g2_nor2b_1 _3148_ (.A(_2226_),
    .B_N(net297),
    .Y(_2233_));
 sg13g2_xnor2_1 _3149_ (.Y(_2234_),
    .A(_2232_),
    .B(_2226_));
 sg13g2_xor2_1 _3150_ (.B(_2234_),
    .A(_2225_),
    .X(_2235_));
 sg13g2_a21oi_1 _3151_ (.A1(_2218_),
    .A2(_2235_),
    .Y(_2236_),
    .B1(_2217_));
 sg13g2_nand2_1 _3152_ (.Y(_2237_),
    .A(net721),
    .B(net311));
 sg13g2_and4_1 _3153_ (.A(\core.a_q[11] ),
    .B(net725),
    .C(net721),
    .D(net738),
    .X(_2238_));
 sg13g2_nand2_1 _3154_ (.Y(_2239_),
    .A(net721),
    .B(net738));
 sg13g2_a21oi_1 _3155_ (.A1(_2205_),
    .A2(_2239_),
    .Y(_2240_),
    .B1(_2238_));
 sg13g2_nor3_1 _3156_ (.A(_2196_),
    .B(_2205_),
    .C(net324),
    .Y(_2241_));
 sg13g2_xor2_1 _3157_ (.B(_2206_),
    .A(_2240_),
    .X(_2242_));
 sg13g2_nand2_1 _3158_ (.Y(_2243_),
    .A(net713),
    .B(net741));
 sg13g2_nand2_1 _3159_ (.Y(_2244_),
    .A(net716),
    .B(net739));
 sg13g2_nand2_2 _3160_ (.Y(_2245_),
    .A(net715),
    .B(\core.a_q[8] ));
 sg13g2_xor2_1 _3161_ (.B(_2245_),
    .A(_2210_),
    .X(_2246_));
 sg13g2_nand2b_1 _3162_ (.Y(_2247_),
    .B(_2246_),
    .A_N(_2243_));
 sg13g2_xnor2_1 _3163_ (.Y(_2248_),
    .A(_2246_),
    .B(_2243_));
 sg13g2_xnor2_1 _3164_ (.Y(_2249_),
    .A(_2242_),
    .B(_2248_));
 sg13g2_nor2_1 _3165_ (.A(_2215_),
    .B(net291),
    .Y(_2250_));
 sg13g2_xor2_1 _3166_ (.B(_2215_),
    .A(_2249_),
    .X(_2251_));
 sg13g2_o21ai_1 _3167_ (.B1(_2230_),
    .Y(_2252_),
    .A1(_2227_),
    .A2(net298));
 sg13g2_o21ai_1 _3168_ (.B1(_2212_),
    .Y(_2253_),
    .A1(_2209_),
    .A2(_2213_));
 sg13g2_nand2_1 _3169_ (.Y(_2254_),
    .A(net709),
    .B(net749));
 sg13g2_nand2_2 _3170_ (.Y(_2255_),
    .A(net710),
    .B(net747));
 sg13g2_xor2_1 _3171_ (.B(_2255_),
    .A(_2228_),
    .X(_2256_));
 sg13g2_nand2b_1 _3172_ (.Y(_2257_),
    .B(_2256_),
    .A_N(_2254_));
 sg13g2_xnor2_1 _3173_ (.Y(_2258_),
    .A(_2256_),
    .B(_2254_));
 sg13g2_xnor2_1 _3174_ (.Y(_2259_),
    .A(_2253_),
    .B(_2258_));
 sg13g2_nor2b_1 _3175_ (.A(net322),
    .B_N(_2252_),
    .Y(_0292_));
 sg13g2_xnor2_1 _3176_ (.Y(_0293_),
    .A(_2252_),
    .B(_2259_));
 sg13g2_xnor2_1 _3177_ (.Y(_0294_),
    .A(_0293_),
    .B(_2251_));
 sg13g2_nor2_1 _3178_ (.A(_2236_),
    .B(_0294_),
    .Y(_0295_));
 sg13g2_a21o_1 _3179_ (.A2(net301),
    .A1(_2225_),
    .B1(_2233_),
    .X(_0296_));
 sg13g2_xor2_1 _3180_ (.B(_0294_),
    .A(_2236_),
    .X(_0297_));
 sg13g2_a21oi_1 _3181_ (.A1(_0296_),
    .A2(net289),
    .Y(_0298_),
    .B1(_0295_));
 sg13g2_a21o_1 _3182_ (.A2(net307),
    .A1(_2253_),
    .B1(_0292_),
    .X(_0299_));
 sg13g2_a21oi_1 _3183_ (.A1(net288),
    .A2(_0293_),
    .Y(_0300_),
    .B1(_2250_));
 sg13g2_a21o_1 _3184_ (.A2(net296),
    .A1(net318),
    .B1(_2241_),
    .X(_0301_));
 sg13g2_nand2_1 _3185_ (.Y(_0302_),
    .A(net711),
    .B(net741));
 sg13g2_nand2_2 _3186_ (.Y(_0303_),
    .A(net713),
    .B(net740));
 sg13g2_xor2_1 _3187_ (.B(_0303_),
    .A(_2244_),
    .X(_0304_));
 sg13g2_nand2b_1 _3188_ (.Y(_0305_),
    .B(_0304_),
    .A_N(_0302_));
 sg13g2_xnor2_1 _3189_ (.Y(_0306_),
    .A(_0302_),
    .B(_0304_));
 sg13g2_nand2_2 _3190_ (.Y(_0307_),
    .A(net718),
    .B(net738));
 sg13g2_a21oi_1 _3191_ (.A1(net725),
    .A2(net738),
    .Y(_0308_),
    .B1(_2237_));
 sg13g2_xnor2_1 _3192_ (.Y(_0309_),
    .A(_0307_),
    .B(_0308_));
 sg13g2_xor2_1 _3193_ (.B(_0309_),
    .A(_0306_),
    .X(_0310_));
 sg13g2_nand2_1 _3194_ (.Y(_0311_),
    .A(_0301_),
    .B(_0310_));
 sg13g2_xnor2_1 _3195_ (.Y(_0312_),
    .A(_0301_),
    .B(_0310_));
 sg13g2_o21ai_1 _3196_ (.B1(_2257_),
    .Y(_0313_),
    .A1(_2228_),
    .A2(_2255_));
 sg13g2_o21ai_1 _3197_ (.B1(_2247_),
    .Y(_0314_),
    .A1(_2210_),
    .A2(net320));
 sg13g2_nand2_1 _3198_ (.Y(_0315_),
    .A(\core.V[9] ),
    .B(net748));
 sg13g2_nand2_2 _3199_ (.Y(_0316_),
    .A(net709),
    .B(net744));
 sg13g2_nor2_1 _3200_ (.A(_2255_),
    .B(_0316_),
    .Y(_0317_));
 sg13g2_or2_1 _3201_ (.X(_0318_),
    .B(_0316_),
    .A(_2255_));
 sg13g2_a22oi_1 _3202_ (.Y(_0319_),
    .B1(net747),
    .B2(net709),
    .A2(net744),
    .A1(net710));
 sg13g2_or2_1 _3203_ (.X(_0320_),
    .B(_0319_),
    .A(_0317_));
 sg13g2_xor2_1 _3204_ (.B(_0320_),
    .A(_0315_),
    .X(_0321_));
 sg13g2_xnor2_1 _3205_ (.Y(_0322_),
    .A(_0314_),
    .B(_0321_));
 sg13g2_nor2b_1 _3206_ (.A(_0322_),
    .B_N(_0313_),
    .Y(_0323_));
 sg13g2_xor2_1 _3207_ (.B(_0322_),
    .A(_0313_),
    .X(_0324_));
 sg13g2_xor2_1 _3208_ (.B(_0324_),
    .A(_0312_),
    .X(_0325_));
 sg13g2_nor2b_1 _3209_ (.A(_0300_),
    .B_N(_0325_),
    .Y(_0326_));
 sg13g2_xnor2_1 _3210_ (.Y(_0327_),
    .A(_0300_),
    .B(_0325_));
 sg13g2_xnor2_1 _3211_ (.Y(_0328_),
    .A(_0299_),
    .B(_0327_));
 sg13g2_nor2_1 _3212_ (.A(_0298_),
    .B(_0328_),
    .Y(_0329_));
 sg13g2_xnor2_1 _3213_ (.Y(_0330_),
    .A(_2196_),
    .B(_2203_));
 sg13g2_inv_1 _3214_ (.Y(_0331_),
    .A(_0330_));
 sg13g2_and4_1 _3215_ (.A(net745),
    .B(net718),
    .C(net743),
    .D(net715),
    .X(_0332_));
 sg13g2_nand2_1 _3216_ (.Y(_0333_),
    .A(net713),
    .B(net748));
 sg13g2_a22oi_1 _3217_ (.Y(_0334_),
    .B1(net746),
    .B2(net715),
    .A2(net742),
    .A1(net718));
 sg13g2_nor3_1 _3218_ (.A(_0332_),
    .B(_0333_),
    .C(_0334_),
    .Y(_0335_));
 sg13g2_or2_1 _3219_ (.X(_0336_),
    .B(_0335_),
    .A(net323));
 sg13g2_nand2_1 _3220_ (.Y(_0337_),
    .A(net726),
    .B(net739));
 sg13g2_or2_1 _3221_ (.X(_0338_),
    .B(_0337_),
    .A(_2198_));
 sg13g2_nand2_1 _3222_ (.Y(_0339_),
    .A(net720),
    .B(net741));
 sg13g2_and2_1 _3223_ (.A(_2198_),
    .B(_0337_),
    .X(_0340_));
 sg13g2_xor2_1 _3224_ (.B(_0337_),
    .A(_2198_),
    .X(_0341_));
 sg13g2_o21ai_1 _3225_ (.B1(_0338_),
    .Y(_0342_),
    .A1(_0340_),
    .A2(_0339_));
 sg13g2_xnor2_1 _3226_ (.Y(_0343_),
    .A(_2223_),
    .B(_2222_));
 sg13g2_and2_1 _3227_ (.A(net303),
    .B(net295),
    .X(_0344_));
 sg13g2_xor2_1 _3228_ (.B(_0343_),
    .A(_0342_),
    .X(_0345_));
 sg13g2_xnor2_1 _3229_ (.Y(_0346_),
    .A(_0345_),
    .B(_0336_));
 sg13g2_or2_1 _3230_ (.X(_0347_),
    .B(_0331_),
    .A(_0346_));
 sg13g2_xnor2_1 _3231_ (.Y(_0348_),
    .A(_2235_),
    .B(_2218_));
 sg13g2_nor2_1 _3232_ (.A(_0347_),
    .B(net304),
    .Y(_0349_));
 sg13g2_a21o_1 _3233_ (.A2(net292),
    .A1(_0336_),
    .B1(_0344_),
    .X(_0350_));
 sg13g2_xor2_1 _3234_ (.B(_0348_),
    .A(_0347_),
    .X(_0351_));
 sg13g2_a21oi_1 _3235_ (.A1(_0350_),
    .A2(_0351_),
    .Y(_0352_),
    .B1(_0349_));
 sg13g2_xnor2_1 _3236_ (.Y(_0353_),
    .A(_0297_),
    .B(_0296_));
 sg13g2_nor2_1 _3237_ (.A(_0352_),
    .B(_0353_),
    .Y(_0354_));
 sg13g2_inv_1 _3238_ (.Y(_0355_),
    .A(_0354_));
 sg13g2_xnor2_1 _3239_ (.Y(_0356_),
    .A(_0351_),
    .B(_0350_));
 sg13g2_nand2_1 _3240_ (.Y(_0357_),
    .A(net726),
    .B(net741));
 sg13g2_nor2_1 _3241_ (.A(net317),
    .B(_0357_),
    .Y(_0358_));
 sg13g2_o21ai_1 _3242_ (.B1(_0333_),
    .Y(_0359_),
    .A1(_0334_),
    .A2(_0332_));
 sg13g2_nor2b_2 _3243_ (.A(_0335_),
    .B_N(_0359_),
    .Y(_0360_));
 sg13g2_and4_1 _3244_ (.A(net718),
    .B(net720),
    .C(net742),
    .D(net746),
    .X(_0361_));
 sg13g2_nand2_1 _3245_ (.Y(_0362_),
    .A(net715),
    .B(net748));
 sg13g2_a22oi_1 _3246_ (.Y(_0363_),
    .B1(net745),
    .B2(net718),
    .A2(net743),
    .A1(net720));
 sg13g2_or3_1 _3247_ (.A(_0361_),
    .B(_0362_),
    .C(_0363_),
    .X(_0364_));
 sg13g2_nor2b_1 _3248_ (.A(_0361_),
    .B_N(_0364_),
    .Y(_0365_));
 sg13g2_xor2_1 _3249_ (.B(_0360_),
    .A(_0358_),
    .X(_0366_));
 sg13g2_nor2b_1 _3250_ (.A(_0365_),
    .B_N(net293),
    .Y(_0367_));
 sg13g2_a21o_1 _3251_ (.A2(_0360_),
    .A1(_0358_),
    .B1(_0367_),
    .X(_0368_));
 sg13g2_xnor2_1 _3252_ (.Y(_0369_),
    .A(_0339_),
    .B(_0341_));
 sg13g2_xnor2_1 _3253_ (.Y(_0370_),
    .A(_0366_),
    .B(_0365_));
 sg13g2_nand2_2 _3254_ (.Y(_0371_),
    .A(_0370_),
    .B(_0369_));
 sg13g2_xnor2_1 _3255_ (.Y(_0372_),
    .A(_0330_),
    .B(_0346_));
 sg13g2_nor2b_1 _3256_ (.A(net300),
    .B_N(_0372_),
    .Y(_0373_));
 sg13g2_inv_1 _3257_ (.Y(_0374_),
    .A(_0373_));
 sg13g2_xnor2_1 _3258_ (.Y(_0375_),
    .A(_0371_),
    .B(_0372_));
 sg13g2_and4_1 _3259_ (.A(net720),
    .B(net723),
    .C(net742),
    .D(net745),
    .X(_0376_));
 sg13g2_nand4_1 _3260_ (.B(net723),
    .C(net742),
    .A(net720),
    .Y(_0377_),
    .D(net745));
 sg13g2_a22oi_1 _3261_ (.Y(_0378_),
    .B1(net745),
    .B2(net720),
    .A2(net723),
    .A1(net742));
 sg13g2_and4_1 _3262_ (.A(net723),
    .B(net726),
    .C(net745),
    .D(net748),
    .X(_0379_));
 sg13g2_o21ai_1 _3263_ (.B1(_0379_),
    .Y(_0380_),
    .A1(_0376_),
    .A2(net302));
 sg13g2_or2_1 _3264_ (.X(_0381_),
    .B(_0380_),
    .A(_0357_));
 sg13g2_nand2_1 _3265_ (.Y(_0382_),
    .A(net718),
    .B(net748));
 sg13g2_or3_1 _3266_ (.A(_0376_),
    .B(_0378_),
    .C(_0382_),
    .X(_0383_));
 sg13g2_o21ai_1 _3267_ (.B1(_0382_),
    .Y(_0384_),
    .A1(_0376_),
    .A2(_0378_));
 sg13g2_nand4_1 _3268_ (.B(net727),
    .C(net330),
    .A(net723),
    .Y(_0385_),
    .D(net745));
 sg13g2_nand2_1 _3269_ (.Y(_0386_),
    .A(net720),
    .B(net748));
 sg13g2_a22oi_1 _3270_ (.Y(_0387_),
    .B1(net745),
    .B2(net723),
    .A2(net330),
    .A1(net726));
 sg13g2_a21oi_1 _3271_ (.A1(_0385_),
    .A2(_0386_),
    .Y(_0388_),
    .B1(_0387_));
 sg13g2_nand3_1 _3272_ (.B(_0384_),
    .C(_0388_),
    .A(_0383_),
    .Y(_0389_));
 sg13g2_nor2_1 _3273_ (.A(_0381_),
    .B(_0389_),
    .Y(_0390_));
 sg13g2_a22oi_1 _3274_ (.Y(_0391_),
    .B1(net741),
    .B2(net723),
    .A2(net740),
    .A1(net727));
 sg13g2_or2_1 _3275_ (.X(_0392_),
    .B(_0391_),
    .A(_0358_));
 sg13g2_o21ai_1 _3276_ (.B1(_0377_),
    .Y(_0393_),
    .A1(_0378_),
    .A2(_0382_));
 sg13g2_o21ai_1 _3277_ (.B1(_0362_),
    .Y(_0394_),
    .A1(_0361_),
    .A2(_0363_));
 sg13g2_a21oi_1 _3278_ (.A1(_0364_),
    .A2(_0394_),
    .Y(_0395_),
    .B1(_0393_));
 sg13g2_and3_1 _3279_ (.X(_0396_),
    .A(_0364_),
    .B(_0393_),
    .C(_0394_));
 sg13g2_o21ai_1 _3280_ (.B1(_0392_),
    .Y(_0397_),
    .A1(_0395_),
    .A2(_0396_));
 sg13g2_or3_1 _3281_ (.A(_0392_),
    .B(_0395_),
    .C(_0396_),
    .X(_0398_));
 sg13g2_a21oi_1 _3282_ (.A1(_0383_),
    .A2(_0384_),
    .Y(_0399_),
    .B1(_0388_));
 sg13g2_nand2_1 _3283_ (.Y(_0400_),
    .A(_0381_),
    .B(_0399_));
 sg13g2_nand3_1 _3284_ (.B(_0380_),
    .C(_0389_),
    .A(_0357_),
    .Y(_0401_));
 sg13g2_and4_1 _3285_ (.A(_0397_),
    .B(_0398_),
    .C(_0400_),
    .D(_0401_),
    .X(_0402_));
 sg13g2_nand2b_1 _3286_ (.Y(_0403_),
    .B(_0398_),
    .A_N(_0396_));
 sg13g2_nor3_1 _3287_ (.A(_0390_),
    .B(_0402_),
    .C(_0403_),
    .Y(_0404_));
 sg13g2_xnor2_1 _3288_ (.Y(_0405_),
    .A(_0369_),
    .B(_0370_));
 sg13g2_o21ai_1 _3289_ (.B1(_0403_),
    .Y(_0406_),
    .A1(_0390_),
    .A2(_0402_));
 sg13g2_a21oi_1 _3290_ (.A1(_0405_),
    .A2(_0406_),
    .Y(_0407_),
    .B1(_0404_));
 sg13g2_o21ai_1 _3291_ (.B1(_0407_),
    .Y(_0408_),
    .A1(_0375_),
    .A2(_0368_));
 sg13g2_nand2_1 _3292_ (.Y(_0409_),
    .A(_0368_),
    .B(_0375_));
 sg13g2_a21o_1 _3293_ (.A2(_0409_),
    .A1(_0408_),
    .B1(_0356_),
    .X(_0410_));
 sg13g2_a21o_1 _3294_ (.A2(_0356_),
    .A1(_0408_),
    .B1(_0374_),
    .X(_0411_));
 sg13g2_xnor2_1 _3295_ (.Y(_0412_),
    .A(_0352_),
    .B(_0353_));
 sg13g2_a21o_2 _3296_ (.A2(_0411_),
    .A1(_0410_),
    .B1(_0412_),
    .X(_0413_));
 sg13g2_xnor2_1 _3297_ (.Y(_0414_),
    .A(_0298_),
    .B(_0328_));
 sg13g2_a21oi_2 _3298_ (.B1(_0414_),
    .Y(_0415_),
    .A2(_0355_),
    .A1(_0413_));
 sg13g2_a21oi_2 _3299_ (.B1(_0326_),
    .Y(_0416_),
    .A2(_0327_),
    .A1(_0299_));
 sg13g2_a21o_1 _3300_ (.A2(_0321_),
    .A1(_0314_),
    .B1(_0323_),
    .X(_0417_));
 sg13g2_o21ai_1 _3301_ (.B1(_0311_),
    .Y(_0418_),
    .A1(_0312_),
    .A2(_0324_));
 sg13g2_a22oi_1 _3302_ (.Y(_0419_),
    .B1(_0306_),
    .B2(_0309_),
    .A2(net325),
    .A1(_1924_));
 sg13g2_nand2_1 _3303_ (.Y(_0420_),
    .A(net710),
    .B(\core.a_q[7] ));
 sg13g2_nand2_1 _3304_ (.Y(_0421_),
    .A(net711),
    .B(net739));
 sg13g2_nor2_1 _3305_ (.A(_0303_),
    .B(_0421_),
    .Y(_0422_));
 sg13g2_or2_1 _3306_ (.X(_0423_),
    .B(_0421_),
    .A(_0303_));
 sg13g2_a22oi_1 _3307_ (.Y(_0424_),
    .B1(net740),
    .B2(net711),
    .A2(net739),
    .A1(net713));
 sg13g2_nor2_1 _3308_ (.A(_0422_),
    .B(_0424_),
    .Y(_0425_));
 sg13g2_xnor2_1 _3309_ (.Y(_0426_),
    .A(_0420_),
    .B(_0425_));
 sg13g2_nand2_1 _3310_ (.Y(_0427_),
    .A(net716),
    .B(net738));
 sg13g2_nand3_1 _3311_ (.B(net310),
    .C(_2239_),
    .A(net719),
    .Y(_0428_));
 sg13g2_xor2_1 _3312_ (.B(_0428_),
    .A(_0427_),
    .X(_0429_));
 sg13g2_xnor2_1 _3313_ (.Y(_0430_),
    .A(_0426_),
    .B(_0429_));
 sg13g2_or2_1 _3314_ (.X(_0431_),
    .B(_0430_),
    .A(_0419_));
 sg13g2_xnor2_1 _3315_ (.Y(_0432_),
    .A(_0419_),
    .B(_0430_));
 sg13g2_o21ai_1 _3316_ (.B1(_0318_),
    .Y(_0433_),
    .A1(_0315_),
    .A2(_0320_));
 sg13g2_o21ai_1 _3317_ (.B1(_0305_),
    .Y(_0434_),
    .A1(_2244_),
    .A2(_0303_));
 sg13g2_nand2_1 _3318_ (.Y(_0435_),
    .A(\core.V[10] ),
    .B(net749));
 sg13g2_nand2_1 _3319_ (.Y(_0436_),
    .A(\core.V[9] ),
    .B(net744));
 sg13g2_nand2_1 _3320_ (.Y(_0437_),
    .A(\core.V[9] ),
    .B(net315));
 sg13g2_xor2_1 _3321_ (.B(_0437_),
    .A(_0316_),
    .X(_0438_));
 sg13g2_nand2b_1 _3322_ (.Y(_0439_),
    .B(_0438_),
    .A_N(_0435_));
 sg13g2_xnor2_1 _3323_ (.Y(_0440_),
    .A(_0435_),
    .B(_0438_));
 sg13g2_xnor2_1 _3324_ (.Y(_0441_),
    .A(_0434_),
    .B(_0440_));
 sg13g2_nor2b_1 _3325_ (.A(_0441_),
    .B_N(_0433_),
    .Y(_0442_));
 sg13g2_xor2_1 _3326_ (.B(_0441_),
    .A(_0433_),
    .X(_0443_));
 sg13g2_xnor2_1 _3327_ (.Y(_0444_),
    .A(_0432_),
    .B(_0443_));
 sg13g2_inv_1 _3328_ (.Y(_0445_),
    .A(_0444_));
 sg13g2_xor2_1 _3329_ (.B(_0444_),
    .A(_0418_),
    .X(_0446_));
 sg13g2_nor2b_1 _3330_ (.A(_0446_),
    .B_N(_0417_),
    .Y(_0447_));
 sg13g2_xor2_1 _3331_ (.B(_0446_),
    .A(_0417_),
    .X(_0448_));
 sg13g2_xor2_1 _3332_ (.B(_0448_),
    .A(_0416_),
    .X(_0449_));
 sg13g2_o21ai_1 _3333_ (.B1(_0449_),
    .Y(_0450_),
    .A1(_0415_),
    .A2(_0329_));
 sg13g2_or3_1 _3334_ (.A(_0329_),
    .B(_0415_),
    .C(_0449_),
    .X(_0451_));
 sg13g2_and3_1 _3335_ (.X(_0452_),
    .A(_1920_),
    .B(_0450_),
    .C(_0451_));
 sg13g2_nand3_1 _3336_ (.B(_0450_),
    .C(_0451_),
    .A(_1920_),
    .Y(_0453_));
 sg13g2_and3_1 _3337_ (.X(_0454_),
    .A(_0355_),
    .B(_0413_),
    .C(_0414_));
 sg13g2_nor3_2 _3338_ (.A(\core.w[1] ),
    .B(_0415_),
    .C(_0454_),
    .Y(_0455_));
 sg13g2_nand3_1 _3339_ (.B(_0411_),
    .C(_0412_),
    .A(_0410_),
    .Y(_0456_));
 sg13g2_nand2_2 _3340_ (.Y(_0457_),
    .A(_0413_),
    .B(_0456_));
 sg13g2_nand2_2 _3341_ (.Y(_0458_),
    .A(net708),
    .B(_0457_));
 sg13g2_o21ai_1 _3342_ (.B1(\core.w[1] ),
    .Y(_0459_),
    .A1(_0415_),
    .A2(_0454_));
 sg13g2_nor2b_2 _3343_ (.A(_0455_),
    .B_N(_0459_),
    .Y(_0460_));
 sg13g2_a21oi_1 _3344_ (.A1(_0458_),
    .A2(_0459_),
    .Y(_0461_),
    .B1(_0455_));
 sg13g2_a21oi_2 _3345_ (.B1(_1920_),
    .Y(_0462_),
    .A2(_0450_),
    .A1(_0451_));
 sg13g2_nor2_1 _3346_ (.A(_0452_),
    .B(_0462_),
    .Y(_0463_));
 sg13g2_o21ai_1 _3347_ (.B1(_0453_),
    .Y(_0464_),
    .A1(_0462_),
    .A2(_0461_));
 sg13g2_o21ai_1 _3348_ (.B1(_0450_),
    .Y(_0465_),
    .A1(_0416_),
    .A2(_0448_));
 sg13g2_a21oi_1 _3349_ (.A1(_0418_),
    .A2(_0445_),
    .Y(_0466_),
    .B1(_0447_));
 sg13g2_o21ai_1 _3350_ (.B1(_0431_),
    .Y(_0467_),
    .A1(_0432_),
    .A2(_0443_));
 sg13g2_xnor2_1 _3351_ (.Y(_0468_),
    .A(_1919_),
    .B(_0467_));
 sg13g2_a21oi_1 _3352_ (.A1(_0434_),
    .A2(_0440_),
    .Y(_0469_),
    .B1(_0442_));
 sg13g2_nand2_1 _3353_ (.Y(_0470_),
    .A(\core.V[11] ),
    .B(net749));
 sg13g2_nand2_1 _3354_ (.Y(_0471_),
    .A(\core.V[10] ),
    .B(net316));
 sg13g2_xnor2_1 _3355_ (.Y(_0472_),
    .A(_0436_),
    .B(_0471_));
 sg13g2_xnor2_1 _3356_ (.Y(_0473_),
    .A(_0470_),
    .B(_0472_));
 sg13g2_o21ai_1 _3357_ (.B1(_0439_),
    .Y(_0474_),
    .A1(_0316_),
    .A2(_0437_));
 sg13g2_o21ai_1 _3358_ (.B1(_0423_),
    .Y(_0475_),
    .A1(_0420_),
    .A2(_0424_));
 sg13g2_nor3_1 _3359_ (.A(net716),
    .B(_2237_),
    .C(_0307_),
    .Y(_0476_));
 sg13g2_a21oi_1 _3360_ (.A1(_0426_),
    .A2(_0429_),
    .Y(_0477_),
    .B1(_0476_));
 sg13g2_xnor2_1 _3361_ (.Y(_0478_),
    .A(_0475_),
    .B(_0477_));
 sg13g2_nand2_1 _3362_ (.Y(_0479_),
    .A(net710),
    .B(\core.a_q[8] ));
 sg13g2_xnor2_1 _3363_ (.Y(_0480_),
    .A(_0421_),
    .B(_0479_));
 sg13g2_nand2_1 _3364_ (.Y(_0481_),
    .A(net713),
    .B(net738));
 sg13g2_nand2_1 _3365_ (.Y(_0482_),
    .A(net709),
    .B(net741));
 sg13g2_xor2_1 _3366_ (.B(_0482_),
    .A(_0481_),
    .X(_0483_));
 sg13g2_xnor2_1 _3367_ (.Y(_0484_),
    .A(_0480_),
    .B(_0483_));
 sg13g2_nand3_1 _3368_ (.B(\core.a_q[11] ),
    .C(_0307_),
    .A(net716),
    .Y(_0485_));
 sg13g2_xnor2_1 _3369_ (.Y(_0486_),
    .A(_0473_),
    .B(_0484_));
 sg13g2_xnor2_1 _3370_ (.Y(_0487_),
    .A(_0474_),
    .B(_0485_));
 sg13g2_xnor2_1 _3371_ (.Y(_0488_),
    .A(_0486_),
    .B(_0487_));
 sg13g2_xnor2_1 _3372_ (.Y(_0489_),
    .A(_0478_),
    .B(_0488_));
 sg13g2_xnor2_1 _3373_ (.Y(_0490_),
    .A(_0469_),
    .B(_0489_));
 sg13g2_xnor2_1 _3374_ (.Y(_0491_),
    .A(_0468_),
    .B(_0490_));
 sg13g2_xnor2_1 _3375_ (.Y(_0492_),
    .A(_0466_),
    .B(_0491_));
 sg13g2_xnor2_1 _3376_ (.Y(_0493_),
    .A(_0492_),
    .B(_0465_));
 sg13g2_xor2_1 _3377_ (.B(_0464_),
    .A(_0493_),
    .X(_0494_));
 sg13g2_xnor2_1 _3378_ (.Y(_0495_),
    .A(_0493_),
    .B(_0464_));
 sg13g2_xnor2_1 _3379_ (.Y(_0496_),
    .A(_0461_),
    .B(_0463_));
 sg13g2_xor2_1 _3380_ (.B(_0457_),
    .A(net708),
    .X(_0497_));
 sg13g2_nand2_2 _3381_ (.Y(_0498_),
    .A(_0460_),
    .B(_0497_));
 sg13g2_nand3_1 _3382_ (.B(_1927_),
    .C(_0000_),
    .A(_1926_),
    .Y(_0499_));
 sg13g2_or3_1 _3383_ (.A(net730),
    .B(net731),
    .C(_0499_),
    .X(_0500_));
 sg13g2_nand3b_1 _3384_ (.B(net684),
    .C(net685),
    .Y(_0501_),
    .A_N(_0500_));
 sg13g2_nor2_1 _3385_ (.A(net683),
    .B(_0501_),
    .Y(_0502_));
 sg13g2_nor4_2 _3386_ (.A(_0502_),
    .B(_0496_),
    .C(_0498_),
    .Y(_0503_),
    .D(net628));
 sg13g2_nand2_1 _3387_ (.Y(_0504_),
    .A(net733),
    .B(net286));
 sg13g2_and2_1 _3388_ (.A(net627),
    .B(_0498_),
    .X(_0505_));
 sg13g2_nand3_1 _3389_ (.B(_0496_),
    .C(_0498_),
    .A(net627),
    .Y(_0506_));
 sg13g2_a21o_1 _3390_ (.A2(_0498_),
    .A1(net627),
    .B1(_0496_),
    .X(_0507_));
 sg13g2_nand2_1 _3391_ (.Y(_0508_),
    .A(_0506_),
    .B(_0507_));
 sg13g2_inv_1 _3392_ (.Y(_0509_),
    .A(_0508_));
 sg13g2_a21o_1 _3393_ (.A2(_0507_),
    .A1(_0506_),
    .B1(net735),
    .X(_0510_));
 sg13g2_nand4_1 _3394_ (.B(net735),
    .C(_0506_),
    .A(net736),
    .Y(_0511_),
    .D(_0507_));
 sg13g2_xnor2_1 _3395_ (.Y(_0512_),
    .A(_1969_),
    .B(_0508_));
 sg13g2_and2_1 _3396_ (.A(_0510_),
    .B(_0511_),
    .X(_0513_));
 sg13g2_xnor2_1 _3397_ (.Y(_0514_),
    .A(\core.TauW_q[5] ),
    .B(_0503_));
 sg13g2_nand3_1 _3398_ (.B(_0511_),
    .C(_0510_),
    .A(_0514_),
    .Y(_0515_));
 sg13g2_nand3b_1 _3399_ (.B(net685),
    .C(net687),
    .Y(_0516_),
    .A_N(_2195_));
 sg13g2_a21oi_2 _3400_ (.B1(_0516_),
    .Y(_0517_),
    .A2(_0504_),
    .A1(_0515_));
 sg13g2_a21o_2 _3401_ (.A2(_0515_),
    .A1(_0504_),
    .B1(_0516_),
    .X(_0518_));
 sg13g2_nor2_1 _3402_ (.A(_0503_),
    .B(_0517_),
    .Y(_0519_));
 sg13g2_xnor2_1 _3403_ (.Y(_0520_),
    .A(_0513_),
    .B(_0514_));
 sg13g2_a21oi_2 _3404_ (.B1(_0519_),
    .Y(_0521_),
    .A2(_0520_),
    .A1(_0517_));
 sg13g2_xor2_1 _3405_ (.B(_0460_),
    .A(_0458_),
    .X(_0522_));
 sg13g2_nand2b_1 _3406_ (.Y(_0523_),
    .B(_0522_),
    .A_N(_0497_));
 sg13g2_a22oi_1 _3407_ (.Y(_0524_),
    .B1(_0523_),
    .B2(_0505_),
    .A2(_0522_),
    .A1(net628));
 sg13g2_and2_1 _3408_ (.A(net736),
    .B(_0524_),
    .X(_0525_));
 sg13g2_mux2_1 _3409_ (.A0(_0509_),
    .A1(_0512_),
    .S(_0517_),
    .X(_0526_));
 sg13g2_xnor2_1 _3410_ (.Y(_0527_),
    .A(_0526_),
    .B(net733));
 sg13g2_nand2_1 _3411_ (.Y(_0528_),
    .A(net684),
    .B(_0526_));
 sg13g2_o21ai_1 _3412_ (.B1(_0528_),
    .Y(_0529_),
    .A1(_0527_),
    .A2(_0525_));
 sg13g2_xnor2_1 _3413_ (.Y(_0530_),
    .A(net732),
    .B(_0521_));
 sg13g2_a22oi_1 _3414_ (.Y(_0531_),
    .B1(_0530_),
    .B2(_0529_),
    .A2(_0521_),
    .A1(_0003_));
 sg13g2_nor2_2 _3415_ (.A(_0500_),
    .B(_0531_),
    .Y(_0532_));
 sg13g2_xor2_1 _3416_ (.B(_0530_),
    .A(net285),
    .X(_0533_));
 sg13g2_mux2_1 _3417_ (.A0(_0521_),
    .A1(_0533_),
    .S(_0532_),
    .X(_0534_));
 sg13g2_nand2_1 _3418_ (.Y(_0535_),
    .A(_0004_),
    .B(_0534_));
 sg13g2_nor3_2 _3419_ (.A(_0531_),
    .B(_0500_),
    .C(net683),
    .Y(_0536_));
 sg13g2_xnor2_1 _3420_ (.Y(_0537_),
    .A(_0524_),
    .B(_0536_));
 sg13g2_and2_1 _3421_ (.A(net684),
    .B(_0537_),
    .X(_0538_));
 sg13g2_inv_1 _3422_ (.Y(_0539_),
    .A(_0538_));
 sg13g2_xnor2_1 _3423_ (.Y(_0540_),
    .A(_0537_),
    .B(net684));
 sg13g2_nand2_1 _3424_ (.Y(_0541_),
    .A(net736),
    .B(_0497_));
 sg13g2_or2_1 _3425_ (.X(_0542_),
    .B(_0497_),
    .A(net736));
 sg13g2_nand2b_1 _3426_ (.Y(_0543_),
    .B(_1969_),
    .A_N(_0542_));
 sg13g2_nand3b_1 _3427_ (.B(_0541_),
    .C(_0543_),
    .Y(_0544_),
    .A_N(_0540_));
 sg13g2_xor2_1 _3428_ (.B(_0527_),
    .A(_0525_),
    .X(_0545_));
 sg13g2_mux2_1 _3429_ (.A0(_0526_),
    .A1(_0545_),
    .S(_0532_),
    .X(_0546_));
 sg13g2_xnor2_1 _3430_ (.Y(_0547_),
    .A(_1971_),
    .B(_0546_));
 sg13g2_inv_1 _3431_ (.Y(_0548_),
    .A(_0547_));
 sg13g2_a21oi_2 _3432_ (.B1(_0548_),
    .Y(_0549_),
    .A2(_0539_),
    .A1(_0544_));
 sg13g2_and2_1 _3433_ (.A(net685),
    .B(_0546_),
    .X(_0550_));
 sg13g2_nor2_1 _3434_ (.A(_0549_),
    .B(_0550_),
    .Y(_0551_));
 sg13g2_xnor2_1 _3435_ (.Y(_0552_),
    .A(net687),
    .B(_0534_));
 sg13g2_inv_1 _3436_ (.Y(_0553_),
    .A(_0552_));
 sg13g2_o21ai_1 _3437_ (.B1(_0553_),
    .Y(_0554_),
    .A1(_0550_),
    .A2(_0549_));
 sg13g2_a21oi_2 _3438_ (.B1(_2195_),
    .Y(_0555_),
    .A2(_0535_),
    .A1(_0554_));
 sg13g2_a21o_1 _3439_ (.A2(_0554_),
    .A1(_0535_),
    .B1(_2195_),
    .X(_0556_));
 sg13g2_xnor2_1 _3440_ (.Y(_0557_),
    .A(_0540_),
    .B(_0541_));
 sg13g2_mux2_2 _3441_ (.A0(_0537_),
    .A1(_0557_),
    .S(_0555_),
    .X(_0558_));
 sg13g2_nand2_1 _3442_ (.Y(_0559_),
    .A(_0534_),
    .B(_0556_));
 sg13g2_xnor2_1 _3443_ (.Y(_0560_),
    .A(_0551_),
    .B(_0552_));
 sg13g2_o21ai_1 _3444_ (.B1(_0559_),
    .Y(_0561_),
    .A1(_0556_),
    .A2(_0560_));
 sg13g2_nand2_1 _3445_ (.Y(_0562_),
    .A(_0005_),
    .B(_0561_));
 sg13g2_nor2_1 _3446_ (.A(_0546_),
    .B(_0555_),
    .Y(_0563_));
 sg13g2_nand3_1 _3447_ (.B(_0544_),
    .C(_0548_),
    .A(_0539_),
    .Y(_0564_));
 sg13g2_nand2b_1 _3448_ (.Y(_0565_),
    .B(_0564_),
    .A_N(_0549_));
 sg13g2_a21oi_2 _3449_ (.B1(_0563_),
    .Y(_0566_),
    .A2(_0565_),
    .A1(_0555_));
 sg13g2_and2_1 _3450_ (.A(_1928_),
    .B(_0566_),
    .X(_0567_));
 sg13g2_nor2_1 _3451_ (.A(net686),
    .B(_0558_),
    .Y(_0568_));
 sg13g2_nand2_1 _3452_ (.Y(_0569_),
    .A(net686),
    .B(_0558_));
 sg13g2_a221oi_1 _3453_ (.B2(_0554_),
    .C1(_2195_),
    .B1(_0535_),
    .A1(net736),
    .Y(_0570_),
    .A2(_0497_));
 sg13g2_a22oi_1 _3454_ (.Y(_0571_),
    .B1(_0570_),
    .B2(_0542_),
    .A2(_0556_),
    .A1(_0497_));
 sg13g2_inv_1 _3455_ (.Y(_0572_),
    .A(_0571_));
 sg13g2_nand2_1 _3456_ (.Y(_0573_),
    .A(_1930_),
    .B(_0571_));
 sg13g2_and2_1 _3457_ (.A(_0569_),
    .B(_0573_),
    .X(_0574_));
 sg13g2_a21o_1 _3458_ (.A2(_0573_),
    .A1(_0569_),
    .B1(_0568_),
    .X(_0575_));
 sg13g2_xnor2_1 _3459_ (.Y(_0576_),
    .A(_1970_),
    .B(_0571_));
 sg13g2_xnor2_1 _3460_ (.Y(_0577_),
    .A(_0558_),
    .B(\core.TauW_q[6] ));
 sg13g2_nand3_1 _3461_ (.B(_0576_),
    .C(_1931_),
    .A(_0577_),
    .Y(_0578_));
 sg13g2_xnor2_1 _3462_ (.Y(_0579_),
    .A(_0004_),
    .B(_0566_));
 sg13g2_inv_1 _3463_ (.Y(_0580_),
    .A(_0579_));
 sg13g2_a21oi_2 _3464_ (.B1(_0579_),
    .Y(_0581_),
    .A2(_0575_),
    .A1(_0578_));
 sg13g2_xor2_1 _3465_ (.B(_0561_),
    .A(net729),
    .X(_0582_));
 sg13g2_inv_1 _3466_ (.Y(_0583_),
    .A(_0582_));
 sg13g2_o21ai_1 _3467_ (.B1(_0583_),
    .Y(_0584_),
    .A1(_0581_),
    .A2(_0567_));
 sg13g2_a21oi_2 _3468_ (.B1(_0499_),
    .Y(_0585_),
    .A2(_0562_),
    .A1(_0584_));
 sg13g2_nand2_1 _3469_ (.Y(_0586_),
    .A(net734),
    .B(_0576_));
 sg13g2_nand2_1 _3470_ (.Y(_0587_),
    .A(_0573_),
    .B(_0586_));
 sg13g2_xor2_1 _3471_ (.B(_0587_),
    .A(_0577_),
    .X(_0588_));
 sg13g2_mux2_1 _3472_ (.A0(_0558_),
    .A1(_0588_),
    .S(net626),
    .X(_0589_));
 sg13g2_inv_1 _3473_ (.Y(_0590_),
    .A(_0589_));
 sg13g2_nor2_1 _3474_ (.A(\core.TauW_q[7] ),
    .B(_0590_),
    .Y(_0591_));
 sg13g2_nor2_2 _3475_ (.A(\core.TauW_q[5] ),
    .B(net736),
    .Y(_0592_));
 sg13g2_nand2_2 _3476_ (.Y(_0593_),
    .A(net684),
    .B(net683));
 sg13g2_and2_1 _3477_ (.A(_1969_),
    .B(_0585_),
    .X(_0594_));
 sg13g2_a21oi_1 _3478_ (.A1(_0002_),
    .A2(_0594_),
    .Y(_0595_),
    .B1(_0592_));
 sg13g2_xnor2_1 _3479_ (.Y(_0596_),
    .A(net734),
    .B(_0576_));
 sg13g2_mux2_1 _3480_ (.A0(_0572_),
    .A1(_0596_),
    .S(net626),
    .X(_0597_));
 sg13g2_xnor2_1 _3481_ (.Y(_0598_),
    .A(_1971_),
    .B(_0597_));
 sg13g2_nand2b_1 _3482_ (.Y(_0599_),
    .B(net685),
    .A_N(_0597_));
 sg13g2_o21ai_1 _3483_ (.B1(_0599_),
    .Y(_0600_),
    .A1(_0598_),
    .A2(_0595_));
 sg13g2_xnor2_1 _3484_ (.Y(_0601_),
    .A(\core.TauW_q[7] ),
    .B(_0589_));
 sg13g2_a21oi_2 _3485_ (.B1(_0591_),
    .Y(_0602_),
    .A2(_0600_),
    .A1(_0601_));
 sg13g2_nor2_1 _3486_ (.A(_0566_),
    .B(net626),
    .Y(_0603_));
 sg13g2_a21oi_1 _3487_ (.A1(_0574_),
    .A2(_0586_),
    .Y(_0604_),
    .B1(_0568_));
 sg13g2_xnor2_1 _3488_ (.Y(_0605_),
    .A(_0580_),
    .B(_0604_));
 sg13g2_a21oi_2 _3489_ (.B1(_0603_),
    .Y(_0606_),
    .A2(_0605_),
    .A1(net626));
 sg13g2_xnor2_1 _3490_ (.Y(_0607_),
    .A(_0005_),
    .B(_0606_));
 sg13g2_nand2b_1 _3491_ (.Y(_0608_),
    .B(_0606_),
    .A_N(net729));
 sg13g2_o21ai_1 _3492_ (.B1(_0608_),
    .Y(_0609_),
    .A1(_0607_),
    .A2(_0602_));
 sg13g2_a21oi_1 _3493_ (.A1(_0580_),
    .A2(_0604_),
    .Y(_0610_),
    .B1(_0567_));
 sg13g2_xnor2_1 _3494_ (.Y(_0611_),
    .A(_0582_),
    .B(_0610_));
 sg13g2_nand2_1 _3495_ (.Y(_0612_),
    .A(net626),
    .B(_0611_));
 sg13g2_o21ai_1 _3496_ (.B1(_0612_),
    .Y(_0613_),
    .A1(_0561_),
    .A2(net626));
 sg13g2_xnor2_1 _3497_ (.Y(_0614_),
    .A(\core.TauW_q[9] ),
    .B(_0613_));
 sg13g2_inv_1 _3498_ (.Y(_0615_),
    .A(_0614_));
 sg13g2_nand2b_1 _3499_ (.Y(_0616_),
    .B(_0006_),
    .A_N(_0613_));
 sg13g2_inv_1 _3500_ (.Y(_0617_),
    .A(_0616_));
 sg13g2_a21oi_2 _3501_ (.B1(_0617_),
    .Y(_0618_),
    .A2(_0609_),
    .A1(_0615_));
 sg13g2_or2_2 _3502_ (.X(_0619_),
    .B(_0618_),
    .A(_2194_));
 sg13g2_inv_2 _3503_ (.Y(_0620_),
    .A(_0619_));
 sg13g2_xnor2_1 _3504_ (.Y(_0621_),
    .A(_0600_),
    .B(_0601_));
 sg13g2_mux2_1 _3505_ (.A0(_0621_),
    .A1(_0590_),
    .S(_0619_),
    .X(_0622_));
 sg13g2_nand2_1 _3506_ (.Y(_0623_),
    .A(net729),
    .B(_0622_));
 sg13g2_nor2_1 _3507_ (.A(net729),
    .B(_0622_),
    .Y(_0624_));
 sg13g2_xnor2_1 _3508_ (.Y(_0625_),
    .A(net729),
    .B(_0622_));
 sg13g2_xnor2_1 _3509_ (.Y(_0626_),
    .A(_0595_),
    .B(_0598_));
 sg13g2_mux2_1 _3510_ (.A0(_0626_),
    .A1(_0597_),
    .S(_0619_),
    .X(_0627_));
 sg13g2_nand2_1 _3511_ (.Y(_0628_),
    .A(_0004_),
    .B(_0627_));
 sg13g2_nand2b_1 _3512_ (.Y(_0629_),
    .B(_1972_),
    .A_N(_0627_));
 sg13g2_and2_1 _3513_ (.A(_0628_),
    .B(_0629_),
    .X(_0630_));
 sg13g2_inv_1 _3514_ (.Y(_0631_),
    .A(_0630_));
 sg13g2_nor2_1 _3515_ (.A(_0625_),
    .B(_0630_),
    .Y(_0632_));
 sg13g2_o21ai_1 _3516_ (.B1(_0594_),
    .Y(_0633_),
    .A1(_0618_),
    .A2(_2194_));
 sg13g2_nor2_1 _3517_ (.A(net734),
    .B(net626),
    .Y(_0634_));
 sg13g2_xnor2_1 _3518_ (.Y(_0635_),
    .A(_1970_),
    .B(_0634_));
 sg13g2_or3_1 _3519_ (.A(_2194_),
    .B(_0618_),
    .C(_0635_),
    .X(_0636_));
 sg13g2_nand2_1 _3520_ (.Y(_0637_),
    .A(_0633_),
    .B(_0636_));
 sg13g2_a21oi_2 _3521_ (.B1(net732),
    .Y(_0638_),
    .A2(_0633_),
    .A1(_0636_));
 sg13g2_and3_1 _3522_ (.X(_0639_),
    .A(net732),
    .B(_0633_),
    .C(_0636_));
 sg13g2_nand3_1 _3523_ (.B(_0633_),
    .C(_0636_),
    .A(net732),
    .Y(_0640_));
 sg13g2_nand2b_1 _3524_ (.Y(_0641_),
    .B(_0640_),
    .A_N(_0638_));
 sg13g2_nor3_1 _3525_ (.A(net734),
    .B(_2194_),
    .C(_0618_),
    .Y(_0642_));
 sg13g2_nand2_1 _3526_ (.Y(_0643_),
    .A(_1969_),
    .B(_0620_));
 sg13g2_xnor2_1 _3527_ (.Y(_0644_),
    .A(_0002_),
    .B(_0642_));
 sg13g2_or4_1 _3528_ (.A(net737),
    .B(_0639_),
    .C(_0638_),
    .D(_0644_),
    .X(_0645_));
 sg13g2_and2_1 _3529_ (.A(net684),
    .B(_0642_),
    .X(_0646_));
 sg13g2_a21oi_1 _3530_ (.A1(_0640_),
    .A2(_0646_),
    .Y(_0647_),
    .B1(_0638_));
 sg13g2_nand2_1 _3531_ (.Y(_0648_),
    .A(_0645_),
    .B(_0647_));
 sg13g2_a221oi_1 _3532_ (.B2(_0645_),
    .C1(_0625_),
    .B1(_0647_),
    .A1(_0628_),
    .Y(_0649_),
    .A2(_0629_));
 sg13g2_nor2_1 _3533_ (.A(net731),
    .B(_0627_),
    .Y(_0650_));
 sg13g2_a21o_1 _3534_ (.A2(_0650_),
    .A1(_0623_),
    .B1(_0624_),
    .X(_0651_));
 sg13g2_xnor2_1 _3535_ (.Y(_0652_),
    .A(_0602_),
    .B(_0607_));
 sg13g2_nand2_1 _3536_ (.Y(_0653_),
    .A(_0606_),
    .B(_0619_));
 sg13g2_o21ai_1 _3537_ (.B1(_0653_),
    .Y(_0654_),
    .A1(_0619_),
    .A2(_0652_));
 sg13g2_xor2_1 _3538_ (.B(_0654_),
    .A(_0006_),
    .X(_0655_));
 sg13g2_o21ai_1 _3539_ (.B1(_0655_),
    .Y(_0656_),
    .A1(_0651_),
    .A2(_0649_));
 sg13g2_nand2_1 _3540_ (.Y(_0657_),
    .A(_1927_),
    .B(_0654_));
 sg13g2_xnor2_1 _3541_ (.Y(_0658_),
    .A(_0609_),
    .B(_0615_));
 sg13g2_mux2_1 _3542_ (.A0(_0658_),
    .A1(_0613_),
    .S(_0619_),
    .X(_0659_));
 sg13g2_xnor2_1 _3543_ (.Y(_0660_),
    .A(\core.TauW_q[10] ),
    .B(_0659_));
 sg13g2_a21o_1 _3544_ (.A2(_0656_),
    .A1(_0657_),
    .B1(_0660_),
    .X(_0661_));
 sg13g2_nand2b_1 _3545_ (.Y(_0662_),
    .B(_0007_),
    .A_N(_0659_));
 sg13g2_nor2_1 _3546_ (.A(_0645_),
    .B(_0660_),
    .Y(_0663_));
 sg13g2_nand4_1 _3547_ (.B(_0632_),
    .C(_0655_),
    .A(_1925_),
    .Y(_0664_),
    .D(_0663_));
 sg13g2_a22oi_1 _3548_ (.Y(_0665_),
    .B1(_0664_),
    .B2(_1968_),
    .A2(_0662_),
    .A1(_0661_));
 sg13g2_nand2_1 _3549_ (.Y(_0666_),
    .A(_1969_),
    .B(net621));
 sg13g2_nor2_1 _3550_ (.A(_0659_),
    .B(net622),
    .Y(_0667_));
 sg13g2_nand3_1 _3551_ (.B(_0657_),
    .C(_0660_),
    .A(_0656_),
    .Y(_0668_));
 sg13g2_and2_1 _3552_ (.A(_0661_),
    .B(_0668_),
    .X(_0669_));
 sg13g2_a21oi_2 _3553_ (.B1(_0667_),
    .Y(_0670_),
    .A2(_0669_),
    .A1(net622));
 sg13g2_and2_1 _3554_ (.A(_1968_),
    .B(_0670_),
    .X(_0671_));
 sg13g2_inv_1 _3555_ (.Y(_0672_),
    .A(_0671_));
 sg13g2_nor2_1 _3556_ (.A(_1968_),
    .B(_0670_),
    .Y(_0673_));
 sg13g2_a21oi_1 _3557_ (.A1(_0631_),
    .A2(_0648_),
    .Y(_0674_),
    .B1(_0650_));
 sg13g2_xor2_1 _3558_ (.B(_0674_),
    .A(_0625_),
    .X(_0675_));
 sg13g2_nand2_1 _3559_ (.Y(_0676_),
    .A(net622),
    .B(_0675_));
 sg13g2_o21ai_1 _3560_ (.B1(_0676_),
    .Y(_0677_),
    .A1(_0622_),
    .A2(_0665_));
 sg13g2_nand2_1 _3561_ (.Y(_0678_),
    .A(_1927_),
    .B(_0677_));
 sg13g2_nor2_1 _3562_ (.A(_0592_),
    .B(_0646_),
    .Y(_0679_));
 sg13g2_xor2_1 _3563_ (.B(_0679_),
    .A(_0641_),
    .X(_0680_));
 sg13g2_mux2_1 _3564_ (.A0(_0637_),
    .A1(_0680_),
    .S(net621),
    .X(_0681_));
 sg13g2_nand2_1 _3565_ (.Y(_0682_),
    .A(_0004_),
    .B(_0681_));
 sg13g2_nand2_1 _3566_ (.Y(_0683_),
    .A(net735),
    .B(_1970_));
 sg13g2_o21ai_1 _3567_ (.B1(_0683_),
    .Y(_0684_),
    .A1(net735),
    .A2(_0644_));
 sg13g2_inv_1 _3568_ (.Y(_0685_),
    .A(_0684_));
 sg13g2_mux2_1 _3569_ (.A0(_0643_),
    .A1(_0685_),
    .S(net621),
    .X(_0686_));
 sg13g2_inv_1 _3570_ (.Y(_0687_),
    .A(_0686_));
 sg13g2_o21ai_1 _3571_ (.B1(_0593_),
    .Y(_0688_),
    .A1(_1970_),
    .A2(_0666_));
 sg13g2_xnor2_1 _3572_ (.Y(_0689_),
    .A(_0003_),
    .B(_0686_));
 sg13g2_a22oi_1 _3573_ (.Y(_0690_),
    .B1(_0688_),
    .B2(_0689_),
    .A2(_0687_),
    .A1(net686));
 sg13g2_xnor2_1 _3574_ (.Y(_0691_),
    .A(net687),
    .B(_0681_));
 sg13g2_o21ai_1 _3575_ (.B1(_0682_),
    .Y(_0692_),
    .A1(_0691_),
    .A2(_0690_));
 sg13g2_xnor2_1 _3576_ (.Y(_0693_),
    .A(_0630_),
    .B(_0648_));
 sg13g2_nor2_1 _3577_ (.A(_0627_),
    .B(net622),
    .Y(_0694_));
 sg13g2_a21oi_2 _3578_ (.B1(_0694_),
    .Y(_0695_),
    .A2(_0693_),
    .A1(net621));
 sg13g2_xnor2_1 _3579_ (.Y(_0696_),
    .A(_1973_),
    .B(_0695_));
 sg13g2_inv_1 _3580_ (.Y(_0697_),
    .A(_0696_));
 sg13g2_nor2_1 _3581_ (.A(net729),
    .B(_0695_),
    .Y(_0698_));
 sg13g2_a21oi_2 _3582_ (.B1(_0698_),
    .Y(_0699_),
    .A2(_0692_),
    .A1(_0697_));
 sg13g2_xnor2_1 _3583_ (.Y(_0700_),
    .A(_1927_),
    .B(_0677_));
 sg13g2_o21ai_1 _3584_ (.B1(_0678_),
    .Y(_0701_),
    .A1(_0700_),
    .A2(_0699_));
 sg13g2_or3_1 _3585_ (.A(_0649_),
    .B(_0651_),
    .C(_0655_),
    .X(_0702_));
 sg13g2_nand2_1 _3586_ (.Y(_0703_),
    .A(_0656_),
    .B(_0702_));
 sg13g2_nor2_1 _3587_ (.A(_0654_),
    .B(net622),
    .Y(_0704_));
 sg13g2_a21oi_2 _3588_ (.B1(_0704_),
    .Y(_0705_),
    .A2(_0703_),
    .A1(net622));
 sg13g2_xor2_1 _3589_ (.B(_0705_),
    .A(_0007_),
    .X(_0706_));
 sg13g2_and2_1 _3590_ (.A(_1926_),
    .B(_0705_),
    .X(_0707_));
 sg13g2_a21o_1 _3591_ (.A2(_0706_),
    .A1(_0701_),
    .B1(_0707_),
    .X(_0708_));
 sg13g2_a221oi_1 _3592_ (.B2(_0706_),
    .C1(_0673_),
    .B1(_0701_),
    .A1(_1926_),
    .Y(_0709_),
    .A2(_0705_));
 sg13g2_nor2_2 _3593_ (.A(_0671_),
    .B(_0709_),
    .Y(_0710_));
 sg13g2_nor2_1 _3594_ (.A(net734),
    .B(net621),
    .Y(_0711_));
 sg13g2_xnor2_1 _3595_ (.Y(_0712_),
    .A(_0002_),
    .B(_0711_));
 sg13g2_a221oi_1 _3596_ (.B2(_0708_),
    .C1(_0673_),
    .B1(_0672_),
    .A1(_1969_),
    .Y(_0713_),
    .A2(net621));
 sg13g2_o21ai_1 _3597_ (.B1(_0666_),
    .Y(_0714_),
    .A1(net620),
    .A2(net618));
 sg13g2_nor3_2 _3598_ (.A(net620),
    .B(net618),
    .C(_0712_),
    .Y(_0715_));
 sg13g2_or3_1 _3599_ (.A(net620),
    .B(net618),
    .C(_0712_),
    .X(_0716_));
 sg13g2_xor2_1 _3600_ (.B(_0706_),
    .A(_0701_),
    .X(_0717_));
 sg13g2_mux2_1 _3601_ (.A0(_0705_),
    .A1(_0717_),
    .S(_0710_),
    .X(_0718_));
 sg13g2_nor2_1 _3602_ (.A(_0000_),
    .B(_0718_),
    .Y(_0719_));
 sg13g2_xnor2_1 _3603_ (.Y(_0720_),
    .A(_0690_),
    .B(_0691_));
 sg13g2_o21ai_1 _3604_ (.B1(_0681_),
    .Y(_0721_),
    .A1(net618),
    .A2(net620));
 sg13g2_or3_1 _3605_ (.A(net620),
    .B(net618),
    .C(_0720_),
    .X(_0722_));
 sg13g2_and2_1 _3606_ (.A(_0721_),
    .B(_0722_),
    .X(_0723_));
 sg13g2_and3_1 _3607_ (.X(_0724_),
    .A(_0721_),
    .B(\core.TauW_q[8] ),
    .C(_0722_));
 sg13g2_nand2_1 _3608_ (.Y(_0725_),
    .A(net729),
    .B(_0723_));
 sg13g2_a21oi_2 _3609_ (.B1(net730),
    .Y(_0726_),
    .A2(_0722_),
    .A1(_0721_));
 sg13g2_or2_1 _3610_ (.X(_0727_),
    .B(_0726_),
    .A(_0724_));
 sg13g2_xnor2_1 _3611_ (.Y(_0728_),
    .A(_0688_),
    .B(_0689_));
 sg13g2_o21ai_1 _3612_ (.B1(_0687_),
    .Y(_0729_),
    .A1(net620),
    .A2(net618));
 sg13g2_or3_1 _3613_ (.A(net620),
    .B(_0728_),
    .C(net618),
    .X(_0730_));
 sg13g2_and2_1 _3614_ (.A(_0729_),
    .B(_0730_),
    .X(_0731_));
 sg13g2_a21oi_1 _3615_ (.A1(_0729_),
    .A2(_0730_),
    .Y(_0732_),
    .B1(_1972_));
 sg13g2_and3_1 _3616_ (.X(_0733_),
    .A(_1972_),
    .B(_0729_),
    .C(_0730_));
 sg13g2_or2_1 _3617_ (.X(_0734_),
    .B(_0733_),
    .A(_0732_));
 sg13g2_nor4_2 _3618_ (.A(_0733_),
    .B(_0726_),
    .C(_0732_),
    .Y(_0735_),
    .D(_0724_));
 sg13g2_a21oi_1 _3619_ (.A1(_0714_),
    .A2(_0716_),
    .Y(_0736_),
    .B1(net686));
 sg13g2_o21ai_1 _3620_ (.B1(net732),
    .Y(_0737_),
    .A1(_0713_),
    .A2(_0715_));
 sg13g2_nor3_1 _3621_ (.A(net732),
    .B(_0713_),
    .C(_0715_),
    .Y(_0738_));
 sg13g2_nor3_2 _3622_ (.A(net734),
    .B(net620),
    .C(net618),
    .Y(_0739_));
 sg13g2_and2_1 _3623_ (.A(net684),
    .B(_0739_),
    .X(_0740_));
 sg13g2_a21o_1 _3624_ (.A2(_0740_),
    .A1(_0737_),
    .B1(_0738_),
    .X(_0741_));
 sg13g2_a21oi_1 _3625_ (.A1(_0737_),
    .A2(_0740_),
    .Y(_0742_),
    .B1(_0738_));
 sg13g2_nor2_1 _3626_ (.A(net731),
    .B(_0731_),
    .Y(_0743_));
 sg13g2_a221oi_1 _3627_ (.B2(_0725_),
    .C1(_0726_),
    .B1(_0743_),
    .A1(_0741_),
    .Y(_0744_),
    .A2(_0735_));
 sg13g2_nor2_1 _3628_ (.A(_0736_),
    .B(_0738_),
    .Y(_0745_));
 sg13g2_xnor2_1 _3629_ (.Y(_0746_),
    .A(_1970_),
    .B(_0739_));
 sg13g2_nand4_1 _3630_ (.B(net683),
    .C(_0745_),
    .A(_0735_),
    .Y(_0747_),
    .D(_0746_));
 sg13g2_xor2_1 _3631_ (.B(_0700_),
    .A(_0699_),
    .X(_0748_));
 sg13g2_mux2_2 _3632_ (.A0(_0677_),
    .A1(_0748_),
    .S(_0710_),
    .X(_0749_));
 sg13g2_nand2_1 _3633_ (.Y(_0750_),
    .A(_1926_),
    .B(_0749_));
 sg13g2_nor2_1 _3634_ (.A(_1926_),
    .B(_0749_),
    .Y(_0751_));
 sg13g2_xnor2_1 _3635_ (.Y(_0752_),
    .A(\core.TauW_q[10] ),
    .B(_0749_));
 sg13g2_xnor2_1 _3636_ (.Y(_0753_),
    .A(_0692_),
    .B(_0697_));
 sg13g2_or3_1 _3637_ (.A(_0671_),
    .B(net290),
    .C(_0753_),
    .X(_0754_));
 sg13g2_o21ai_1 _3638_ (.B1(_0754_),
    .Y(_0755_),
    .A1(_0695_),
    .A2(_0710_));
 sg13g2_xor2_1 _3639_ (.B(_0755_),
    .A(_0006_),
    .X(_0756_));
 sg13g2_nand2_1 _3640_ (.Y(_0757_),
    .A(_0752_),
    .B(_0756_));
 sg13g2_a21o_1 _3641_ (.A2(_0744_),
    .A1(_0747_),
    .B1(_0757_),
    .X(_0758_));
 sg13g2_and2_1 _3642_ (.A(_1927_),
    .B(_0755_),
    .X(_0759_));
 sg13g2_nand2b_1 _3643_ (.Y(_0760_),
    .B(_0759_),
    .A_N(_0751_));
 sg13g2_and2_1 _3644_ (.A(_0750_),
    .B(_0760_),
    .X(_0761_));
 sg13g2_a21oi_2 _3645_ (.B1(_0719_),
    .Y(_0762_),
    .A2(_0758_),
    .A1(_0761_));
 sg13g2_a21o_2 _3646_ (.A2(_0761_),
    .A1(_0758_),
    .B1(_0719_),
    .X(_0763_));
 sg13g2_and2_1 _3647_ (.A(_0000_),
    .B(_0718_),
    .X(_0764_));
 sg13g2_nor2_1 _3648_ (.A(_0670_),
    .B(_0710_),
    .Y(_0765_));
 sg13g2_a21oi_2 _3649_ (.B1(_0765_),
    .Y(_0766_),
    .A2(_0708_),
    .A1(_0673_));
 sg13g2_nor2b_2 _3650_ (.A(_0764_),
    .B_N(_0766_),
    .Y(_0767_));
 sg13g2_nand2b_2 _3651_ (.Y(_0768_),
    .B(_0766_),
    .A_N(_0764_));
 sg13g2_nor2_2 _3652_ (.A(_0768_),
    .B(_0762_),
    .Y(_0769_));
 sg13g2_nand2_2 _3653_ (.Y(_0770_),
    .A(_0763_),
    .B(_0767_));
 sg13g2_nor4_2 _3654_ (.A(_0713_),
    .B(_0715_),
    .C(_0762_),
    .Y(_0771_),
    .D(_0768_));
 sg13g2_nor2_1 _3655_ (.A(_0592_),
    .B(_0740_),
    .Y(_0772_));
 sg13g2_xnor2_1 _3656_ (.Y(_0773_),
    .A(_0745_),
    .B(_0772_));
 sg13g2_a21oi_2 _3657_ (.B1(_0771_),
    .Y(_0774_),
    .A2(_0773_),
    .A1(_0770_));
 sg13g2_a21o_1 _3658_ (.A2(_0773_),
    .A1(_0770_),
    .B1(_0771_),
    .X(_0775_));
 sg13g2_nand2_1 _3659_ (.Y(_0776_),
    .A(_1969_),
    .B(_0746_));
 sg13g2_nand2_1 _3660_ (.Y(_0777_),
    .A(_0683_),
    .B(_0776_));
 sg13g2_nand3_1 _3661_ (.B(_0763_),
    .C(_0767_),
    .A(_0739_),
    .Y(_0778_));
 sg13g2_o21ai_1 _3662_ (.B1(_0777_),
    .Y(_0779_),
    .A1(_0768_),
    .A2(_0762_));
 sg13g2_nand2_1 _3663_ (.Y(_0780_),
    .A(_0778_),
    .B(_0779_));
 sg13g2_inv_1 _3664_ (.Y(_0781_),
    .A(_0780_));
 sg13g2_a21oi_2 _3665_ (.B1(_1971_),
    .Y(_0782_),
    .A2(_0778_),
    .A1(_0779_));
 sg13g2_nand3_1 _3666_ (.B(_0778_),
    .C(_0779_),
    .A(_1971_),
    .Y(_0783_));
 sg13g2_nor2b_1 _3667_ (.A(_0782_),
    .B_N(_0783_),
    .Y(_0784_));
 sg13g2_a21oi_2 _3668_ (.B1(\core.TauW_q[5] ),
    .Y(_0785_),
    .A2(_0769_),
    .A1(net736));
 sg13g2_nand3b_1 _3669_ (.B(_0785_),
    .C(_0783_),
    .Y(_0786_),
    .A_N(_0782_));
 sg13g2_a22oi_1 _3670_ (.Y(_0787_),
    .B1(_0780_),
    .B2(net685),
    .A2(_0775_),
    .A1(_1928_));
 sg13g2_and2_1 _3671_ (.A(_0786_),
    .B(_0787_),
    .X(_0788_));
 sg13g2_nor2_1 _3672_ (.A(net687),
    .B(_0775_),
    .Y(_0789_));
 sg13g2_nand3b_1 _3673_ (.B(_0763_),
    .C(_0767_),
    .Y(_0790_),
    .A_N(_0723_));
 sg13g2_nand3_1 _3674_ (.B(net734),
    .C(net733),
    .A(net685),
    .Y(_0791_));
 sg13g2_a21oi_1 _3675_ (.A1(_0742_),
    .A2(_0791_),
    .Y(_0792_),
    .B1(_0734_));
 sg13g2_nor2_1 _3676_ (.A(_0743_),
    .B(_0792_),
    .Y(_0793_));
 sg13g2_xor2_1 _3677_ (.B(_0793_),
    .A(_0727_),
    .X(_0794_));
 sg13g2_o21ai_1 _3678_ (.B1(_0794_),
    .Y(_0795_),
    .A1(_0762_),
    .A2(_0768_));
 sg13g2_and2_1 _3679_ (.A(_0790_),
    .B(_0795_),
    .X(_0796_));
 sg13g2_nand3_1 _3680_ (.B(_0790_),
    .C(_0795_),
    .A(\core.TauW_q[9] ),
    .Y(_0797_));
 sg13g2_nor2_1 _3681_ (.A(\core.TauW_q[9] ),
    .B(_0796_),
    .Y(_0798_));
 sg13g2_a21o_1 _3682_ (.A2(_0795_),
    .A1(_0790_),
    .B1(\core.TauW_q[9] ),
    .X(_0799_));
 sg13g2_nand2_1 _3683_ (.Y(_0800_),
    .A(_0797_),
    .B(_0799_));
 sg13g2_nand3_1 _3684_ (.B(_0742_),
    .C(_0791_),
    .A(_0734_),
    .Y(_0801_));
 sg13g2_nand2b_1 _3685_ (.Y(_0802_),
    .B(_0801_),
    .A_N(_0792_));
 sg13g2_nor3_1 _3686_ (.A(_0731_),
    .B(_0762_),
    .C(_0768_),
    .Y(_0803_));
 sg13g2_a21oi_1 _3687_ (.A1(_0763_),
    .A2(_0767_),
    .Y(_0804_),
    .B1(_0802_));
 sg13g2_nor2_1 _3688_ (.A(_0803_),
    .B(_0804_),
    .Y(_0805_));
 sg13g2_inv_1 _3689_ (.Y(_0806_),
    .A(_0805_));
 sg13g2_o21ai_1 _3690_ (.B1(_0005_),
    .Y(_0807_),
    .A1(_0803_),
    .A2(_0804_));
 sg13g2_or3_1 _3691_ (.A(_0005_),
    .B(_0803_),
    .C(_0804_),
    .X(_0808_));
 sg13g2_nand2_1 _3692_ (.Y(_0809_),
    .A(_0807_),
    .B(_0808_));
 sg13g2_nand4_1 _3693_ (.B(_0799_),
    .C(_0807_),
    .A(_0797_),
    .Y(_0810_),
    .D(_0808_));
 sg13g2_a221oi_1 _3694_ (.B2(_0786_),
    .C1(_0810_),
    .B1(_0787_),
    .A1(net731),
    .Y(_0811_),
    .A2(_0774_));
 sg13g2_nor2_1 _3695_ (.A(net730),
    .B(_0805_),
    .Y(_0812_));
 sg13g2_a21o_1 _3696_ (.A2(_0812_),
    .A1(_0797_),
    .B1(_0798_),
    .X(_0813_));
 sg13g2_or2_1 _3697_ (.X(_0814_),
    .B(_0813_),
    .A(_0811_));
 sg13g2_nand4_1 _3698_ (.B(net733),
    .C(_0735_),
    .A(net734),
    .Y(_0815_),
    .D(_0745_));
 sg13g2_nand2_1 _3699_ (.Y(_0816_),
    .A(_0744_),
    .B(_0815_));
 sg13g2_a21oi_1 _3700_ (.A1(_0756_),
    .A2(_0816_),
    .Y(_0817_),
    .B1(_0759_));
 sg13g2_xnor2_1 _3701_ (.Y(_0818_),
    .A(_0752_),
    .B(_0817_));
 sg13g2_mux2_2 _3702_ (.A0(_0749_),
    .A1(_0818_),
    .S(_0770_),
    .X(_0819_));
 sg13g2_nor2_1 _3703_ (.A(_1925_),
    .B(_0819_),
    .Y(_0820_));
 sg13g2_xnor2_1 _3704_ (.Y(_0821_),
    .A(_1925_),
    .B(_0819_));
 sg13g2_nand3_1 _3705_ (.B(_0763_),
    .C(_0767_),
    .A(_0755_),
    .Y(_0822_));
 sg13g2_xnor2_1 _3706_ (.Y(_0823_),
    .A(_0756_),
    .B(_0816_));
 sg13g2_o21ai_1 _3707_ (.B1(_0822_),
    .Y(_0824_),
    .A1(_0823_),
    .A2(_0769_));
 sg13g2_inv_1 _3708_ (.Y(_0825_),
    .A(_0824_));
 sg13g2_xor2_1 _3709_ (.B(_0824_),
    .A(_0007_),
    .X(_0826_));
 sg13g2_nor2b_2 _3710_ (.A(_0821_),
    .B_N(_0826_),
    .Y(_0827_));
 sg13g2_o21ai_1 _3711_ (.B1(_0827_),
    .Y(_0828_),
    .A1(_0813_),
    .A2(_0811_));
 sg13g2_nor3_1 _3712_ (.A(\core.TauW_q[10] ),
    .B(_0820_),
    .C(_0825_),
    .Y(_0829_));
 sg13g2_a21oi_1 _3713_ (.A1(_1925_),
    .A2(_0819_),
    .Y(_0830_),
    .B1(_0829_));
 sg13g2_or2_1 _3714_ (.X(_0831_),
    .B(_0764_),
    .A(_0719_));
 sg13g2_a21oi_1 _3715_ (.A1(_0750_),
    .A2(_0817_),
    .Y(_0832_),
    .B1(_0751_));
 sg13g2_nor2b_1 _3716_ (.A(_0831_),
    .B_N(_0832_),
    .Y(_0833_));
 sg13g2_nor2_1 _3717_ (.A(_0764_),
    .B(_0833_),
    .Y(_0834_));
 sg13g2_nand2_1 _3718_ (.Y(_0835_),
    .A(_0762_),
    .B(_0766_));
 sg13g2_mux2_1 _3719_ (.A0(_0766_),
    .A1(_0835_),
    .S(_0834_),
    .X(_0836_));
 sg13g2_nand2_1 _3720_ (.Y(_0837_),
    .A(_0718_),
    .B(_0769_));
 sg13g2_xor2_1 _3721_ (.B(_0832_),
    .A(_0831_),
    .X(_0838_));
 sg13g2_o21ai_1 _3722_ (.B1(_0837_),
    .Y(_0839_),
    .A1(_0769_),
    .A2(_0838_));
 sg13g2_nor2b_1 _3723_ (.A(_0839_),
    .B_N(_0836_),
    .Y(_0840_));
 sg13g2_nand3_1 _3724_ (.B(_0830_),
    .C(_0840_),
    .A(_0828_),
    .Y(_0841_));
 sg13g2_xnor2_1 _3725_ (.Y(_0842_),
    .A(net687),
    .B(_0774_));
 sg13g2_o21ai_1 _3726_ (.B1(_0786_),
    .Y(_0843_),
    .A1(net732),
    .A2(_0781_));
 sg13g2_xnor2_1 _3727_ (.Y(_0844_),
    .A(_0842_),
    .B(_0843_));
 sg13g2_mux2_2 _3728_ (.A0(_0774_),
    .A1(_0844_),
    .S(net614),
    .X(_0845_));
 sg13g2_nor2_1 _3729_ (.A(net683),
    .B(_0769_),
    .Y(_0846_));
 sg13g2_xor2_1 _3730_ (.B(net735),
    .A(\core.TauW_q[5] ),
    .X(_0847_));
 sg13g2_xnor2_1 _3731_ (.Y(_0848_),
    .A(_0846_),
    .B(_0847_));
 sg13g2_mux2_1 _3732_ (.A0(_0846_),
    .A1(_0848_),
    .S(net615),
    .X(_0849_));
 sg13g2_nor2_1 _3733_ (.A(_0003_),
    .B(_0849_),
    .Y(_0850_));
 sg13g2_and2_1 _3734_ (.A(net736),
    .B(net615),
    .X(_0851_));
 sg13g2_a21oi_1 _3735_ (.A1(net733),
    .A2(_0851_),
    .Y(_0852_),
    .B1(_0592_));
 sg13g2_a221oi_1 _3736_ (.B2(net733),
    .C1(_0592_),
    .B1(_0851_),
    .A1(_0849_),
    .Y(_0853_),
    .A2(_0003_));
 sg13g2_xnor2_1 _3737_ (.Y(_0854_),
    .A(_0784_),
    .B(_0785_));
 sg13g2_mux2_2 _3738_ (.A0(_0781_),
    .A1(_0854_),
    .S(net614),
    .X(_0855_));
 sg13g2_xnor2_1 _3739_ (.Y(_0856_),
    .A(_1972_),
    .B(_0855_));
 sg13g2_or3_1 _3740_ (.A(_0856_),
    .B(_0853_),
    .C(_0850_),
    .X(_0857_));
 sg13g2_nor2_1 _3741_ (.A(net731),
    .B(_0855_),
    .Y(_0858_));
 sg13g2_nor2_1 _3742_ (.A(net730),
    .B(_0845_),
    .Y(_0859_));
 sg13g2_nor2_1 _3743_ (.A(_0858_),
    .B(_0859_),
    .Y(_0860_));
 sg13g2_and2_1 _3744_ (.A(net730),
    .B(_0845_),
    .X(_0861_));
 sg13g2_a21o_1 _3745_ (.A2(_0860_),
    .A1(_0857_),
    .B1(_0861_),
    .X(_0862_));
 sg13g2_a221oi_1 _3746_ (.B2(_0787_),
    .C1(_0809_),
    .B1(_0786_),
    .A1(net731),
    .Y(_0863_),
    .A2(_0774_));
 sg13g2_nor2_1 _3747_ (.A(_0812_),
    .B(_0863_),
    .Y(_0864_));
 sg13g2_xnor2_1 _3748_ (.Y(_0865_),
    .A(_0800_),
    .B(_0864_));
 sg13g2_mux2_2 _3749_ (.A0(_0796_),
    .A1(_0865_),
    .S(net615),
    .X(_0866_));
 sg13g2_xnor2_1 _3750_ (.Y(_0867_),
    .A(\core.TauW_q[10] ),
    .B(_0866_));
 sg13g2_o21ai_1 _3751_ (.B1(_0809_),
    .Y(_0868_),
    .A1(_0788_),
    .A2(_0789_));
 sg13g2_nor2b_1 _3752_ (.A(_0863_),
    .B_N(_0868_),
    .Y(_0869_));
 sg13g2_mux2_1 _3753_ (.A0(_0806_),
    .A1(_0869_),
    .S(net614),
    .X(_0870_));
 sg13g2_inv_1 _3754_ (.Y(_0871_),
    .A(_0870_));
 sg13g2_xnor2_1 _3755_ (.Y(_0872_),
    .A(_0006_),
    .B(_0870_));
 sg13g2_or2_1 _3756_ (.X(_0873_),
    .B(_0872_),
    .A(_0867_));
 sg13g2_a221oi_1 _3757_ (.B2(_0857_),
    .C1(_0873_),
    .B1(_0860_),
    .A1(net730),
    .Y(_0874_),
    .A2(_0845_));
 sg13g2_nand2_1 _3758_ (.Y(_0875_),
    .A(_1927_),
    .B(_0870_));
 sg13g2_a21o_1 _3759_ (.A2(_0866_),
    .A1(\core.TauW_q[10] ),
    .B1(_0875_),
    .X(_0876_));
 sg13g2_o21ai_1 _3760_ (.B1(_0876_),
    .Y(_0877_),
    .A1(\core.TauW_q[10] ),
    .A2(_0866_));
 sg13g2_or2_1 _3761_ (.X(_0878_),
    .B(_0877_),
    .A(_0874_));
 sg13g2_xor2_1 _3762_ (.B(_0826_),
    .A(_0814_),
    .X(_0879_));
 sg13g2_nand2_1 _3763_ (.Y(_0880_),
    .A(net614),
    .B(_0879_));
 sg13g2_o21ai_1 _3764_ (.B1(_0880_),
    .Y(_0881_),
    .A1(_0825_),
    .A2(net614));
 sg13g2_nand2b_1 _3765_ (.Y(_0882_),
    .B(_1968_),
    .A_N(_0881_));
 sg13g2_o21ai_1 _3766_ (.B1(_0882_),
    .Y(_0883_),
    .A1(_0877_),
    .A2(_0874_));
 sg13g2_nand2_1 _3767_ (.Y(_0884_),
    .A(_0000_),
    .B(_0881_));
 sg13g2_a22oi_1 _3768_ (.Y(_0885_),
    .B1(_0826_),
    .B2(_0814_),
    .A2(_0824_),
    .A1(_1926_));
 sg13g2_xnor2_1 _3769_ (.Y(_0886_),
    .A(_0821_),
    .B(_0885_));
 sg13g2_nand3_1 _3770_ (.B(_0830_),
    .C(_0836_),
    .A(_0828_),
    .Y(_0887_));
 sg13g2_nand2b_1 _3771_ (.Y(_0888_),
    .B(_0887_),
    .A_N(_0840_));
 sg13g2_nor2_1 _3772_ (.A(_0819_),
    .B(net614),
    .Y(_0889_));
 sg13g2_a21oi_1 _3773_ (.A1(net614),
    .A2(_0886_),
    .Y(_0890_),
    .B1(_0889_));
 sg13g2_nand2_1 _3774_ (.Y(_0891_),
    .A(_0884_),
    .B(_0888_));
 sg13g2_nor2_2 _3775_ (.A(_0890_),
    .B(_0891_),
    .Y(_0892_));
 sg13g2_nand2_2 _3776_ (.Y(_0893_),
    .A(_0892_),
    .B(_0883_));
 sg13g2_or2_1 _3777_ (.X(_0894_),
    .B(_0861_),
    .A(_0859_));
 sg13g2_o21ai_1 _3778_ (.B1(_0857_),
    .Y(_0895_),
    .A1(net731),
    .A2(_0855_));
 sg13g2_xor2_1 _3779_ (.B(_0895_),
    .A(_0894_),
    .X(_0896_));
 sg13g2_mux2_1 _3780_ (.A0(_0845_),
    .A1(_0896_),
    .S(_0893_),
    .X(_0897_));
 sg13g2_xor2_1 _3781_ (.B(_0897_),
    .A(_0006_),
    .X(_0898_));
 sg13g2_o21ai_1 _3782_ (.B1(_0856_),
    .Y(_0899_),
    .A1(_0850_),
    .A2(_0853_));
 sg13g2_nand2_1 _3783_ (.Y(_0900_),
    .A(_0857_),
    .B(_0899_));
 sg13g2_mux2_1 _3784_ (.A0(_0855_),
    .A1(_0900_),
    .S(_0893_),
    .X(_0901_));
 sg13g2_nand2_1 _3785_ (.Y(_0902_),
    .A(_1973_),
    .B(_0901_));
 sg13g2_xnor2_1 _3786_ (.Y(_0903_),
    .A(_1973_),
    .B(_0901_));
 sg13g2_nor2_2 _3787_ (.A(_0903_),
    .B(_0898_),
    .Y(_0904_));
 sg13g2_xor2_1 _3788_ (.B(_0851_),
    .A(_0847_),
    .X(_0905_));
 sg13g2_and3_1 _3789_ (.X(_0906_),
    .A(_0851_),
    .B(_0883_),
    .C(_0892_));
 sg13g2_a21oi_1 _3790_ (.A1(_0883_),
    .A2(_0892_),
    .Y(_0907_),
    .B1(_0905_));
 sg13g2_or3_1 _3791_ (.A(_0003_),
    .B(_0906_),
    .C(_0907_),
    .X(_0908_));
 sg13g2_o21ai_1 _3792_ (.B1(_0003_),
    .Y(_0909_),
    .A1(_0906_),
    .A2(_0907_));
 sg13g2_nand3b_1 _3793_ (.B(_0883_),
    .C(_0892_),
    .Y(_0910_),
    .A_N(_0849_));
 sg13g2_xnor2_1 _3794_ (.Y(_0911_),
    .A(_0003_),
    .B(_0849_));
 sg13g2_xor2_1 _3795_ (.B(_0911_),
    .A(_0852_),
    .X(_0912_));
 sg13g2_a21o_1 _3796_ (.A2(_0892_),
    .A1(_0883_),
    .B1(_0912_),
    .X(_0913_));
 sg13g2_nand3_1 _3797_ (.B(_0910_),
    .C(_0913_),
    .A(net687),
    .Y(_0914_));
 sg13g2_a21oi_1 _3798_ (.A1(_0910_),
    .A2(_0913_),
    .Y(_0915_),
    .B1(net687));
 sg13g2_a21o_1 _3799_ (.A2(_0913_),
    .A1(_0910_),
    .B1(net687),
    .X(_0916_));
 sg13g2_nand4_1 _3800_ (.B(_0909_),
    .C(_0914_),
    .A(_0908_),
    .Y(_0917_),
    .D(_0916_));
 sg13g2_a21oi_1 _3801_ (.A1(_0883_),
    .A2(_0892_),
    .Y(_0918_),
    .B1(net683));
 sg13g2_nand2_1 _3802_ (.Y(_0919_),
    .A(net684),
    .B(_0918_));
 sg13g2_o21ai_1 _3803_ (.B1(net733),
    .Y(_0920_),
    .A1(\core.TauW_q[5] ),
    .A2(net683));
 sg13g2_o21ai_1 _3804_ (.B1(_0919_),
    .Y(_0921_),
    .A1(_0918_),
    .A2(_0920_));
 sg13g2_nor3_1 _3805_ (.A(net685),
    .B(_0906_),
    .C(_0907_),
    .Y(_0922_));
 sg13g2_o21ai_1 _3806_ (.B1(_0914_),
    .Y(_0923_),
    .A1(_0915_),
    .A2(_0922_));
 sg13g2_o21ai_1 _3807_ (.B1(_0923_),
    .Y(_0924_),
    .A1(_0917_),
    .A2(_0921_));
 sg13g2_nor2_1 _3808_ (.A(_0898_),
    .B(_0902_),
    .Y(_0925_));
 sg13g2_a221oi_1 _3809_ (.B2(_0904_),
    .C1(_0925_),
    .B1(_0924_),
    .A1(\core.TauW_q[9] ),
    .Y(_0926_),
    .A2(_0897_));
 sg13g2_xnor2_1 _3810_ (.Y(_0927_),
    .A(_0862_),
    .B(_0872_));
 sg13g2_mux2_1 _3811_ (.A0(_0871_),
    .A1(_0927_),
    .S(_0893_),
    .X(_0928_));
 sg13g2_xor2_1 _3812_ (.B(_0928_),
    .A(_0007_),
    .X(_0929_));
 sg13g2_nand2_1 _3813_ (.Y(_0930_),
    .A(\core.TauW_q[10] ),
    .B(_0928_));
 sg13g2_o21ai_1 _3814_ (.B1(_0930_),
    .Y(_0931_),
    .A1(_0929_),
    .A2(_0926_));
 sg13g2_nor2_1 _3815_ (.A(_0866_),
    .B(_0893_),
    .Y(_0932_));
 sg13g2_o21ai_1 _3816_ (.B1(_0875_),
    .Y(_0933_),
    .A1(_0862_),
    .A2(_0872_));
 sg13g2_xnor2_1 _3817_ (.Y(_0934_),
    .A(_0867_),
    .B(_0933_));
 sg13g2_a21oi_1 _3818_ (.A1(_0893_),
    .A2(_0934_),
    .Y(_0935_),
    .B1(_0932_));
 sg13g2_nor2_1 _3819_ (.A(\core.TauW_q[11] ),
    .B(_0935_),
    .Y(_0936_));
 sg13g2_nor4_1 _3820_ (.A(_0593_),
    .B(_0898_),
    .C(_0903_),
    .D(_0929_),
    .Y(_0937_));
 sg13g2_nor2b_1 _3821_ (.A(_0917_),
    .B_N(_0937_),
    .Y(_0938_));
 sg13g2_nor2_1 _3822_ (.A(_0936_),
    .B(_0938_),
    .Y(_0939_));
 sg13g2_a22oi_1 _3823_ (.Y(_0940_),
    .B1(_0931_),
    .B2(_0939_),
    .A2(_0935_),
    .A1(\core.TauW_q[11] ));
 sg13g2_xnor2_1 _3824_ (.Y(_0941_),
    .A(_0000_),
    .B(_0878_));
 sg13g2_nand2_1 _3825_ (.Y(_0942_),
    .A(_0881_),
    .B(_0941_));
 sg13g2_o21ai_1 _3826_ (.B1(_0890_),
    .Y(_0943_),
    .A1(_0000_),
    .A2(_0878_));
 sg13g2_nand3_1 _3827_ (.B(_0942_),
    .C(_0943_),
    .A(_0888_),
    .Y(_0944_));
 sg13g2_nor2_1 _3828_ (.A(_0940_),
    .B(_0944_),
    .Y(_0945_));
 sg13g2_o21ai_1 _3829_ (.B1(net681),
    .Y(_0946_),
    .A1(_0516_),
    .A2(_0593_));
 sg13g2_nand2_1 _3830_ (.Y(_0947_),
    .A(net472),
    .B(net770));
 sg13g2_o21ai_1 _3831_ (.B1(_0947_),
    .Y(_0063_),
    .A1(_0945_),
    .A2(net646));
 sg13g2_nand2_1 _3832_ (.Y(_0948_),
    .A(net498),
    .B(net767));
 sg13g2_nor2_1 _3833_ (.A(net628),
    .B(_0945_),
    .Y(_0949_));
 sg13g2_xnor2_1 _3834_ (.Y(_0950_),
    .A(_0893_),
    .B(_0949_));
 sg13g2_o21ai_1 _3835_ (.B1(_0948_),
    .Y(_0064_),
    .A1(net646),
    .A2(_0950_));
 sg13g2_nor3_1 _3836_ (.A(_0893_),
    .B(_0940_),
    .C(_0944_),
    .Y(_0951_));
 sg13g2_nor2_2 _3837_ (.A(net628),
    .B(_0951_),
    .Y(_0952_));
 sg13g2_xnor2_1 _3838_ (.Y(_0953_),
    .A(net615),
    .B(_0952_));
 sg13g2_nand2_1 _3839_ (.Y(_0954_),
    .A(net542),
    .B(net767));
 sg13g2_o21ai_1 _3840_ (.B1(_0954_),
    .Y(_0065_),
    .A1(net646),
    .A2(_0953_));
 sg13g2_a21oi_1 _3841_ (.A1(net627),
    .A2(net615),
    .Y(_0955_),
    .B1(_0952_));
 sg13g2_xnor2_1 _3842_ (.Y(_0956_),
    .A(_0769_),
    .B(_0955_));
 sg13g2_nand2_1 _3843_ (.Y(_0957_),
    .A(net559),
    .B(net767));
 sg13g2_o21ai_1 _3844_ (.B1(_0957_),
    .Y(_0066_),
    .A1(net646),
    .A2(_0956_));
 sg13g2_nand2_1 _3845_ (.Y(_0958_),
    .A(net505),
    .B(net768));
 sg13g2_or2_1 _3846_ (.X(_0959_),
    .B(net614),
    .A(_0770_));
 sg13g2_nor4_2 _3847_ (.A(_0893_),
    .B(_0959_),
    .C(_0944_),
    .Y(_0960_),
    .D(_0940_));
 sg13g2_nor2_1 _3848_ (.A(net282),
    .B(_0960_),
    .Y(_0961_));
 sg13g2_xnor2_1 _3849_ (.Y(_0962_),
    .A(_0710_),
    .B(_0961_));
 sg13g2_o21ai_1 _3850_ (.B1(_0958_),
    .Y(_0067_),
    .A1(net645),
    .A2(_0962_));
 sg13g2_a21oi_1 _3851_ (.A1(net627),
    .A2(_0710_),
    .Y(_0963_),
    .B1(_0961_));
 sg13g2_xor2_1 _3852_ (.B(_0963_),
    .A(net622),
    .X(_0964_));
 sg13g2_nand2_1 _3853_ (.Y(_0965_),
    .A(net593),
    .B(net769));
 sg13g2_o21ai_1 _3854_ (.B1(_0965_),
    .Y(_0068_),
    .A1(net645),
    .A2(_0964_));
 sg13g2_nor2_1 _3855_ (.A(net621),
    .B(_0710_),
    .Y(_0966_));
 sg13g2_and2_1 _3856_ (.A(_0966_),
    .B(_0960_),
    .X(_0967_));
 sg13g2_nor2_1 _3857_ (.A(net283),
    .B(_0967_),
    .Y(_0968_));
 sg13g2_xnor2_1 _3858_ (.Y(_0969_),
    .A(_0620_),
    .B(_0968_));
 sg13g2_nand2_1 _3859_ (.Y(_0970_),
    .A(net539),
    .B(net769));
 sg13g2_o21ai_1 _3860_ (.B1(_0970_),
    .Y(_0069_),
    .A1(net645),
    .A2(_0969_));
 sg13g2_nand2_1 _3861_ (.Y(_0971_),
    .A(net556),
    .B(net768));
 sg13g2_a21oi_2 _3862_ (.B1(net282),
    .Y(_0972_),
    .A2(_0967_),
    .A1(_0619_));
 sg13g2_xnor2_1 _3863_ (.Y(_0973_),
    .A(_0972_),
    .B(net626));
 sg13g2_o21ai_1 _3864_ (.B1(_0971_),
    .Y(_0070_),
    .A1(net645),
    .A2(_0973_));
 sg13g2_nand2_1 _3865_ (.Y(_0974_),
    .A(net581),
    .B(net768));
 sg13g2_nor4_1 _3866_ (.A(_0585_),
    .B(_0620_),
    .C(net621),
    .D(_0710_),
    .Y(_0975_));
 sg13g2_a21oi_2 _3867_ (.B1(net628),
    .Y(_0976_),
    .A2(_0960_),
    .A1(_0975_));
 sg13g2_xnor2_1 _3868_ (.Y(_0977_),
    .A(_0555_),
    .B(_0976_));
 sg13g2_o21ai_1 _3869_ (.B1(_0974_),
    .Y(_0071_),
    .A1(net645),
    .A2(_0977_));
 sg13g2_a21o_1 _3870_ (.A2(_0555_),
    .A1(net627),
    .B1(_0976_),
    .X(_0978_));
 sg13g2_xnor2_1 _3871_ (.Y(_0979_),
    .A(_0532_),
    .B(_0978_));
 sg13g2_nand2_1 _3872_ (.Y(_0980_),
    .A(net605),
    .B(net768));
 sg13g2_o21ai_1 _3873_ (.B1(_0980_),
    .Y(_0072_),
    .A1(net646),
    .A2(_0979_));
 sg13g2_nand2_1 _3874_ (.Y(_0981_),
    .A(net514),
    .B(net768));
 sg13g2_o21ai_1 _3875_ (.B1(net627),
    .Y(_0982_),
    .A1(_0532_),
    .A2(_0555_));
 sg13g2_nor2b_2 _3876_ (.A(_0976_),
    .B_N(_0982_),
    .Y(_0983_));
 sg13g2_xnor2_1 _3877_ (.Y(_0984_),
    .A(_0518_),
    .B(_0983_));
 sg13g2_o21ai_1 _3878_ (.B1(_0981_),
    .Y(_0073_),
    .A1(net645),
    .A2(_0984_));
 sg13g2_o21ai_1 _3879_ (.B1(_0983_),
    .Y(_0985_),
    .A1(net628),
    .A2(_0518_));
 sg13g2_nor2_1 _3880_ (.A(net737),
    .B(_0501_),
    .Y(_0986_));
 sg13g2_nand2b_1 _3881_ (.Y(_0987_),
    .B(net683),
    .A_N(_0501_));
 sg13g2_or4_1 _3882_ (.A(net628),
    .B(_0496_),
    .C(_0498_),
    .D(_0501_),
    .X(_0988_));
 sg13g2_a22oi_1 _3883_ (.Y(_0989_),
    .B1(_0987_),
    .B2(_0988_),
    .A2(net287),
    .A1(_1969_));
 sg13g2_xnor2_1 _3884_ (.Y(_0990_),
    .A(_0985_),
    .B(_0989_));
 sg13g2_nand2_1 _3885_ (.Y(_0991_),
    .A(net469),
    .B(net768));
 sg13g2_o21ai_1 _3886_ (.B1(_0991_),
    .Y(_0074_),
    .A1(_0990_),
    .A2(net645));
 sg13g2_nor2_1 _3887_ (.A(net628),
    .B(net646),
    .Y(_0992_));
 sg13g2_a21o_1 _3888_ (.A2(net768),
    .A1(net817),
    .B1(_0992_),
    .X(_0075_));
 sg13g2_a21oi_1 _3889_ (.A1(net284),
    .A2(_0986_),
    .Y(_0993_),
    .B1(net645));
 sg13g2_o21ai_1 _3890_ (.B1(_0993_),
    .Y(_0994_),
    .A1(net627),
    .A2(_0986_));
 sg13g2_o21ai_1 _3891_ (.B1(_0994_),
    .Y(_0076_),
    .A1(_1977_),
    .A2(_2139_));
 sg13g2_a21o_1 _3892_ (.A2(net768),
    .A1(net578),
    .B1(_0992_),
    .X(_0077_));
 sg13g2_o21ai_1 _3893_ (.B1(_0994_),
    .Y(_0078_),
    .A1(_1979_),
    .A2(_2139_));
 sg13g2_nor2_2 _3894_ (.A(\core.drive[0] ),
    .B(\core.drive[1] ),
    .Y(_0995_));
 sg13g2_and3_1 _3895_ (.X(_0996_),
    .A(_0023_),
    .B(net760),
    .C(_0995_));
 sg13g2_nor2_1 _3896_ (.A(\core.C_q[10] ),
    .B(\core.C_q[9] ),
    .Y(_0997_));
 sg13g2_nand4_1 _3897_ (.B(_1953_),
    .C(_0025_),
    .A(_1952_),
    .Y(_0998_),
    .D(_0997_));
 sg13g2_or3_1 _3898_ (.A(\core.C_q[6] ),
    .B(net756),
    .C(_0998_),
    .X(_0999_));
 sg13g2_o21ai_1 _3899_ (.B1(_0996_),
    .Y(_1000_),
    .A1(_0026_),
    .A2(_0999_));
 sg13g2_nor2_1 _3900_ (.A(\core.C_q[11] ),
    .B(\core.C_q[10] ),
    .Y(_1001_));
 sg13g2_nand3_1 _3901_ (.B(_1952_),
    .C(_1001_),
    .A(_1951_),
    .Y(_1002_));
 sg13g2_nor3_2 _3902_ (.A(net337),
    .B(\core.C_q[6] ),
    .C(_1002_),
    .Y(_1003_));
 sg13g2_nor2_2 _3903_ (.A(_0023_),
    .B(net760),
    .Y(_1004_));
 sg13g2_xnor2_1 _3904_ (.Y(_1005_),
    .A(\core.drive[2] ),
    .B(_0995_));
 sg13g2_a21oi_2 _3905_ (.B1(_1004_),
    .Y(_1006_),
    .A2(_1005_),
    .A1(net760));
 sg13g2_xnor2_1 _3906_ (.Y(_1007_),
    .A(_1006_),
    .B(net757));
 sg13g2_nor2_1 _3907_ (.A(net759),
    .B(_1006_),
    .Y(_1008_));
 sg13g2_nor3_2 _3908_ (.A(net754),
    .B(_1007_),
    .C(_1008_),
    .Y(_1009_));
 sg13g2_nor2b_2 _3909_ (.A(_1009_),
    .B_N(_1003_),
    .Y(_1010_));
 sg13g2_o21ai_1 _3910_ (.B1(net754),
    .Y(_1011_),
    .A1(_1008_),
    .A2(_1007_));
 sg13g2_a21oi_1 _3911_ (.A1(_1010_),
    .A2(net335),
    .Y(_1012_),
    .B1(_1000_));
 sg13g2_nand2_2 _3912_ (.Y(_1013_),
    .A(_1011_),
    .B(_1000_));
 sg13g2_nand2_1 _3913_ (.Y(_1014_),
    .A(_1010_),
    .B(_1013_));
 sg13g2_nand3b_1 _3914_ (.B(_1013_),
    .C(_1010_),
    .Y(_1015_),
    .A_N(net334));
 sg13g2_a21o_1 _3915_ (.A2(_1010_),
    .A1(_1013_),
    .B1(_1006_),
    .X(_1016_));
 sg13g2_and2_1 _3916_ (.A(_1015_),
    .B(_1016_),
    .X(_1017_));
 sg13g2_nor2_1 _3917_ (.A(net756),
    .B(_1017_),
    .Y(_1018_));
 sg13g2_nand2_1 _3918_ (.Y(_1019_),
    .A(net345),
    .B(\core.drive[1] ));
 sg13g2_nand3b_1 _3919_ (.B(_1019_),
    .C(net762),
    .Y(_1020_),
    .A_N(_0995_));
 sg13g2_o21ai_1 _3920_ (.B1(_1020_),
    .Y(_1021_),
    .A1(net762),
    .A2(_0024_));
 sg13g2_nor2_1 _3921_ (.A(net757),
    .B(_1021_),
    .Y(_1022_));
 sg13g2_nand3_1 _3922_ (.B(_1015_),
    .C(net753),
    .A(_1016_),
    .Y(_1023_));
 sg13g2_a21o_1 _3923_ (.A2(_1015_),
    .A1(_1016_),
    .B1(net753),
    .X(_1024_));
 sg13g2_nand2_1 _3924_ (.Y(_1025_),
    .A(_1023_),
    .B(_1024_));
 sg13g2_a21oi_2 _3925_ (.B1(_1022_),
    .Y(_1026_),
    .A2(_1023_),
    .A1(_1024_));
 sg13g2_nor2_2 _3926_ (.A(_1018_),
    .B(_1026_),
    .Y(_1027_));
 sg13g2_a21o_1 _3927_ (.A2(net682),
    .A1(_1027_),
    .B1(_0998_),
    .X(_1028_));
 sg13g2_nor2_1 _3928_ (.A(net682),
    .B(_1027_),
    .Y(_1029_));
 sg13g2_o21ai_1 _3929_ (.B1(net752),
    .Y(_1030_),
    .A1(_1018_),
    .A2(_1026_));
 sg13g2_o21ai_1 _3930_ (.B1(_1012_),
    .Y(_1031_),
    .A1(_1028_),
    .A2(_1029_));
 sg13g2_nor2b_2 _3931_ (.A(_1012_),
    .B_N(_1030_),
    .Y(_1032_));
 sg13g2_or2_1 _3932_ (.X(_1033_),
    .B(_1032_),
    .A(_1028_));
 sg13g2_inv_1 _3933_ (.Y(_1034_),
    .A(_1033_));
 sg13g2_nor3_2 _3934_ (.A(_0026_),
    .B(_1032_),
    .C(_1028_),
    .Y(_1035_));
 sg13g2_xor2_1 _3935_ (.B(_1035_),
    .A(_1021_),
    .X(_1036_));
 sg13g2_nand2_1 _3936_ (.Y(_1037_),
    .A(net753),
    .B(_1036_));
 sg13g2_nor2_1 _3937_ (.A(_1955_),
    .B(net343),
    .Y(_1038_));
 sg13g2_xnor2_1 _3938_ (.Y(_1039_),
    .A(_1036_),
    .B(net753));
 sg13g2_o21ai_1 _3939_ (.B1(_1037_),
    .Y(_1040_),
    .A1(_1039_),
    .A2(_1038_));
 sg13g2_xnor2_1 _3940_ (.Y(_1041_),
    .A(_1022_),
    .B(_1025_));
 sg13g2_nand2b_1 _3941_ (.Y(_1042_),
    .B(_1041_),
    .A_N(_1033_));
 sg13g2_o21ai_1 _3942_ (.B1(_1042_),
    .Y(_1043_),
    .A1(_1034_),
    .A2(_1017_));
 sg13g2_xnor2_1 _3943_ (.Y(_1044_),
    .A(_1043_),
    .B(net682));
 sg13g2_a22oi_1 _3944_ (.Y(_1045_),
    .B1(_1040_),
    .B2(_1044_),
    .A2(_1043_),
    .A1(_1954_));
 sg13g2_a21oi_2 _3945_ (.B1(_1002_),
    .Y(_1046_),
    .A2(_1045_),
    .A1(_1966_));
 sg13g2_nand2b_1 _3946_ (.Y(_1047_),
    .B(_0022_),
    .A_N(_1045_));
 sg13g2_a21oi_1 _3947_ (.A1(_1046_),
    .A2(_1047_),
    .Y(_1048_),
    .B1(_1031_));
 sg13g2_o21ai_1 _3948_ (.B1(_1031_),
    .Y(_1049_),
    .A1(_1045_),
    .A2(_1966_));
 sg13g2_nand2_2 _3949_ (.Y(_1050_),
    .A(_1049_),
    .B(_1046_));
 sg13g2_inv_1 _3950_ (.Y(_1051_),
    .A(_1050_));
 sg13g2_a21o_1 _3951_ (.A2(_1049_),
    .A1(_1046_),
    .B1(_1967_),
    .X(_1052_));
 sg13g2_xnor2_1 _3952_ (.Y(_1053_),
    .A(net758),
    .B(net343));
 sg13g2_nand3_1 _3953_ (.B(_1053_),
    .C(_1049_),
    .A(_1046_),
    .Y(_1054_));
 sg13g2_nand2_1 _3954_ (.Y(_1055_),
    .A(_1052_),
    .B(_1054_));
 sg13g2_or2_1 _3955_ (.X(_1056_),
    .B(_1055_),
    .A(net755));
 sg13g2_a21oi_1 _3956_ (.A1(_1052_),
    .A2(_1054_),
    .Y(_1057_),
    .B1(_1964_));
 sg13g2_and3_1 _3957_ (.X(_1058_),
    .A(_1054_),
    .B(_1052_),
    .C(_1964_));
 sg13g2_nor2_1 _3958_ (.A(_1057_),
    .B(_1058_),
    .Y(_1059_));
 sg13g2_o21ai_1 _3959_ (.B1(_1955_),
    .Y(_1060_),
    .A1(_1057_),
    .A2(_1058_));
 sg13g2_xor2_1 _3960_ (.B(net333),
    .A(_1038_),
    .X(_1061_));
 sg13g2_mux2_2 _3961_ (.A0(_1061_),
    .A1(_1036_),
    .S(_1050_),
    .X(_1062_));
 sg13g2_xnor2_1 _3962_ (.Y(_1063_),
    .A(net682),
    .B(_1062_));
 sg13g2_xnor2_1 _3963_ (.Y(_1064_),
    .A(_1062_),
    .B(net752));
 sg13g2_a21oi_2 _3964_ (.B1(_1064_),
    .Y(_1065_),
    .A2(_1060_),
    .A1(_1056_));
 sg13g2_and2_1 _3965_ (.A(_1954_),
    .B(_1062_),
    .X(_1066_));
 sg13g2_nand2_1 _3966_ (.Y(_1067_),
    .A(_1043_),
    .B(_1050_));
 sg13g2_xnor2_1 _3967_ (.Y(_1068_),
    .A(net332),
    .B(_1044_));
 sg13g2_o21ai_1 _3968_ (.B1(_1067_),
    .Y(_1069_),
    .A1(_1050_),
    .A2(_1068_));
 sg13g2_xnor2_1 _3969_ (.Y(_1070_),
    .A(_1966_),
    .B(_1069_));
 sg13g2_inv_1 _3970_ (.Y(_1071_),
    .A(_1070_));
 sg13g2_o21ai_1 _3971_ (.B1(_1070_),
    .Y(_1072_),
    .A1(_1066_),
    .A2(_1065_));
 sg13g2_nand2_1 _3972_ (.Y(_1073_),
    .A(net751),
    .B(_1048_));
 sg13g2_nand2_1 _3973_ (.Y(_1074_),
    .A(_1953_),
    .B(_1069_));
 sg13g2_and2_1 _3974_ (.A(_1073_),
    .B(_1074_),
    .X(_1075_));
 sg13g2_or2_1 _3975_ (.X(_1076_),
    .B(_1048_),
    .A(net751));
 sg13g2_nand3_1 _3976_ (.B(_0997_),
    .C(_1076_),
    .A(_0025_),
    .Y(_1077_));
 sg13g2_a21o_2 _3977_ (.A2(_1072_),
    .A1(_1075_),
    .B1(_1077_),
    .X(_1078_));
 sg13g2_inv_2 _3978_ (.Y(_1079_),
    .A(_1078_));
 sg13g2_nand2_1 _3979_ (.Y(_1080_),
    .A(_1073_),
    .B(_1076_));
 sg13g2_o21ai_1 _3980_ (.B1(_1056_),
    .Y(_1081_),
    .A1(_1963_),
    .A2(_1059_));
 sg13g2_a21oi_1 _3981_ (.A1(_1063_),
    .A2(_1081_),
    .Y(_1082_),
    .B1(_1066_));
 sg13g2_o21ai_1 _3982_ (.B1(_1074_),
    .Y(_1083_),
    .A1(_1071_),
    .A2(_1082_));
 sg13g2_xnor2_1 _3983_ (.Y(_1084_),
    .A(_1080_),
    .B(_1083_));
 sg13g2_mux2_1 _3984_ (.A0(_1048_),
    .A1(_1084_),
    .S(_1079_),
    .X(_1085_));
 sg13g2_nand2_1 _3985_ (.Y(_1086_),
    .A(_1062_),
    .B(_1078_));
 sg13g2_xnor2_1 _3986_ (.Y(_1087_),
    .A(_1063_),
    .B(_1081_));
 sg13g2_o21ai_1 _3987_ (.B1(_1086_),
    .Y(_1088_),
    .A1(_1078_),
    .A2(_1087_));
 sg13g2_nor2_2 _3988_ (.A(net756),
    .B(net759),
    .Y(_1089_));
 sg13g2_a21oi_1 _3989_ (.A1(net759),
    .A2(_1078_),
    .Y(_1090_),
    .B1(net756));
 sg13g2_xnor2_1 _3990_ (.Y(_1091_),
    .A(_1963_),
    .B(_1059_));
 sg13g2_mux2_1 _3991_ (.A0(_1091_),
    .A1(_1055_),
    .S(_1078_),
    .X(_1092_));
 sg13g2_inv_1 _3992_ (.Y(_1093_),
    .A(_1092_));
 sg13g2_xnor2_1 _3993_ (.Y(_1094_),
    .A(_1092_),
    .B(net752));
 sg13g2_nor2_1 _3994_ (.A(\core.C_q[6] ),
    .B(_1092_),
    .Y(_1095_));
 sg13g2_a21o_1 _3995_ (.A2(_1090_),
    .A1(_1094_),
    .B1(_1095_),
    .X(_1096_));
 sg13g2_xnor2_1 _3996_ (.Y(_1097_),
    .A(_1966_),
    .B(_1088_));
 sg13g2_a22oi_1 _3997_ (.Y(_1098_),
    .B1(_1096_),
    .B2(_1097_),
    .A2(_1088_),
    .A1(_1953_));
 sg13g2_xnor2_1 _3998_ (.Y(_1099_),
    .A(_1071_),
    .B(_1082_));
 sg13g2_nand2_1 _3999_ (.Y(_1100_),
    .A(_1069_),
    .B(_1078_));
 sg13g2_o21ai_1 _4000_ (.B1(_1100_),
    .Y(_1101_),
    .A1(_1078_),
    .A2(_1099_));
 sg13g2_xnor2_1 _4001_ (.Y(_1102_),
    .A(_0029_),
    .B(_1101_));
 sg13g2_nand2_1 _4002_ (.Y(_1103_),
    .A(_1952_),
    .B(_1101_));
 sg13g2_o21ai_1 _4003_ (.B1(_1103_),
    .Y(_1104_),
    .A1(_1102_),
    .A2(_1098_));
 sg13g2_o21ai_1 _4004_ (.B1(_1001_),
    .Y(_1105_),
    .A1(_1104_),
    .A2(net750));
 sg13g2_and2_1 _4005_ (.A(net750),
    .B(_1104_),
    .X(_1106_));
 sg13g2_o21ai_1 _4006_ (.B1(_1085_),
    .Y(_1107_),
    .A1(_1105_),
    .A2(_1106_));
 sg13g2_a21oi_2 _4007_ (.B1(_1085_),
    .Y(_1108_),
    .A2(_1104_),
    .A1(net750));
 sg13g2_nor2_2 _4008_ (.A(_1108_),
    .B(_1105_),
    .Y(_1109_));
 sg13g2_inv_2 _4009_ (.Y(_1110_),
    .A(_1109_));
 sg13g2_xnor2_1 _4010_ (.Y(_1111_),
    .A(_1098_),
    .B(_1102_));
 sg13g2_nor2_1 _4011_ (.A(_1101_),
    .B(_1109_),
    .Y(_1112_));
 sg13g2_a21oi_2 _4012_ (.B1(_1112_),
    .Y(_1113_),
    .A2(_1111_),
    .A1(_1109_));
 sg13g2_and2_1 _4013_ (.A(_1951_),
    .B(_1113_),
    .X(_1114_));
 sg13g2_nand2_1 _4014_ (.Y(_1115_),
    .A(net759),
    .B(_1079_));
 sg13g2_nand2b_1 _4015_ (.Y(_1116_),
    .B(net757),
    .A_N(net755));
 sg13g2_xnor2_1 _4016_ (.Y(_1117_),
    .A(net755),
    .B(net757));
 sg13g2_xor2_1 _4017_ (.B(net757),
    .A(net755),
    .X(_1118_));
 sg13g2_nor3_2 _4018_ (.A(_1108_),
    .B(_1105_),
    .C(_1118_),
    .Y(_1119_));
 sg13g2_xnor2_1 _4019_ (.Y(_1120_),
    .A(_1119_),
    .B(_1115_));
 sg13g2_nor2_1 _4020_ (.A(_0028_),
    .B(_1120_),
    .Y(_1121_));
 sg13g2_nor3_2 _4021_ (.A(_1955_),
    .B(_1105_),
    .C(_1108_),
    .Y(_1122_));
 sg13g2_a21oi_1 _4022_ (.A1(net754),
    .A2(_1122_),
    .Y(_1123_),
    .B1(_1089_));
 sg13g2_a221oi_1 _4023_ (.B2(net754),
    .C1(_1089_),
    .B1(_1122_),
    .A1(_1120_),
    .Y(_1124_),
    .A2(net752));
 sg13g2_xor2_1 _4024_ (.B(_1094_),
    .A(_1090_),
    .X(_1125_));
 sg13g2_mux2_1 _4025_ (.A0(_1093_),
    .A1(_1125_),
    .S(_1109_),
    .X(_1126_));
 sg13g2_xnor2_1 _4026_ (.Y(_1127_),
    .A(_0022_),
    .B(_1126_));
 sg13g2_nor3_2 _4027_ (.A(_1121_),
    .B(_1127_),
    .C(_1124_),
    .Y(_1128_));
 sg13g2_and2_1 _4028_ (.A(_1953_),
    .B(_1126_),
    .X(_1129_));
 sg13g2_xnor2_1 _4029_ (.Y(_1130_),
    .A(_1096_),
    .B(_1097_));
 sg13g2_nor3_1 _4030_ (.A(_1105_),
    .B(_1108_),
    .C(_1130_),
    .Y(_1131_));
 sg13g2_a21oi_2 _4031_ (.B1(_1131_),
    .Y(_1132_),
    .A2(_1110_),
    .A1(_1088_));
 sg13g2_xnor2_1 _4032_ (.Y(_1133_),
    .A(_0029_),
    .B(_1132_));
 sg13g2_o21ai_1 _4033_ (.B1(_1133_),
    .Y(_1134_),
    .A1(_1129_),
    .A2(_1128_));
 sg13g2_or2_1 _4034_ (.X(_1135_),
    .B(_1132_),
    .A(\core.C_q[8] ));
 sg13g2_xor2_1 _4035_ (.B(_1113_),
    .A(_0030_),
    .X(_1136_));
 sg13g2_inv_1 _4036_ (.Y(_1137_),
    .A(_1136_));
 sg13g2_a21oi_2 _4037_ (.B1(_1137_),
    .Y(_1138_),
    .A2(_1134_),
    .A1(_1135_));
 sg13g2_nor3_1 _4038_ (.A(_0031_),
    .B(_1114_),
    .C(_1138_),
    .Y(_1139_));
 sg13g2_nor2_2 _4039_ (.A(_1962_),
    .B(_1139_),
    .Y(_1140_));
 sg13g2_o21ai_1 _4040_ (.B1(_0031_),
    .Y(_1141_),
    .A1(_1138_),
    .A2(_1114_));
 sg13g2_a21oi_2 _4041_ (.B1(_1107_),
    .Y(_1142_),
    .A2(_1141_),
    .A1(_1140_));
 sg13g2_nand2_2 _4042_ (.Y(_1143_),
    .A(_1107_),
    .B(_1141_));
 sg13g2_nand2_2 _4043_ (.Y(_1144_),
    .A(_1140_),
    .B(_1143_));
 sg13g2_inv_1 _4044_ (.Y(_1145_),
    .A(net625));
 sg13g2_nand3_1 _4045_ (.B(_1140_),
    .C(_1143_),
    .A(_1117_),
    .Y(_1146_));
 sg13g2_xnor2_1 _4046_ (.Y(_1147_),
    .A(_1122_),
    .B(_1146_));
 sg13g2_xnor2_1 _4047_ (.Y(_1148_),
    .A(_1965_),
    .B(_1147_));
 sg13g2_a21oi_1 _4048_ (.A1(net759),
    .A2(_1144_),
    .Y(_1149_),
    .B1(net756));
 sg13g2_a22oi_1 _4049_ (.Y(_1150_),
    .B1(_1148_),
    .B2(_1149_),
    .A2(_1147_),
    .A1(_1954_));
 sg13g2_xnor2_1 _4050_ (.Y(_1151_),
    .A(_1965_),
    .B(_1120_));
 sg13g2_xnor2_1 _4051_ (.Y(_1152_),
    .A(_1123_),
    .B(_1151_));
 sg13g2_mux2_2 _4052_ (.A0(_1152_),
    .A1(_1120_),
    .S(net625),
    .X(_1153_));
 sg13g2_xnor2_1 _4053_ (.Y(_1154_),
    .A(net336),
    .B(_1153_));
 sg13g2_inv_2 _4054_ (.Y(_1155_),
    .A(_1154_));
 sg13g2_nand2_1 _4055_ (.Y(_1156_),
    .A(_0022_),
    .B(_1153_));
 sg13g2_o21ai_1 _4056_ (.B1(_1156_),
    .Y(_1157_),
    .A1(_1155_),
    .A2(_1150_));
 sg13g2_o21ai_1 _4057_ (.B1(_1127_),
    .Y(_1158_),
    .A1(_1121_),
    .A2(_1124_));
 sg13g2_nor2b_1 _4058_ (.A(_1128_),
    .B_N(_1158_),
    .Y(_1159_));
 sg13g2_mux2_2 _4059_ (.A0(_1159_),
    .A1(_1126_),
    .S(net625),
    .X(_1160_));
 sg13g2_xor2_1 _4060_ (.B(_1160_),
    .A(_0029_),
    .X(_1161_));
 sg13g2_a22oi_1 _4061_ (.Y(_1162_),
    .B1(_1157_),
    .B2(_1161_),
    .A2(_1160_),
    .A1(_1952_));
 sg13g2_or3_1 _4062_ (.A(_1128_),
    .B(_1129_),
    .C(_1133_),
    .X(_1163_));
 sg13g2_nand2_1 _4063_ (.Y(_1164_),
    .A(_1134_),
    .B(_1163_));
 sg13g2_mux2_1 _4064_ (.A0(_1164_),
    .A1(_1132_),
    .S(net625),
    .X(_1165_));
 sg13g2_xnor2_1 _4065_ (.Y(_1166_),
    .A(net750),
    .B(_1165_));
 sg13g2_inv_1 _4066_ (.Y(_1167_),
    .A(_1166_));
 sg13g2_or2_1 _4067_ (.X(_1168_),
    .B(_1165_),
    .A(\core.C_q[9] ));
 sg13g2_o21ai_1 _4068_ (.B1(_1168_),
    .Y(_1169_),
    .A1(_1167_),
    .A2(_1162_));
 sg13g2_nand2_1 _4069_ (.Y(_1170_),
    .A(_1113_),
    .B(net625));
 sg13g2_nand3_1 _4070_ (.B(_1135_),
    .C(_1137_),
    .A(_1134_),
    .Y(_1171_));
 sg13g2_nand2b_1 _4071_ (.Y(_1172_),
    .B(_1171_),
    .A_N(_1138_));
 sg13g2_o21ai_1 _4072_ (.B1(_1170_),
    .Y(_1173_),
    .A1(net625),
    .A2(_1172_));
 sg13g2_xor2_1 _4073_ (.B(_1173_),
    .A(_0031_),
    .X(_1174_));
 sg13g2_a22oi_1 _4074_ (.Y(_1175_),
    .B1(_1169_),
    .B2(_1174_),
    .A2(_1173_),
    .A1(_1950_));
 sg13g2_xnor2_1 _4075_ (.Y(_1176_),
    .A(_0025_),
    .B(_1175_));
 sg13g2_inv_1 _4076_ (.Y(_1177_),
    .A(_1176_));
 sg13g2_nand2_1 _4077_ (.Y(_1178_),
    .A(_1142_),
    .B(_1177_));
 sg13g2_nand2_1 _4078_ (.Y(_1179_),
    .A(_0025_),
    .B(_1142_));
 sg13g2_a22oi_1 _4079_ (.Y(_1180_),
    .B1(_1179_),
    .B2(_1175_),
    .A2(_1107_),
    .A1(_1962_));
 sg13g2_inv_1 _4080_ (.Y(_1181_),
    .A(net624));
 sg13g2_xnor2_1 _4081_ (.Y(_1182_),
    .A(_1169_),
    .B(_1174_));
 sg13g2_nor2_1 _4082_ (.A(_1173_),
    .B(net623),
    .Y(_1183_));
 sg13g2_a21oi_2 _4083_ (.B1(_1183_),
    .Y(_1184_),
    .A2(_1182_),
    .A1(net623));
 sg13g2_nand2_1 _4084_ (.Y(_1185_),
    .A(_0025_),
    .B(_1184_));
 sg13g2_inv_1 _4085_ (.Y(_1186_),
    .A(_1185_));
 sg13g2_xnor2_1 _4086_ (.Y(_1187_),
    .A(_1962_),
    .B(_1184_));
 sg13g2_nand2_1 _4087_ (.Y(_1188_),
    .A(net758),
    .B(_1145_));
 sg13g2_a221oi_1 _4088_ (.B2(_1179_),
    .C1(_1118_),
    .B1(_1175_),
    .A1(_1962_),
    .Y(_1189_),
    .A2(_1107_));
 sg13g2_xnor2_1 _4089_ (.Y(_1190_),
    .A(_1188_),
    .B(_1189_));
 sg13g2_xnor2_1 _4090_ (.Y(_1191_),
    .A(net752),
    .B(_1190_));
 sg13g2_and2_2 _4091_ (.A(net758),
    .B(net624),
    .X(_1192_));
 sg13g2_a21oi_1 _4092_ (.A1(net755),
    .A2(net757),
    .Y(_1193_),
    .B1(net753));
 sg13g2_mux2_1 _4093_ (.A0(_1116_),
    .A1(_1193_),
    .S(_1192_),
    .X(_1194_));
 sg13g2_nand2_1 _4094_ (.Y(_1195_),
    .A(_1954_),
    .B(_1190_));
 sg13g2_o21ai_1 _4095_ (.B1(_1195_),
    .Y(_1196_),
    .A1(_1194_),
    .A2(_1191_));
 sg13g2_nor2_1 _4096_ (.A(_1147_),
    .B(net624),
    .Y(_1197_));
 sg13g2_xnor2_1 _4097_ (.Y(_1198_),
    .A(_1148_),
    .B(_1149_));
 sg13g2_a21oi_2 _4098_ (.B1(_1197_),
    .Y(_1199_),
    .A2(_1198_),
    .A1(net624));
 sg13g2_inv_1 _4099_ (.Y(_1200_),
    .A(_1199_));
 sg13g2_xnor2_1 _4100_ (.Y(_1201_),
    .A(_1966_),
    .B(_1199_));
 sg13g2_a22oi_1 _4101_ (.Y(_1202_),
    .B1(_1196_),
    .B2(_1201_),
    .A2(_1199_),
    .A1(_1953_));
 sg13g2_xnor2_1 _4102_ (.Y(_1203_),
    .A(_1150_),
    .B(_1155_));
 sg13g2_nor2_1 _4103_ (.A(_1153_),
    .B(net623),
    .Y(_1204_));
 sg13g2_a21oi_2 _4104_ (.B1(_1204_),
    .Y(_1205_),
    .A2(_1203_),
    .A1(net623));
 sg13g2_xnor2_1 _4105_ (.Y(_1206_),
    .A(net751),
    .B(_1205_));
 sg13g2_nand2_1 _4106_ (.Y(_1207_),
    .A(_1952_),
    .B(_1205_));
 sg13g2_o21ai_1 _4107_ (.B1(_1207_),
    .Y(_1208_),
    .A1(_1206_),
    .A2(_1202_));
 sg13g2_xnor2_1 _4108_ (.Y(_1209_),
    .A(_1157_),
    .B(_1161_));
 sg13g2_nand2_1 _4109_ (.Y(_1210_),
    .A(net623),
    .B(_1209_));
 sg13g2_o21ai_1 _4110_ (.B1(_1210_),
    .Y(_1211_),
    .A1(_1160_),
    .A2(net623));
 sg13g2_inv_1 _4111_ (.Y(_1212_),
    .A(_1211_));
 sg13g2_xnor2_1 _4112_ (.Y(_1213_),
    .A(net750),
    .B(_1211_));
 sg13g2_a22oi_1 _4113_ (.Y(_1214_),
    .B1(_1208_),
    .B2(_1213_),
    .A2(_1212_),
    .A1(_1951_));
 sg13g2_xnor2_1 _4114_ (.Y(_1215_),
    .A(_1162_),
    .B(_1166_));
 sg13g2_nand2_1 _4115_ (.Y(_1216_),
    .A(net623),
    .B(_1215_));
 sg13g2_o21ai_1 _4116_ (.B1(_1216_),
    .Y(_1217_),
    .A1(_1165_),
    .A2(net623));
 sg13g2_xor2_1 _4117_ (.B(_1217_),
    .A(_0031_),
    .X(_1218_));
 sg13g2_inv_1 _4118_ (.Y(_1219_),
    .A(_1218_));
 sg13g2_nand2_1 _4119_ (.Y(_1220_),
    .A(_1950_),
    .B(_1217_));
 sg13g2_o21ai_1 _4120_ (.B1(_1220_),
    .Y(_1221_),
    .A1(_1219_),
    .A2(_1214_));
 sg13g2_nand2_1 _4121_ (.Y(_1222_),
    .A(_1187_),
    .B(_1221_));
 sg13g2_a21o_1 _4122_ (.A2(_1222_),
    .A1(_1185_),
    .B1(_1178_),
    .X(_1223_));
 sg13g2_a221oi_1 _4123_ (.B2(_1187_),
    .C1(_1186_),
    .B1(_1221_),
    .A1(_1142_),
    .Y(_1224_),
    .A2(_1177_));
 sg13g2_nand3_1 _4124_ (.B(_1185_),
    .C(_1222_),
    .A(_1178_),
    .Y(_1225_));
 sg13g2_xor2_1 _4125_ (.B(_1213_),
    .A(_1208_),
    .X(_1226_));
 sg13g2_nand2_1 _4126_ (.Y(_1227_),
    .A(_1225_),
    .B(_1226_));
 sg13g2_o21ai_1 _4127_ (.B1(_1227_),
    .Y(_1228_),
    .A1(_1211_),
    .A2(_1225_));
 sg13g2_and2_1 _4128_ (.A(_1950_),
    .B(_1228_),
    .X(_1229_));
 sg13g2_nand2_1 _4129_ (.Y(_1230_),
    .A(_1205_),
    .B(net619));
 sg13g2_xnor2_1 _4130_ (.Y(_1231_),
    .A(_1202_),
    .B(_1206_));
 sg13g2_o21ai_1 _4131_ (.B1(_1230_),
    .Y(_1232_),
    .A1(net619),
    .A2(_1231_));
 sg13g2_nand2_1 _4132_ (.Y(_1233_),
    .A(_1951_),
    .B(_1232_));
 sg13g2_or3_1 _4133_ (.A(_1118_),
    .B(_1192_),
    .C(_1224_),
    .X(_1234_));
 sg13g2_o21ai_1 _4134_ (.B1(_1192_),
    .Y(_1235_),
    .A1(_1118_),
    .A2(_1224_));
 sg13g2_nand2_1 _4135_ (.Y(_1236_),
    .A(_1234_),
    .B(_1235_));
 sg13g2_a21o_1 _4136_ (.A2(_1235_),
    .A1(_1234_),
    .B1(net682),
    .X(_1237_));
 sg13g2_nand3_1 _4137_ (.B(_1234_),
    .C(_1235_),
    .A(net682),
    .Y(_1238_));
 sg13g2_nand2_1 _4138_ (.Y(_1239_),
    .A(_1237_),
    .B(_1238_));
 sg13g2_a21oi_1 _4139_ (.A1(net758),
    .A2(net619),
    .Y(_1240_),
    .B1(net755));
 sg13g2_nand3_1 _4140_ (.B(_1238_),
    .C(_1240_),
    .A(_1237_),
    .Y(_1241_));
 sg13g2_nand2_1 _4141_ (.Y(_1242_),
    .A(_1954_),
    .B(_1236_));
 sg13g2_a21oi_1 _4142_ (.A1(net753),
    .A2(_1192_),
    .Y(_1243_),
    .B1(_1089_));
 sg13g2_xnor2_1 _4143_ (.Y(_1244_),
    .A(_1191_),
    .B(_1243_));
 sg13g2_nand2_2 _4144_ (.Y(_1245_),
    .A(_1190_),
    .B(net619));
 sg13g2_o21ai_1 _4145_ (.B1(_1245_),
    .Y(_1246_),
    .A1(_1224_),
    .A2(_1244_));
 sg13g2_xnor2_1 _4146_ (.Y(_1247_),
    .A(_0022_),
    .B(_1246_));
 sg13g2_a21o_1 _4147_ (.A2(_1242_),
    .A1(_1241_),
    .B1(_1247_),
    .X(_1248_));
 sg13g2_nand2_1 _4148_ (.Y(_1249_),
    .A(_1953_),
    .B(_1246_));
 sg13g2_xnor2_1 _4149_ (.Y(_1250_),
    .A(_1196_),
    .B(_1201_));
 sg13g2_mux2_2 _4150_ (.A0(_1250_),
    .A1(_1200_),
    .S(net619),
    .X(_1251_));
 sg13g2_xnor2_1 _4151_ (.Y(_1252_),
    .A(net751),
    .B(_1251_));
 sg13g2_inv_1 _4152_ (.Y(_1253_),
    .A(_1252_));
 sg13g2_a21o_1 _4153_ (.A2(_1249_),
    .A1(_1248_),
    .B1(_1253_),
    .X(_1254_));
 sg13g2_or2_1 _4154_ (.X(_1255_),
    .B(_1251_),
    .A(\core.C_q[8] ));
 sg13g2_xor2_1 _4155_ (.B(_1232_),
    .A(net750),
    .X(_1256_));
 sg13g2_inv_1 _4156_ (.Y(_1257_),
    .A(_1256_));
 sg13g2_a21o_1 _4157_ (.A2(_1254_),
    .A1(_1255_),
    .B1(_1257_),
    .X(_1258_));
 sg13g2_xor2_1 _4158_ (.B(_1228_),
    .A(_0031_),
    .X(_1259_));
 sg13g2_inv_1 _4159_ (.Y(_1260_),
    .A(_1259_));
 sg13g2_a21oi_2 _4160_ (.B1(_1260_),
    .Y(_1261_),
    .A2(_1233_),
    .A1(_1258_));
 sg13g2_nor2_1 _4161_ (.A(_1229_),
    .B(_1261_),
    .Y(_1262_));
 sg13g2_xnor2_1 _4162_ (.Y(_1263_),
    .A(_1214_),
    .B(_1219_));
 sg13g2_nand2_1 _4163_ (.Y(_1264_),
    .A(_1217_),
    .B(net619));
 sg13g2_o21ai_1 _4164_ (.B1(_1264_),
    .Y(_1265_),
    .A1(net619),
    .A2(_1263_));
 sg13g2_xnor2_1 _4165_ (.Y(_1266_),
    .A(_1962_),
    .B(_1265_));
 sg13g2_o21ai_1 _4166_ (.B1(_1266_),
    .Y(_1267_),
    .A1(_1261_),
    .A2(_1229_));
 sg13g2_nand2_1 _4167_ (.Y(_1268_),
    .A(_1949_),
    .B(_1265_));
 sg13g2_and2_1 _4168_ (.A(_1267_),
    .B(_1268_),
    .X(_1269_));
 sg13g2_nor2_1 _4169_ (.A(_1184_),
    .B(_1225_),
    .Y(_1270_));
 sg13g2_xnor2_1 _4170_ (.Y(_1271_),
    .A(_1187_),
    .B(_1221_));
 sg13g2_a21oi_1 _4171_ (.A1(_1225_),
    .A2(_1271_),
    .Y(_1272_),
    .B1(_1270_));
 sg13g2_inv_1 _4172_ (.Y(_1273_),
    .A(_1272_));
 sg13g2_and2_1 _4173_ (.A(_1269_),
    .B(_1273_),
    .X(_1274_));
 sg13g2_nor2_2 _4174_ (.A(_1223_),
    .B(_1274_),
    .Y(_1275_));
 sg13g2_and4_1 _4175_ (.A(_1223_),
    .B(_1267_),
    .C(_1268_),
    .D(_1273_),
    .X(_1276_));
 sg13g2_nand4_1 _4176_ (.B(_1223_),
    .C(_1268_),
    .A(_1267_),
    .Y(_1277_),
    .D(_1273_));
 sg13g2_nand3_1 _4177_ (.B(_1258_),
    .C(_1260_),
    .A(_1233_),
    .Y(_1278_));
 sg13g2_nand2b_1 _4178_ (.Y(_1279_),
    .B(_1278_),
    .A_N(_1261_));
 sg13g2_nand2_1 _4179_ (.Y(_1280_),
    .A(_1228_),
    .B(net616));
 sg13g2_o21ai_1 _4180_ (.B1(_1280_),
    .Y(_1281_),
    .A1(net616),
    .A2(_1279_));
 sg13g2_nor2_1 _4181_ (.A(_0025_),
    .B(_1281_),
    .Y(_1282_));
 sg13g2_nand2b_1 _4182_ (.Y(_1283_),
    .B(_1962_),
    .A_N(_1281_));
 sg13g2_xnor2_1 _4183_ (.Y(_1284_),
    .A(_1239_),
    .B(_1240_));
 sg13g2_mux2_1 _4184_ (.A0(_1236_),
    .A1(_1284_),
    .S(_1277_),
    .X(_1285_));
 sg13g2_xnor2_1 _4185_ (.Y(_1286_),
    .A(_0022_),
    .B(_1285_));
 sg13g2_inv_2 _4186_ (.Y(_1287_),
    .A(_1286_));
 sg13g2_nand2_1 _4187_ (.Y(_1288_),
    .A(net758),
    .B(_1225_));
 sg13g2_and3_1 _4188_ (.X(_1289_),
    .A(_1117_),
    .B(_1277_),
    .C(_1288_));
 sg13g2_a21oi_2 _4189_ (.B1(_1288_),
    .Y(_1290_),
    .A2(_1277_),
    .A1(_1117_));
 sg13g2_or2_1 _4190_ (.X(_1291_),
    .B(_1290_),
    .A(_1289_));
 sg13g2_inv_1 _4191_ (.Y(_1292_),
    .A(_1291_));
 sg13g2_nor3_1 _4192_ (.A(net752),
    .B(_1289_),
    .C(_1290_),
    .Y(_1293_));
 sg13g2_o21ai_1 _4193_ (.B1(net752),
    .Y(_1294_),
    .A1(_1289_),
    .A2(_1290_));
 sg13g2_nor2_1 _4194_ (.A(_1955_),
    .B(net617),
    .Y(_1295_));
 sg13g2_a21oi_1 _4195_ (.A1(net753),
    .A2(_1295_),
    .Y(_1296_),
    .B1(_1089_));
 sg13g2_o21ai_1 _4196_ (.B1(_1294_),
    .Y(_1297_),
    .A1(_1293_),
    .A2(_1296_));
 sg13g2_and2_1 _4197_ (.A(_1953_),
    .B(_1285_),
    .X(_1298_));
 sg13g2_a21o_1 _4198_ (.A2(_1297_),
    .A1(_1287_),
    .B1(_1298_),
    .X(_1299_));
 sg13g2_nand2_1 _4199_ (.Y(_1300_),
    .A(_1246_),
    .B(net616));
 sg13g2_nand3_1 _4200_ (.B(_1242_),
    .C(_1247_),
    .A(_1241_),
    .Y(_1301_));
 sg13g2_nand2_1 _4201_ (.Y(_1302_),
    .A(_1248_),
    .B(_1301_));
 sg13g2_o21ai_1 _4202_ (.B1(_1300_),
    .Y(_1303_),
    .A1(net616),
    .A2(_1302_));
 sg13g2_xor2_1 _4203_ (.B(_1303_),
    .A(net751),
    .X(_1304_));
 sg13g2_a22oi_1 _4204_ (.Y(_1305_),
    .B1(_1304_),
    .B2(_1299_),
    .A2(_1303_),
    .A1(_1952_));
 sg13g2_nand3_1 _4205_ (.B(_1249_),
    .C(_1253_),
    .A(_1248_),
    .Y(_1306_));
 sg13g2_a21oi_1 _4206_ (.A1(_1254_),
    .A2(_1306_),
    .Y(_1307_),
    .B1(net617));
 sg13g2_a21oi_2 _4207_ (.B1(_1307_),
    .Y(_1308_),
    .A2(net617),
    .A1(_1251_));
 sg13g2_xnor2_1 _4208_ (.Y(_1309_),
    .A(net750),
    .B(_1308_));
 sg13g2_nand2_1 _4209_ (.Y(_1310_),
    .A(_1951_),
    .B(_1308_));
 sg13g2_o21ai_1 _4210_ (.B1(_1310_),
    .Y(_1311_),
    .A1(_1309_),
    .A2(_1305_));
 sg13g2_nand3_1 _4211_ (.B(_1255_),
    .C(_1257_),
    .A(_1254_),
    .Y(_1312_));
 sg13g2_nand2_1 _4212_ (.Y(_1313_),
    .A(_1258_),
    .B(_1312_));
 sg13g2_nand2_1 _4213_ (.Y(_1314_),
    .A(_1232_),
    .B(net616));
 sg13g2_o21ai_1 _4214_ (.B1(_1314_),
    .Y(_1315_),
    .A1(net616),
    .A2(_1313_));
 sg13g2_xor2_1 _4215_ (.B(_1315_),
    .A(_0031_),
    .X(_1316_));
 sg13g2_a22oi_1 _4216_ (.Y(_1317_),
    .B1(_1311_),
    .B2(_1316_),
    .A2(_1315_),
    .A1(_1950_));
 sg13g2_xor2_1 _4217_ (.B(_1266_),
    .A(_1262_),
    .X(_1318_));
 sg13g2_nor2_1 _4218_ (.A(net616),
    .B(_1318_),
    .Y(_1319_));
 sg13g2_a21oi_1 _4219_ (.A1(_1265_),
    .A2(net616),
    .Y(_1320_),
    .B1(_1319_));
 sg13g2_nand2_1 _4220_ (.Y(_1321_),
    .A(_0025_),
    .B(_1281_));
 sg13g2_and2_1 _4221_ (.A(_1320_),
    .B(_1321_),
    .X(_1322_));
 sg13g2_o21ai_1 _4222_ (.B1(_1322_),
    .Y(_1323_),
    .A1(_1317_),
    .A2(_1282_));
 sg13g2_nand2b_1 _4223_ (.Y(_1324_),
    .B(_1274_),
    .A_N(_1223_));
 sg13g2_o21ai_1 _4224_ (.B1(_1324_),
    .Y(_1325_),
    .A1(_1269_),
    .A2(_1273_));
 sg13g2_or2_1 _4225_ (.X(_1326_),
    .B(_1325_),
    .A(_1323_));
 sg13g2_nor3_1 _4226_ (.A(_1275_),
    .B(_1323_),
    .C(_1325_),
    .Y(_1327_));
 sg13g2_or3_2 _4227_ (.A(_1323_),
    .B(_1275_),
    .C(_1325_),
    .X(_1328_));
 sg13g2_xnor2_1 _4228_ (.Y(_1329_),
    .A(_1311_),
    .B(_1316_));
 sg13g2_nand2_1 _4229_ (.Y(_1330_),
    .A(_1315_),
    .B(net613));
 sg13g2_o21ai_1 _4230_ (.B1(_1330_),
    .Y(_1331_),
    .A1(net613),
    .A2(_1329_));
 sg13g2_and2_1 _4231_ (.A(_1949_),
    .B(_1331_),
    .X(_1332_));
 sg13g2_nor2_1 _4232_ (.A(_1949_),
    .B(_1331_),
    .Y(_1333_));
 sg13g2_xnor2_1 _4233_ (.Y(_1334_),
    .A(_1305_),
    .B(_1309_));
 sg13g2_nand2_1 _4234_ (.Y(_1335_),
    .A(_1328_),
    .B(_1334_));
 sg13g2_o21ai_1 _4235_ (.B1(_1335_),
    .Y(_1336_),
    .A1(_1308_),
    .A2(_1328_));
 sg13g2_xor2_1 _4236_ (.B(_1336_),
    .A(_0031_),
    .X(_1337_));
 sg13g2_or3_1 _4237_ (.A(_1332_),
    .B(_1333_),
    .C(_1337_),
    .X(_1338_));
 sg13g2_xnor2_1 _4238_ (.Y(_1339_),
    .A(_1286_),
    .B(_1297_));
 sg13g2_mux2_1 _4239_ (.A0(_1285_),
    .A1(_1339_),
    .S(_1328_),
    .X(_1340_));
 sg13g2_nor2_1 _4240_ (.A(net751),
    .B(_1340_),
    .Y(_1341_));
 sg13g2_nor2b_1 _4241_ (.A(_1293_),
    .B_N(_1294_),
    .Y(_1342_));
 sg13g2_xnor2_1 _4242_ (.Y(_1343_),
    .A(_1296_),
    .B(_1342_));
 sg13g2_nor4_1 _4243_ (.A(_1275_),
    .B(_1292_),
    .C(_1323_),
    .D(_1325_),
    .Y(_1344_));
 sg13g2_a21oi_1 _4244_ (.A1(_1328_),
    .A2(_1343_),
    .Y(_1345_),
    .B1(_1344_));
 sg13g2_nor2_1 _4245_ (.A(net339),
    .B(_1345_),
    .Y(_1346_));
 sg13g2_a21oi_1 _4246_ (.A1(net751),
    .A2(_1340_),
    .Y(_1347_),
    .B1(_1346_));
 sg13g2_nand3b_1 _4247_ (.B(_1328_),
    .C(_1117_),
    .Y(_1348_),
    .A_N(_1295_));
 sg13g2_o21ai_1 _4248_ (.B1(_1295_),
    .Y(_1349_),
    .A1(_1118_),
    .A2(_1327_));
 sg13g2_a21oi_1 _4249_ (.A1(_1348_),
    .A2(_1349_),
    .Y(_1350_),
    .B1(net682));
 sg13g2_and3_1 _4250_ (.X(_1351_),
    .A(_1348_),
    .B(net682),
    .C(_1349_));
 sg13g2_nor3_1 _4251_ (.A(net755),
    .B(_1955_),
    .C(net613),
    .Y(_1352_));
 sg13g2_a21oi_1 _4252_ (.A1(net755),
    .A2(net613),
    .Y(_1353_),
    .B1(_1955_));
 sg13g2_nor2_1 _4253_ (.A(_1964_),
    .B(_1353_),
    .Y(_1354_));
 sg13g2_or4_1 _4254_ (.A(_1350_),
    .B(_1354_),
    .C(_1352_),
    .D(_1351_),
    .X(_1355_));
 sg13g2_nand2_1 _4255_ (.Y(_1356_),
    .A(net338),
    .B(_1345_));
 sg13g2_nand3_1 _4256_ (.B(_1348_),
    .C(_1349_),
    .A(\core.C_q[6] ),
    .Y(_1357_));
 sg13g2_and2_1 _4257_ (.A(_1356_),
    .B(_1357_),
    .X(_1358_));
 sg13g2_a221oi_1 _4258_ (.B2(_1355_),
    .C1(_1346_),
    .B1(_1358_),
    .A1(net751),
    .Y(_1359_),
    .A2(_1340_));
 sg13g2_nand2_1 _4259_ (.Y(_1360_),
    .A(_1303_),
    .B(net613));
 sg13g2_xnor2_1 _4260_ (.Y(_1361_),
    .A(_1299_),
    .B(_1304_));
 sg13g2_o21ai_1 _4261_ (.B1(_1360_),
    .Y(_1362_),
    .A1(net613),
    .A2(_1361_));
 sg13g2_xor2_1 _4262_ (.B(_1362_),
    .A(net750),
    .X(_1363_));
 sg13g2_o21ai_1 _4263_ (.B1(_1363_),
    .Y(_1364_),
    .A1(_1359_),
    .A2(_1341_));
 sg13g2_or2_1 _4264_ (.X(_1365_),
    .B(_1362_),
    .A(_1951_));
 sg13g2_a21oi_2 _4265_ (.B1(_1338_),
    .Y(_1366_),
    .A2(_1364_),
    .A1(_1365_));
 sg13g2_a21oi_1 _4266_ (.A1(net342),
    .A2(_1336_),
    .Y(_1367_),
    .B1(_1333_));
 sg13g2_a21oi_1 _4267_ (.A1(_1949_),
    .A2(_1331_),
    .Y(_1368_),
    .B1(_1367_));
 sg13g2_a21oi_1 _4268_ (.A1(_1283_),
    .A2(_1321_),
    .Y(_1369_),
    .B1(_1317_));
 sg13g2_o21ai_1 _4269_ (.B1(_1323_),
    .Y(_1370_),
    .A1(_1282_),
    .A2(_1320_));
 sg13g2_nand3b_1 _4270_ (.B(_1320_),
    .C(net613),
    .Y(_1371_),
    .A_N(_1281_));
 sg13g2_o21ai_1 _4271_ (.B1(_1371_),
    .Y(_1372_),
    .A1(_1369_),
    .A2(_1370_));
 sg13g2_a21oi_1 _4272_ (.A1(_1323_),
    .A2(_1325_),
    .Y(_1373_),
    .B1(_1275_));
 sg13g2_nand2_1 _4273_ (.Y(_1374_),
    .A(_1372_),
    .B(_1373_));
 sg13g2_nor2b_1 _4274_ (.A(_1341_),
    .B_N(_1089_),
    .Y(_1375_));
 sg13g2_nand4_1 _4275_ (.B(_1356_),
    .C(_1363_),
    .A(_1347_),
    .Y(_1376_),
    .D(_1375_));
 sg13g2_nor4_1 _4276_ (.A(_1338_),
    .B(_1350_),
    .C(_1351_),
    .D(_1376_),
    .Y(_1377_));
 sg13g2_nor2_1 _4277_ (.A(_1374_),
    .B(_1377_),
    .Y(_1378_));
 sg13g2_o21ai_1 _4278_ (.B1(_1378_),
    .Y(_1379_),
    .A1(_1368_),
    .A2(_1366_));
 sg13g2_nand2_1 _4279_ (.Y(_1380_),
    .A(_1003_),
    .B(_1089_));
 sg13g2_a21oi_2 _4280_ (.B1(net765),
    .Y(_1381_),
    .A2(_1089_),
    .A1(_1003_));
 sg13g2_nand2_1 _4281_ (.Y(_1382_),
    .A(net681),
    .B(_1380_));
 sg13g2_a22oi_1 _4282_ (.Y(_1383_),
    .B1(_1379_),
    .B2(_1381_),
    .A2(net764),
    .A1(net569));
 sg13g2_inv_1 _4283_ (.Y(_0079_),
    .A(_1383_));
 sg13g2_nand2_1 _4284_ (.Y(_1384_),
    .A(net762),
    .B(_1379_));
 sg13g2_xnor2_1 _4285_ (.Y(_1385_),
    .A(net613),
    .B(_1384_));
 sg13g2_nand2_1 _4286_ (.Y(_1386_),
    .A(net475),
    .B(net765));
 sg13g2_o21ai_1 _4287_ (.B1(_1386_),
    .Y(_0080_),
    .A1(net643),
    .A2(_1385_));
 sg13g2_nand2_1 _4288_ (.Y(_1387_),
    .A(net447),
    .B(net765));
 sg13g2_o21ai_1 _4289_ (.B1(net762),
    .Y(_1388_),
    .A1(_1326_),
    .A2(_1379_));
 sg13g2_xnor2_1 _4290_ (.Y(_1389_),
    .A(net617),
    .B(_1388_));
 sg13g2_o21ai_1 _4291_ (.B1(_1387_),
    .Y(_0081_),
    .A1(net643),
    .A2(_1389_));
 sg13g2_nor3_1 _4292_ (.A(_1277_),
    .B(_1326_),
    .C(_1379_),
    .Y(_1390_));
 sg13g2_nand2b_1 _4293_ (.Y(_1391_),
    .B(net762),
    .A_N(_1390_));
 sg13g2_xnor2_1 _4294_ (.Y(_1392_),
    .A(net619),
    .B(_1391_));
 sg13g2_nand2_1 _4295_ (.Y(_1393_),
    .A(net455),
    .B(net764));
 sg13g2_o21ai_1 _4296_ (.B1(_1393_),
    .Y(_0082_),
    .A1(net643),
    .A2(_1392_));
 sg13g2_nor4_2 _4297_ (.A(_1225_),
    .B(_1277_),
    .C(_1379_),
    .Y(_1394_),
    .D(_1326_));
 sg13g2_nor2b_1 _4298_ (.A(_1394_),
    .B_N(net762),
    .Y(_1395_));
 sg13g2_xnor2_1 _4299_ (.Y(_1396_),
    .A(net624),
    .B(_1395_));
 sg13g2_nand2_1 _4300_ (.Y(_1397_),
    .A(net444),
    .B(net764));
 sg13g2_o21ai_1 _4301_ (.B1(_1397_),
    .Y(_0083_),
    .A1(net643),
    .A2(_1396_));
 sg13g2_nand2_1 _4302_ (.Y(_1398_),
    .A(_1181_),
    .B(_1394_));
 sg13g2_nand2_1 _4303_ (.Y(_1399_),
    .A(net761),
    .B(_1398_));
 sg13g2_xnor2_1 _4304_ (.Y(_1400_),
    .A(net625),
    .B(_1399_));
 sg13g2_nand2_1 _4305_ (.Y(_1401_),
    .A(net511),
    .B(net766));
 sg13g2_o21ai_1 _4306_ (.B1(_1401_),
    .Y(_0084_),
    .A1(net644),
    .A2(_1400_));
 sg13g2_o21ai_1 _4307_ (.B1(net761),
    .Y(_1402_),
    .A1(_1145_),
    .A2(_1398_));
 sg13g2_xnor2_1 _4308_ (.Y(_1403_),
    .A(_1110_),
    .B(_1402_));
 sg13g2_nand2_1 _4309_ (.Y(_1404_),
    .A(net464),
    .B(net765));
 sg13g2_o21ai_1 _4310_ (.B1(_1404_),
    .Y(_0085_),
    .A1(net644),
    .A2(_1403_));
 sg13g2_nand4_1 _4311_ (.B(net625),
    .C(_1181_),
    .A(_1394_),
    .Y(_1405_),
    .D(_1110_));
 sg13g2_nand2_1 _4312_ (.Y(_1406_),
    .A(net761),
    .B(_1405_));
 sg13g2_xnor2_1 _4313_ (.Y(_1407_),
    .A(_1078_),
    .B(_1406_));
 sg13g2_nand2_1 _4314_ (.Y(_1408_),
    .A(net454),
    .B(net765));
 sg13g2_o21ai_1 _4315_ (.B1(_1408_),
    .Y(_0086_),
    .A1(net643),
    .A2(_1407_));
 sg13g2_o21ai_1 _4316_ (.B1(net761),
    .Y(_1409_),
    .A1(_1079_),
    .A2(_1405_));
 sg13g2_xnor2_1 _4317_ (.Y(_1410_),
    .A(_1050_),
    .B(_1409_));
 sg13g2_nand2_1 _4318_ (.Y(_1411_),
    .A(net536),
    .B(net764));
 sg13g2_o21ai_1 _4319_ (.B1(_1411_),
    .Y(_0087_),
    .A1(net643),
    .A2(_1410_));
 sg13g2_nor3_1 _4320_ (.A(_1051_),
    .B(_1079_),
    .C(_1405_),
    .Y(_1412_));
 sg13g2_nor2b_1 _4321_ (.A(_1412_),
    .B_N(net761),
    .Y(_1413_));
 sg13g2_xnor2_1 _4322_ (.Y(_1414_),
    .A(_1034_),
    .B(_1413_));
 sg13g2_nand2_1 _4323_ (.Y(_1415_),
    .A(net503),
    .B(net765));
 sg13g2_o21ai_1 _4324_ (.B1(_1415_),
    .Y(_0088_),
    .A1(net643),
    .A2(_1414_));
 sg13g2_nor4_2 _4325_ (.A(_1034_),
    .B(_1051_),
    .C(_1405_),
    .Y(_1416_),
    .D(_1079_));
 sg13g2_nand2b_1 _4326_ (.Y(_1417_),
    .B(net761),
    .A_N(_1416_));
 sg13g2_xnor2_1 _4327_ (.Y(_1418_),
    .A(_1014_),
    .B(_1417_));
 sg13g2_nand2_1 _4328_ (.Y(_1419_),
    .A(net504),
    .B(net765));
 sg13g2_o21ai_1 _4329_ (.B1(_1419_),
    .Y(_0089_),
    .A1(net644),
    .A2(_1418_));
 sg13g2_nor2_1 _4330_ (.A(net757),
    .B(_0996_),
    .Y(_1420_));
 sg13g2_nor2_1 _4331_ (.A(_0999_),
    .B(_1420_),
    .Y(_1421_));
 sg13g2_inv_1 _4332_ (.Y(_1422_),
    .A(_1421_));
 sg13g2_nand2_2 _4333_ (.Y(_1423_),
    .A(_1416_),
    .B(_1014_));
 sg13g2_nand2_2 _4334_ (.Y(_1424_),
    .A(_1423_),
    .B(net760));
 sg13g2_xnor2_1 _4335_ (.Y(_1425_),
    .A(_1422_),
    .B(_1424_));
 sg13g2_nand2_1 _4336_ (.Y(_1426_),
    .A(net552),
    .B(net766));
 sg13g2_o21ai_1 _4337_ (.B1(_1426_),
    .Y(_0090_),
    .A1(net644),
    .A2(_1425_));
 sg13g2_and2_1 _4338_ (.A(net760),
    .B(_1381_),
    .X(_1427_));
 sg13g2_o21ai_1 _4339_ (.B1(_1427_),
    .Y(_1428_),
    .A1(_1421_),
    .A2(_1423_));
 sg13g2_o21ai_1 _4340_ (.B1(_1428_),
    .Y(_0091_),
    .A1(_1974_),
    .A2(net681));
 sg13g2_nand2_1 _4341_ (.Y(_1429_),
    .A(net561),
    .B(net766));
 sg13g2_nor2_1 _4342_ (.A(net758),
    .B(_0999_),
    .Y(_1430_));
 sg13g2_nor4_1 _4343_ (.A(net340),
    .B(net344),
    .C(_0996_),
    .D(_1021_),
    .Y(_1431_));
 sg13g2_nor2b_1 _4344_ (.A(_1380_),
    .B_N(_1431_),
    .Y(_1432_));
 sg13g2_a21oi_1 _4345_ (.A1(_1006_),
    .A2(_1432_),
    .Y(_1433_),
    .B1(_1430_));
 sg13g2_nand4_1 _4346_ (.B(_1380_),
    .C(_1014_),
    .A(_1416_),
    .Y(_1434_),
    .D(_1422_));
 sg13g2_nand2_1 _4347_ (.Y(_1435_),
    .A(_1434_),
    .B(net760));
 sg13g2_xnor2_1 _4348_ (.Y(_1436_),
    .A(_1433_),
    .B(_1435_));
 sg13g2_o21ai_1 _4349_ (.B1(_1429_),
    .Y(_0092_),
    .A1(_1436_),
    .A2(net644));
 sg13g2_o21ai_1 _4350_ (.B1(_1427_),
    .Y(_1437_),
    .A1(_1430_),
    .A2(_1434_));
 sg13g2_o21ai_1 _4351_ (.B1(_1437_),
    .Y(_0093_),
    .A1(_1975_),
    .A2(net681));
 sg13g2_a21oi_2 _4352_ (.B1(_1430_),
    .Y(_1438_),
    .A2(net760),
    .A1(_1434_));
 sg13g2_a21o_1 _4353_ (.A2(_1430_),
    .A1(net760),
    .B1(net643),
    .X(_1439_));
 sg13g2_nand2_1 _4354_ (.Y(_1440_),
    .A(net551),
    .B(net766));
 sg13g2_o21ai_1 _4355_ (.B1(_1440_),
    .Y(_0094_),
    .A1(_1439_),
    .A2(_1438_));
 sg13g2_mux2_1 _4356_ (.A0(net728),
    .A1(net818),
    .S(net767),
    .X(_0095_));
 sg13g2_xnor2_1 _4357_ (.Y(_1441_),
    .A(net319),
    .B(net728));
 sg13g2_nand2_1 _4358_ (.Y(_1442_),
    .A(net499),
    .B(net767));
 sg13g2_o21ai_1 _4359_ (.B1(_1442_),
    .Y(_0096_),
    .A1(net767),
    .A2(_1441_));
 sg13g2_nor2b_1 _4360_ (.A(net727),
    .B_N(net725),
    .Y(_1443_));
 sg13g2_xnor2_1 _4361_ (.Y(_1444_),
    .A(net721),
    .B(_1443_));
 sg13g2_nand2_1 _4362_ (.Y(_1445_),
    .A(net431),
    .B(net767));
 sg13g2_o21ai_1 _4363_ (.B1(_1445_),
    .Y(_0097_),
    .A1(net767),
    .A2(_1444_));
 sg13g2_o21ai_1 _4364_ (.B1(net790),
    .Y(_1446_),
    .A1(net693),
    .A2(net758));
 sg13g2_a21oi_1 _4365_ (.A1(net693),
    .A2(_1890_),
    .Y(_0098_),
    .B1(_1446_));
 sg13g2_o21ai_1 _4366_ (.B1(net790),
    .Y(_1447_),
    .A1(net688),
    .A2(net756));
 sg13g2_a21oi_1 _4367_ (.A1(net688),
    .A2(_1888_),
    .Y(_0099_),
    .B1(_1447_));
 sg13g2_o21ai_1 _4368_ (.B1(net790),
    .Y(_1448_),
    .A1(net688),
    .A2(\core.C_q[6] ));
 sg13g2_a21oi_1 _4369_ (.A1(net689),
    .A2(_1886_),
    .Y(_0100_),
    .B1(_1448_));
 sg13g2_a21oi_1 _4370_ (.A1(net692),
    .A2(net576),
    .Y(_1449_),
    .B1(net773));
 sg13g2_o21ai_1 _4371_ (.B1(_1449_),
    .Y(_0101_),
    .A1(net688),
    .A2(net824));
 sg13g2_o21ai_1 _4372_ (.B1(net790),
    .Y(_1450_),
    .A1(net688),
    .A2(\core.C_q[8] ));
 sg13g2_a21oi_1 _4373_ (.A1(net688),
    .A2(_1884_),
    .Y(_0102_),
    .B1(_1450_));
 sg13g2_o21ai_1 _4374_ (.B1(net790),
    .Y(_1451_),
    .A1(net688),
    .A2(\core.C_q[9] ));
 sg13g2_a21oi_1 _4375_ (.A1(net688),
    .A2(_1882_),
    .Y(_0103_),
    .B1(_1451_));
 sg13g2_a21oi_2 _4376_ (.B1(net774),
    .Y(_1452_),
    .A2(net855),
    .A1(net692));
 sg13g2_o21ai_1 _4377_ (.B1(_1452_),
    .Y(_0104_),
    .A1(net689),
    .A2(_1950_));
 sg13g2_a21oi_1 _4378_ (.A1(net692),
    .A2(\core.p_C[7] ),
    .Y(_1453_),
    .B1(net773));
 sg13g2_o21ai_1 _4379_ (.B1(_1453_),
    .Y(_0105_),
    .A1(net689),
    .A2(_1949_));
 sg13g2_o21ai_1 _4380_ (.B1(net790),
    .Y(_1454_),
    .A1(net690),
    .A2(\core.VT_q[4] ));
 sg13g2_a21oi_1 _4381_ (.A1(net691),
    .A2(_1898_),
    .Y(_0106_),
    .B1(_1454_));
 sg13g2_a21oi_1 _4382_ (.A1(net692),
    .A2(\core.p_VT[1] ),
    .Y(_1455_),
    .B1(net773));
 sg13g2_o21ai_1 _4383_ (.B1(_1455_),
    .Y(_0107_),
    .A1(net691),
    .A2(_1947_));
 sg13g2_a21oi_1 _4384_ (.A1(net690),
    .A2(\core.p_VT[2] ),
    .Y(_1456_),
    .B1(net773));
 sg13g2_o21ai_1 _4385_ (.B1(_1456_),
    .Y(_0108_),
    .A1(net690),
    .A2(_1946_));
 sg13g2_a21oi_1 _4386_ (.A1(net690),
    .A2(\core.p_VT[3] ),
    .Y(_1457_),
    .B1(net773));
 sg13g2_o21ai_1 _4387_ (.B1(_1457_),
    .Y(_0109_),
    .A1(net690),
    .A2(_1945_));
 sg13g2_o21ai_1 _4388_ (.B1(net788),
    .Y(_1458_),
    .A1(net690),
    .A2(\core.VT_q[8] ));
 sg13g2_a21oi_1 _4389_ (.A1(net691),
    .A2(_1894_),
    .Y(_0110_),
    .B1(_1458_));
 sg13g2_o21ai_1 _4390_ (.B1(net788),
    .Y(_1459_),
    .A1(net690),
    .A2(\core.VT_q[9] ));
 sg13g2_a21oi_1 _4391_ (.A1(net691),
    .A2(_1892_),
    .Y(_0111_),
    .B1(_1459_));
 sg13g2_a21oi_1 _4392_ (.A1(net706),
    .A2(\core.p_VT[6] ),
    .Y(_1460_),
    .B1(net774));
 sg13g2_o21ai_1 _4393_ (.B1(_1460_),
    .Y(_0112_),
    .A1(net699),
    .A2(_1943_));
 sg13g2_a21oi_1 _4394_ (.A1(net692),
    .A2(net467),
    .Y(_1461_),
    .B1(net773));
 sg13g2_o21ai_1 _4395_ (.B1(_1461_),
    .Y(_0113_),
    .A1(net690),
    .A2(_1942_));
 sg13g2_a21oi_1 _4396_ (.A1(net699),
    .A2(\core.p_Vreset[0] ),
    .Y(_1462_),
    .B1(net774));
 sg13g2_o21ai_1 _4397_ (.B1(_1462_),
    .Y(_0114_),
    .A1(net697),
    .A2(_1941_));
 sg13g2_a21oi_1 _4398_ (.A1(net697),
    .A2(\core.p_Vreset[1] ),
    .Y(_1463_),
    .B1(net774));
 sg13g2_o21ai_1 _4399_ (.B1(_1463_),
    .Y(_0115_),
    .A1(net697),
    .A2(_1940_));
 sg13g2_a21oi_1 _4400_ (.A1(net699),
    .A2(net527),
    .Y(_1464_),
    .B1(net776));
 sg13g2_o21ai_1 _4401_ (.B1(_1464_),
    .Y(_0116_),
    .A1(net699),
    .A2(_1939_));
 sg13g2_a21oi_1 _4402_ (.A1(net699),
    .A2(\core.p_Vreset[3] ),
    .Y(_1465_),
    .B1(net776));
 sg13g2_o21ai_1 _4403_ (.B1(_1465_),
    .Y(_0117_),
    .A1(net697),
    .A2(_1938_));
 sg13g2_a21oi_1 _4404_ (.A1(net700),
    .A2(net473),
    .Y(_1466_),
    .B1(net774));
 sg13g2_o21ai_1 _4405_ (.B1(_1466_),
    .Y(_0118_),
    .A1(net699),
    .A2(_1937_));
 sg13g2_a21oi_1 _4406_ (.A1(net699),
    .A2(\core.p_Vreset[5] ),
    .Y(_1467_),
    .B1(net774));
 sg13g2_o21ai_1 _4407_ (.B1(_1467_),
    .Y(_0119_),
    .A1(net699),
    .A2(_1936_));
 sg13g2_o21ai_1 _4408_ (.B1(net805),
    .Y(_1468_),
    .A1(net700),
    .A2(\core.Vreset_q[10] ));
 sg13g2_a21oi_1 _4409_ (.A1(net700),
    .A2(_1900_),
    .Y(_0120_),
    .B1(_1468_));
 sg13g2_a21oi_1 _4410_ (.A1(net697),
    .A2(net413),
    .Y(_1469_),
    .B1(net774));
 sg13g2_o21ai_1 _4411_ (.B1(_1469_),
    .Y(_0121_),
    .A1(net697),
    .A2(_1935_));
 sg13g2_o21ai_1 _4412_ (.B1(net810),
    .Y(_1470_),
    .A1(net703),
    .A2(\core.b_q[4] ));
 sg13g2_a21oi_1 _4413_ (.A1(net703),
    .A2(_1906_),
    .Y(_0122_),
    .B1(_1470_));
 sg13g2_o21ai_1 _4414_ (.B1(net810),
    .Y(_1471_),
    .A1(net704),
    .A2(\core.b_q[5] ));
 sg13g2_a21oi_1 _4415_ (.A1(net704),
    .A2(_1905_),
    .Y(_0123_),
    .B1(_1471_));
 sg13g2_o21ai_1 _4416_ (.B1(net810),
    .Y(_1472_),
    .A1(net704),
    .A2(\core.b_q[6] ));
 sg13g2_a21oi_1 _4417_ (.A1(net704),
    .A2(_1904_),
    .Y(_0124_),
    .B1(_1472_));
 sg13g2_a21oi_1 _4418_ (.A1(net703),
    .A2(\core.p_b[3] ),
    .Y(_1473_),
    .B1(net775));
 sg13g2_o21ai_1 _4419_ (.B1(_1473_),
    .Y(_0125_),
    .A1(net704),
    .A2(_1934_));
 sg13g2_o21ai_1 _4420_ (.B1(net808),
    .Y(_1474_),
    .A1(net703),
    .A2(\core.b_q[8] ));
 sg13g2_a21oi_1 _4421_ (.A1(net703),
    .A2(_1903_),
    .Y(_0126_),
    .B1(_1474_));
 sg13g2_a21oi_1 _4422_ (.A1(net705),
    .A2(\core.p_b[5] ),
    .Y(_1475_),
    .B1(net775));
 sg13g2_o21ai_1 _4423_ (.B1(_1475_),
    .Y(_0127_),
    .A1(net703),
    .A2(_1933_));
 sg13g2_o21ai_1 _4424_ (.B1(net809),
    .Y(_1476_),
    .A1(net703),
    .A2(\core.b_q[10] ));
 sg13g2_a21oi_1 _4425_ (.A1(net703),
    .A2(_1902_),
    .Y(_0128_),
    .B1(_1476_));
 sg13g2_o21ai_1 _4426_ (.B1(net809),
    .Y(_1477_),
    .A1(net705),
    .A2(\core.b_q[11] ));
 sg13g2_a21oi_1 _4427_ (.A1(net705),
    .A2(_1901_),
    .Y(_0129_),
    .B1(_1477_));
 sg13g2_o21ai_1 _4428_ (.B1(net791),
    .Y(_1478_),
    .A1(net694),
    .A2(net749));
 sg13g2_a21oi_1 _4429_ (.A1(net694),
    .A2(_1913_),
    .Y(_0130_),
    .B1(_1478_));
 sg13g2_a21oi_1 _4430_ (.A1(net696),
    .A2(net843),
    .Y(_1479_),
    .B1(net773));
 sg13g2_o21ai_1 _4431_ (.B1(_1479_),
    .Y(_0131_),
    .A1(net694),
    .A2(_1932_));
 sg13g2_o21ai_1 _4432_ (.B1(net791),
    .Y(_1480_),
    .A1(net694),
    .A2(net744));
 sg13g2_a21oi_1 _4433_ (.A1(net695),
    .A2(_1912_),
    .Y(_0132_),
    .B1(_1480_));
 sg13g2_o21ai_1 _4434_ (.B1(net792),
    .Y(_1481_),
    .A1(net696),
    .A2(\core.a_q[7] ));
 sg13g2_a21oi_1 _4435_ (.A1(net696),
    .A2(_1911_),
    .Y(_0133_),
    .B1(_1481_));
 sg13g2_o21ai_1 _4436_ (.B1(net791),
    .Y(_1482_),
    .A1(net694),
    .A2(net740));
 sg13g2_a21oi_1 _4437_ (.A1(net695),
    .A2(_1910_),
    .Y(_0134_),
    .B1(_1482_));
 sg13g2_o21ai_1 _4438_ (.B1(net791),
    .Y(_1483_),
    .A1(net694),
    .A2(net739));
 sg13g2_a21oi_1 _4439_ (.A1(net694),
    .A2(_1909_),
    .Y(_0135_),
    .B1(_1483_));
 sg13g2_o21ai_1 _4440_ (.B1(net791),
    .Y(_1484_),
    .A1(net694),
    .A2(net588));
 sg13g2_a21oi_1 _4441_ (.A1(net695),
    .A2(_1908_),
    .Y(_0136_),
    .B1(_1484_));
 sg13g2_o21ai_1 _4442_ (.B1(net793),
    .Y(_1485_),
    .A1(net697),
    .A2(net309));
 sg13g2_a21oi_1 _4443_ (.A1(net697),
    .A2(_1907_),
    .Y(_0137_),
    .B1(_1485_));
 sg13g2_o21ai_1 _4444_ (.B1(net805),
    .Y(_1486_),
    .A1(net702),
    .A2(net737));
 sg13g2_a21oi_1 _4445_ (.A1(net702),
    .A2(_1918_),
    .Y(_0138_),
    .B1(_1486_));
 sg13g2_o21ai_1 _4446_ (.B1(net793),
    .Y(_1487_),
    .A1(net698),
    .A2(\core.TauW_q[5] ));
 sg13g2_a21oi_1 _4447_ (.A1(net698),
    .A2(_1917_),
    .Y(_0139_),
    .B1(_1487_));
 sg13g2_a21oi_1 _4448_ (.A1(net701),
    .A2(net839),
    .Y(_1488_),
    .B1(net776));
 sg13g2_o21ai_1 _4449_ (.B1(_1488_),
    .Y(_0140_),
    .A1(net702),
    .A2(net685));
 sg13g2_o21ai_1 _4450_ (.B1(net805),
    .Y(_1489_),
    .A1(net702),
    .A2(\core.TauW_q[7] ));
 sg13g2_a21oi_1 _4451_ (.A1(net702),
    .A2(_1916_),
    .Y(_0141_),
    .B1(_1489_));
 sg13g2_o21ai_1 _4452_ (.B1(net806),
    .Y(_1490_),
    .A1(net701),
    .A2(net729));
 sg13g2_a21oi_1 _4453_ (.A1(net701),
    .A2(_1915_),
    .Y(_0142_),
    .B1(_1490_));
 sg13g2_a21oi_1 _4454_ (.A1(net701),
    .A2(net813),
    .Y(_1491_),
    .B1(net776));
 sg13g2_o21ai_1 _4455_ (.B1(_1491_),
    .Y(_0143_),
    .A1(net701),
    .A2(_1927_));
 sg13g2_a21oi_1 _4456_ (.A1(net701),
    .A2(net835),
    .Y(_1492_),
    .B1(net775));
 sg13g2_o21ai_1 _4457_ (.B1(_1492_),
    .Y(_0144_),
    .A1(net701),
    .A2(_1926_));
 sg13g2_o21ai_1 _4458_ (.B1(net811),
    .Y(_1493_),
    .A1(net701),
    .A2(\core.TauW_q[11] ));
 sg13g2_a21oi_1 _4459_ (.A1(net702),
    .A2(_1914_),
    .Y(_0145_),
    .B1(_1493_));
 sg13g2_o21ai_1 _4460_ (.B1(net807),
    .Y(_1494_),
    .A1(net783),
    .A2(net510));
 sg13g2_a21oi_1 _4461_ (.A1(net783),
    .A2(net636),
    .Y(_0146_),
    .B1(_1494_));
 sg13g2_nor3_1 _4462_ (.A(\core.V[14] ),
    .B(\core.V[13] ),
    .C(net868),
    .Y(_1495_));
 sg13g2_nand2b_2 _4463_ (.Y(_1496_),
    .B(net783),
    .A_N(_1495_));
 sg13g2_nor2_2 _4464_ (.A(net629),
    .B(_1496_),
    .Y(_1497_));
 sg13g2_nand2_1 _4465_ (.Y(_1498_),
    .A(net726),
    .B(net569));
 sg13g2_xor2_1 _4466_ (.B(net569),
    .A(net726),
    .X(_1499_));
 sg13g2_a22oi_1 _4467_ (.Y(_1500_),
    .B1(_1497_),
    .B2(_1499_),
    .A2(net726),
    .A1(net780));
 sg13g2_nor2_1 _4468_ (.A(net771),
    .B(_1500_),
    .Y(_0147_));
 sg13g2_nand2_1 _4469_ (.Y(_1501_),
    .A(net724),
    .B(\core.dV[1] ));
 sg13g2_xor2_1 _4470_ (.B(net475),
    .A(net724),
    .X(_1502_));
 sg13g2_nand2b_1 _4471_ (.Y(_1503_),
    .B(_1502_),
    .A_N(_1498_));
 sg13g2_xnor2_1 _4472_ (.Y(_1504_),
    .A(_1498_),
    .B(_1502_));
 sg13g2_a22oi_1 _4473_ (.Y(_1505_),
    .B1(_1497_),
    .B2(_1504_),
    .A2(net874),
    .A1(net780));
 sg13g2_nor2_1 _4474_ (.A(net771),
    .B(_1505_),
    .Y(_0148_));
 sg13g2_nand2_1 _4475_ (.Y(_1506_),
    .A(_1501_),
    .B(_1503_));
 sg13g2_xnor2_1 _4476_ (.Y(_1507_),
    .A(net722),
    .B(net447));
 sg13g2_a21oi_1 _4477_ (.A1(_1501_),
    .A2(_1503_),
    .Y(_1508_),
    .B1(_1507_));
 sg13g2_xnor2_1 _4478_ (.Y(_1509_),
    .A(_1506_),
    .B(_1507_));
 sg13g2_a22oi_1 _4479_ (.Y(_1510_),
    .B1(_1497_),
    .B2(_1509_),
    .A2(net856),
    .A1(net780));
 sg13g2_nor2_1 _4480_ (.A(net771),
    .B(net857),
    .Y(_0149_));
 sg13g2_a21o_1 _4481_ (.A2(net884),
    .A1(net722),
    .B1(_1508_),
    .X(_1511_));
 sg13g2_xnor2_1 _4482_ (.Y(_1512_),
    .A(net326),
    .B(net455));
 sg13g2_nor2b_1 _4483_ (.A(_1512_),
    .B_N(_1511_),
    .Y(_1513_));
 sg13g2_xnor2_1 _4484_ (.Y(_1514_),
    .A(_1511_),
    .B(_1512_));
 sg13g2_a22oi_1 _4485_ (.Y(_1515_),
    .B1(_1497_),
    .B2(_1514_),
    .A2(net326),
    .A1(net780));
 sg13g2_nor2_1 _4486_ (.A(net771),
    .B(_1515_),
    .Y(_0150_));
 sg13g2_a21o_1 _4487_ (.A2(\core.dV[3] ),
    .A1(net327),
    .B1(_1513_),
    .X(_1516_));
 sg13g2_and2_1 _4488_ (.A(net329),
    .B(\core.dV[4] ),
    .X(_1517_));
 sg13g2_xor2_1 _4489_ (.B(\core.dV[4] ),
    .A(net329),
    .X(_1518_));
 sg13g2_xor2_1 _4490_ (.B(_1518_),
    .A(_1516_),
    .X(_1519_));
 sg13g2_nor2_1 _4491_ (.A(net629),
    .B(_1519_),
    .Y(_1520_));
 sg13g2_nor4_1 _4492_ (.A(\core.V[11] ),
    .B(\core.V[10] ),
    .C(\core.V[9] ),
    .D(net709),
    .Y(_1521_));
 sg13g2_or4_1 _4493_ (.A(net308),
    .B(net712),
    .C(net314),
    .D(net313),
    .X(_1522_));
 sg13g2_nand3_1 _4494_ (.B(_2011_),
    .C(_1521_),
    .A(_1997_),
    .Y(_1523_));
 sg13g2_o21ai_1 _4495_ (.B1(\core.V[14] ),
    .Y(_1524_),
    .A1(_1522_),
    .A2(_1523_));
 sg13g2_nor2_2 _4496_ (.A(\core.V[15] ),
    .B(_1524_),
    .Y(_1525_));
 sg13g2_nor2_2 _4497_ (.A(_1496_),
    .B(_1525_),
    .Y(_1526_));
 sg13g2_o21ai_1 _4498_ (.B1(_1526_),
    .Y(_1527_),
    .A1(net492),
    .A2(net633));
 sg13g2_a21oi_1 _4499_ (.A1(net778),
    .A2(net848),
    .Y(_1528_),
    .B1(net772));
 sg13g2_o21ai_1 _4500_ (.B1(_1528_),
    .Y(_0151_),
    .A1(_1520_),
    .A2(_1527_));
 sg13g2_a21o_1 _4501_ (.A2(_1518_),
    .A1(_1516_),
    .B1(_1517_),
    .X(_1529_));
 sg13g2_nor2_1 _4502_ (.A(net331),
    .B(\core.dV[5] ),
    .Y(_1530_));
 sg13g2_xor2_1 _4503_ (.B(\core.dV[5] ),
    .A(net713),
    .X(_1531_));
 sg13g2_xnor2_1 _4504_ (.Y(_1532_),
    .A(_1529_),
    .B(_1531_));
 sg13g2_o21ai_1 _4505_ (.B1(_1526_),
    .Y(_1533_),
    .A1(net490),
    .A2(net633));
 sg13g2_a21oi_1 _4506_ (.A1(net632),
    .A2(_1532_),
    .Y(_1534_),
    .B1(_1533_));
 sg13g2_a21oi_1 _4507_ (.A1(net778),
    .A2(net879),
    .Y(_1535_),
    .B1(_1534_));
 sg13g2_nand2_1 _4508_ (.Y(_0152_),
    .A(net793),
    .B(_1535_));
 sg13g2_and2_1 _4509_ (.A(net711),
    .B(\core.dV[6] ),
    .X(_1536_));
 sg13g2_xnor2_1 _4510_ (.Y(_1537_),
    .A(net711),
    .B(\core.dV[6] ));
 sg13g2_a21oi_1 _4511_ (.A1(net331),
    .A2(\core.dV[5] ),
    .Y(_1538_),
    .B1(_1529_));
 sg13g2_nor3_2 _4512_ (.A(_1530_),
    .B(_1537_),
    .C(_1538_),
    .Y(_1539_));
 sg13g2_o21ai_1 _4513_ (.B1(_1537_),
    .Y(_1540_),
    .A1(_1530_),
    .A2(_1538_));
 sg13g2_nor2b_2 _4514_ (.A(_1539_),
    .B_N(_1540_),
    .Y(_1541_));
 sg13g2_nor2_1 _4515_ (.A(net840),
    .B(net633),
    .Y(_1542_));
 sg13g2_o21ai_1 _4516_ (.B1(_1526_),
    .Y(_1543_),
    .A1(net629),
    .A2(_1541_));
 sg13g2_a21oi_1 _4517_ (.A1(net779),
    .A2(net712),
    .Y(_1544_),
    .B1(net772));
 sg13g2_o21ai_1 _4518_ (.B1(_1544_),
    .Y(_0153_),
    .A1(_1542_),
    .A2(_1543_));
 sg13g2_nand2_1 _4519_ (.Y(_1545_),
    .A(net710),
    .B(\core.dV[7] ));
 sg13g2_xor2_1 _4520_ (.B(\core.dV[7] ),
    .A(net710),
    .X(_1546_));
 sg13g2_o21ai_1 _4521_ (.B1(_1546_),
    .Y(_1547_),
    .A1(_1536_),
    .A2(_1539_));
 sg13g2_or3_1 _4522_ (.A(_1536_),
    .B(_1539_),
    .C(_1546_),
    .X(_1548_));
 sg13g2_and2_1 _4523_ (.A(_1547_),
    .B(_1548_),
    .X(_1549_));
 sg13g2_nor2_1 _4524_ (.A(net533),
    .B(net633),
    .Y(_1550_));
 sg13g2_o21ai_1 _4525_ (.B1(_1526_),
    .Y(_1551_),
    .A1(net629),
    .A2(_1549_));
 sg13g2_a21oi_1 _4526_ (.A1(net779),
    .A2(net845),
    .Y(_1552_),
    .B1(net772));
 sg13g2_o21ai_1 _4527_ (.B1(_1552_),
    .Y(_0154_),
    .A1(_1550_),
    .A2(_1551_));
 sg13g2_nand2_1 _4528_ (.Y(_1553_),
    .A(net709),
    .B(\core.dV[8] ));
 sg13g2_xnor2_1 _4529_ (.Y(_1554_),
    .A(net709),
    .B(\core.dV[8] ));
 sg13g2_a21o_1 _4530_ (.A2(_1547_),
    .A1(_1545_),
    .B1(_1554_),
    .X(_1555_));
 sg13g2_nand3_1 _4531_ (.B(_1547_),
    .C(_1554_),
    .A(_1545_),
    .Y(_1556_));
 sg13g2_a21oi_2 _4532_ (.B1(net629),
    .Y(_1557_),
    .A2(_1556_),
    .A1(_1555_));
 sg13g2_o21ai_1 _4533_ (.B1(_1526_),
    .Y(_1558_),
    .A1(net865),
    .A2(net632));
 sg13g2_a21oi_1 _4534_ (.A1(net778),
    .A2(net709),
    .Y(_1559_),
    .B1(net772));
 sg13g2_o21ai_1 _4535_ (.B1(_1559_),
    .Y(_0155_),
    .A1(_1557_),
    .A2(_1558_));
 sg13g2_and2_1 _4536_ (.A(_1553_),
    .B(_1555_),
    .X(_1560_));
 sg13g2_nor2_1 _4537_ (.A(\core.V[9] ),
    .B(\core.dV[9] ),
    .Y(_1561_));
 sg13g2_nand2_1 _4538_ (.Y(_1562_),
    .A(\core.V[9] ),
    .B(\core.dV[9] ));
 sg13g2_nand2b_1 _4539_ (.Y(_1563_),
    .B(_1562_),
    .A_N(_1561_));
 sg13g2_xnor2_1 _4540_ (.Y(_1564_),
    .A(_1560_),
    .B(_1563_));
 sg13g2_o21ai_1 _4541_ (.B1(_1526_),
    .Y(_1565_),
    .A1(\core.Vreset_q[9] ),
    .A2(net632));
 sg13g2_a21oi_1 _4542_ (.A1(net632),
    .A2(_1564_),
    .Y(_1566_),
    .B1(_1565_));
 sg13g2_a21oi_1 _4543_ (.A1(net778),
    .A2(net872),
    .Y(_1567_),
    .B1(_1566_));
 sg13g2_nand2_1 _4544_ (.Y(_0156_),
    .A(net791),
    .B(net873));
 sg13g2_and2_1 _4545_ (.A(\core.V[10] ),
    .B(\core.dV[10] ),
    .X(_1568_));
 sg13g2_xor2_1 _4546_ (.B(\core.dV[10] ),
    .A(\core.V[10] ),
    .X(_1569_));
 sg13g2_o21ai_1 _4547_ (.B1(_1562_),
    .Y(_1570_),
    .A1(_1560_),
    .A2(_1561_));
 sg13g2_xnor2_1 _4548_ (.Y(_1571_),
    .A(_1569_),
    .B(_1570_));
 sg13g2_o21ai_1 _4549_ (.B1(_1526_),
    .Y(_1572_),
    .A1(\core.Vreset_q[10] ),
    .A2(net632));
 sg13g2_a21oi_1 _4550_ (.A1(net632),
    .A2(_1571_),
    .Y(_1573_),
    .B1(_1572_));
 sg13g2_a21oi_1 _4551_ (.A1(net778),
    .A2(net861),
    .Y(_1574_),
    .B1(_1573_));
 sg13g2_nor2_1 _4552_ (.A(net771),
    .B(net862),
    .Y(_0157_));
 sg13g2_a21o_1 _4553_ (.A2(net630),
    .A1(_0008_),
    .B1(_1525_),
    .X(_1575_));
 sg13g2_nor2_1 _4554_ (.A(_1496_),
    .B(_1575_),
    .Y(_1576_));
 sg13g2_a21o_1 _4555_ (.A2(_1570_),
    .A1(_1569_),
    .B1(_1568_),
    .X(_1577_));
 sg13g2_xnor2_1 _4556_ (.Y(_1578_),
    .A(\core.V[11] ),
    .B(\core.dV[11] ));
 sg13g2_a21oi_1 _4557_ (.A1(_1577_),
    .A2(_1578_),
    .Y(_1579_),
    .B1(net629));
 sg13g2_o21ai_1 _4558_ (.B1(_1579_),
    .Y(_1580_),
    .A1(_1577_),
    .A2(_1578_));
 sg13g2_a22oi_1 _4559_ (.Y(_1581_),
    .B1(_1576_),
    .B2(_1580_),
    .A2(net875),
    .A1(net778));
 sg13g2_nand2_1 _4560_ (.Y(_0158_),
    .A(net791),
    .B(net876));
 sg13g2_nand2_1 _4561_ (.Y(_1582_),
    .A(\core.V[12] ),
    .B(\core.dV[12] ));
 sg13g2_xnor2_1 _4562_ (.Y(_1583_),
    .A(\core.V[12] ),
    .B(\core.dV[12] ));
 sg13g2_a21o_1 _4563_ (.A2(\core.dV[11] ),
    .A1(\core.V[11] ),
    .B1(_1577_),
    .X(_1584_));
 sg13g2_o21ai_1 _4564_ (.B1(_1584_),
    .Y(_1585_),
    .A1(\core.V[11] ),
    .A2(\core.dV[11] ));
 sg13g2_xnor2_1 _4565_ (.Y(_1586_),
    .A(_1583_),
    .B(_1585_));
 sg13g2_nand2_1 _4566_ (.Y(_1587_),
    .A(net632),
    .B(_1586_));
 sg13g2_a22oi_1 _4567_ (.Y(_1588_),
    .B1(_1576_),
    .B2(_1587_),
    .A2(net846),
    .A1(net778));
 sg13g2_nand2_1 _4568_ (.Y(_0159_),
    .A(net791),
    .B(net847));
 sg13g2_nor2_1 _4569_ (.A(net783),
    .B(net863),
    .Y(_1589_));
 sg13g2_o21ai_1 _4570_ (.B1(_1582_),
    .Y(_1590_),
    .A1(_1583_),
    .A2(_1585_));
 sg13g2_nor2_1 _4571_ (.A(\core.V[13] ),
    .B(\core.dV[13] ),
    .Y(_1591_));
 sg13g2_and2_1 _4572_ (.A(\core.V[13] ),
    .B(\core.dV[13] ),
    .X(_1592_));
 sg13g2_o21ai_1 _4573_ (.B1(_1590_),
    .Y(_1593_),
    .A1(_1591_),
    .A2(_1592_));
 sg13g2_nor3_1 _4574_ (.A(_1590_),
    .B(_1591_),
    .C(_1592_),
    .Y(_1594_));
 sg13g2_nor2_1 _4575_ (.A(net629),
    .B(_1594_),
    .Y(_1595_));
 sg13g2_a21oi_1 _4576_ (.A1(_1593_),
    .A2(_1595_),
    .Y(_1596_),
    .B1(_1575_));
 sg13g2_nor2_1 _4577_ (.A(_1496_),
    .B(_1596_),
    .Y(_1597_));
 sg13g2_o21ai_1 _4578_ (.B1(net793),
    .Y(_0160_),
    .A1(_1589_),
    .A2(_1597_));
 sg13g2_a21oi_1 _4579_ (.A1(net778),
    .A2(\core.V[14] ),
    .Y(_1598_),
    .B1(net772));
 sg13g2_xnor2_1 _4580_ (.Y(_1599_),
    .A(\core.V[14] ),
    .B(\core.dV[14] ));
 sg13g2_nor2_1 _4581_ (.A(_1590_),
    .B(_1592_),
    .Y(_1600_));
 sg13g2_o21ai_1 _4582_ (.B1(_1599_),
    .Y(_1601_),
    .A1(_1591_),
    .A2(_1600_));
 sg13g2_nor3_1 _4583_ (.A(_1591_),
    .B(_1599_),
    .C(_1600_),
    .Y(_1602_));
 sg13g2_nor2_1 _4584_ (.A(net629),
    .B(_1602_),
    .Y(_1603_));
 sg13g2_a221oi_1 _4585_ (.B2(_1603_),
    .C1(_1525_),
    .B1(_1601_),
    .A1(net858),
    .Y(_1604_),
    .A2(net630));
 sg13g2_o21ai_1 _4586_ (.B1(_1598_),
    .Y(_0161_),
    .A1(_1496_),
    .A2(_1604_));
 sg13g2_a21oi_1 _4587_ (.A1(\core.V[14] ),
    .A2(\core.dV[14] ),
    .Y(_1605_),
    .B1(_1602_));
 sg13g2_xor2_1 _4588_ (.B(\core.dV[15] ),
    .A(\core.V[15] ),
    .X(_1606_));
 sg13g2_o21ai_1 _4589_ (.B1(net632),
    .Y(_1607_),
    .A1(_1605_),
    .A2(_1606_));
 sg13g2_a21oi_1 _4590_ (.A1(_1605_),
    .A2(_1606_),
    .Y(_1608_),
    .B1(_1607_));
 sg13g2_nor2_1 _4591_ (.A(_1575_),
    .B(_1608_),
    .Y(_1609_));
 sg13g2_o21ai_1 _4592_ (.B1(net783),
    .Y(_1610_),
    .A1(_1495_),
    .A2(_1609_));
 sg13g2_o21ai_1 _4593_ (.B1(_1610_),
    .Y(_0162_),
    .A1(net681),
    .A2(_2193_));
 sg13g2_a21o_2 _4594_ (.A2(net630),
    .A1(_1990_),
    .B1(net779),
    .X(_1611_));
 sg13g2_a22oi_1 _4595_ (.Y(_1612_),
    .B1(_1611_),
    .B2(net708),
    .A2(_2086_),
    .A1(_2019_));
 sg13g2_o21ai_1 _4596_ (.B1(net792),
    .Y(_1613_),
    .A1(net708),
    .A2(net472));
 sg13g2_nor2_1 _4597_ (.A(_1612_),
    .B(_1613_),
    .Y(_0163_));
 sg13g2_xor2_1 _4598_ (.B(_2020_),
    .A(_2019_),
    .X(_1614_));
 sg13g2_a22oi_1 _4599_ (.Y(_1615_),
    .B1(_1614_),
    .B2(_2086_),
    .A2(_1611_),
    .A1(net867));
 sg13g2_nor2_1 _4600_ (.A(net771),
    .B(_1615_),
    .Y(_0164_));
 sg13g2_xor2_1 _4601_ (.B(_2022_),
    .A(_2018_),
    .X(_1616_));
 sg13g2_a22oi_1 _4602_ (.Y(_1617_),
    .B1(_1616_),
    .B2(_2086_),
    .A2(_1611_),
    .A1(net870));
 sg13g2_nor2_1 _4603_ (.A(net771),
    .B(net871),
    .Y(_0165_));
 sg13g2_nand2b_1 _4604_ (.Y(_1618_),
    .B(_2024_),
    .A_N(_2025_));
 sg13g2_and3_1 _4605_ (.X(_1619_),
    .A(_1990_),
    .B(_2026_),
    .C(_1618_));
 sg13g2_o21ai_1 _4606_ (.B1(net792),
    .Y(_1620_),
    .A1(_1611_),
    .A2(_1619_));
 sg13g2_a21oi_1 _4607_ (.A1(_1919_),
    .A2(_1611_),
    .Y(_0166_),
    .B1(_1620_));
 sg13g2_nor3_2 _4608_ (.A(_1957_),
    .B(net607),
    .C(net707),
    .Y(_1621_));
 sg13g2_o21ai_1 _4609_ (.B1(net804),
    .Y(_1622_),
    .A1(_0016_),
    .A2(_1621_));
 sg13g2_nor2_1 _4610_ (.A(\core.watchdog_cnt[4] ),
    .B(net400),
    .Y(_1623_));
 sg13g2_nand2b_1 _4611_ (.Y(_1624_),
    .B(\core.watchdog_cnt[6] ),
    .A_N(\core.watchdog_cnt[7] ));
 sg13g2_o21ai_1 _4612_ (.B1(_0019_),
    .Y(_1625_),
    .A1(_1623_),
    .A2(_1624_));
 sg13g2_nand3_1 _4613_ (.B(\core.watchdog_cnt[8] ),
    .C(_1625_),
    .A(\core.watchdog_cnt[9] ),
    .Y(_1626_));
 sg13g2_nor4_2 _4614_ (.A(\core.watchdog_cnt[13] ),
    .B(\core.watchdog_cnt[12] ),
    .C(\core.watchdog_cnt[11] ),
    .Y(_1627_),
    .D(\core.watchdog_cnt[10] ));
 sg13g2_nand2_1 _4615_ (.Y(_1628_),
    .A(\core.watchdog_cnt[15] ),
    .B(\core.watchdog_cnt[14] ));
 sg13g2_a21oi_2 _4616_ (.B1(_1628_),
    .Y(_1629_),
    .A2(_1627_),
    .A1(_1626_));
 sg13g2_nor2_1 _4617_ (.A(net679),
    .B(_1629_),
    .Y(_1630_));
 sg13g2_nand3_1 _4618_ (.B(_1621_),
    .C(net641),
    .A(net4),
    .Y(_1631_));
 sg13g2_and3_1 _4619_ (.X(_1632_),
    .A(\core.lstate[0] ),
    .B(net707),
    .C(_0016_));
 sg13g2_and4_1 _4620_ (.A(net5),
    .B(net6),
    .C(net7),
    .D(net8),
    .X(_1633_));
 sg13g2_nand3_1 _4621_ (.B(_1632_),
    .C(_1633_),
    .A(_2161_),
    .Y(_1634_));
 sg13g2_nand2_1 _4622_ (.Y(_1635_),
    .A(net6),
    .B(net7));
 sg13g2_nand4_1 _4623_ (.B(net8),
    .C(_2161_),
    .A(net5),
    .Y(_1636_),
    .D(_1632_));
 sg13g2_nor2_1 _4624_ (.A(_1635_),
    .B(_1636_),
    .Y(_1637_));
 sg13g2_a21oi_1 _4625_ (.A1(_1631_),
    .A2(net676),
    .Y(_0167_),
    .B1(_1622_));
 sg13g2_and2_1 _4626_ (.A(net707),
    .B(_2158_),
    .X(_1638_));
 sg13g2_nand2_2 _4627_ (.Y(_1639_),
    .A(net707),
    .B(_2158_));
 sg13g2_nand3_1 _4628_ (.B(net592),
    .C(net554),
    .A(net560),
    .Y(_1640_));
 sg13g2_nand2b_1 _4629_ (.Y(_1641_),
    .B(net554),
    .A_N(net374));
 sg13g2_or2_1 _4630_ (.X(_1642_),
    .B(_1640_),
    .A(net591));
 sg13g2_and3_1 _4631_ (.X(_1643_),
    .A(net560),
    .B(net563),
    .C(_1638_));
 sg13g2_nor2_1 _4632_ (.A(_1639_),
    .B(_1642_),
    .Y(_1644_));
 sg13g2_or2_1 _4633_ (.X(_1645_),
    .B(_1642_),
    .A(_1639_));
 sg13g2_nand2_2 _4634_ (.Y(_1646_),
    .A(_2160_),
    .B(_1629_));
 sg13g2_inv_1 _4635_ (.Y(_1647_),
    .A(_1646_));
 sg13g2_nand2_1 _4636_ (.Y(_1648_),
    .A(\core.nibble_cnt ),
    .B(_2161_));
 sg13g2_nor3_2 _4637_ (.A(net707),
    .B(_2165_),
    .C(_1648_),
    .Y(_1649_));
 sg13g2_a22oi_1 _4638_ (.Y(_1650_),
    .B1(_1649_),
    .B2(net4),
    .A2(_1646_),
    .A1(_1961_));
 sg13g2_a22oi_1 _4639_ (.Y(_1651_),
    .B1(_1632_),
    .B2(_2162_),
    .A2(_1621_),
    .A1(net4));
 sg13g2_a22oi_1 _4640_ (.Y(_1652_),
    .B1(net677),
    .B2(net4),
    .A2(_2163_),
    .A1(net680));
 sg13g2_a21o_1 _4641_ (.A2(_1652_),
    .A1(_1651_),
    .B1(_1650_),
    .X(_1653_));
 sg13g2_a21oi_1 _4642_ (.A1(_1645_),
    .A2(_1653_),
    .Y(_0168_),
    .B1(_1622_));
 sg13g2_o21ai_1 _4643_ (.B1(net521),
    .Y(_1654_),
    .A1(_2160_),
    .A2(_2163_));
 sg13g2_nand3_1 _4644_ (.B(net677),
    .C(_1648_),
    .A(net4),
    .Y(_1655_));
 sg13g2_nand3_1 _4645_ (.B(_1651_),
    .C(_1655_),
    .A(_2160_),
    .Y(_1656_));
 sg13g2_nand3_1 _4646_ (.B(_1654_),
    .C(_1656_),
    .A(_1646_),
    .Y(_1657_));
 sg13g2_a21oi_1 _4647_ (.A1(_1639_),
    .A2(_1657_),
    .Y(_0169_),
    .B1(_1622_));
 sg13g2_nor2_2 _4648_ (.A(_2167_),
    .B(_1649_),
    .Y(_1658_));
 sg13g2_or2_1 _4649_ (.X(_1659_),
    .B(_1649_),
    .A(_2167_));
 sg13g2_a21oi_1 _4650_ (.A1(net5),
    .A2(net677),
    .Y(_1660_),
    .B1(_1659_));
 sg13g2_o21ai_1 _4651_ (.B1(net801),
    .Y(_1661_),
    .A1(net545),
    .A2(_1658_));
 sg13g2_nor2_1 _4652_ (.A(_1660_),
    .B(_1661_),
    .Y(_0170_));
 sg13g2_a21oi_1 _4653_ (.A1(net6),
    .A2(net677),
    .Y(_1662_),
    .B1(_1659_));
 sg13g2_o21ai_1 _4654_ (.B1(net801),
    .Y(_1663_),
    .A1(net577),
    .A2(_1658_));
 sg13g2_nor2_1 _4655_ (.A(_1662_),
    .B(_1663_),
    .Y(_0171_));
 sg13g2_a21oi_1 _4656_ (.A1(net7),
    .A2(net677),
    .Y(_1664_),
    .B1(_1659_));
 sg13g2_o21ai_1 _4657_ (.B1(net801),
    .Y(_1665_),
    .A1(net557),
    .A2(_1658_));
 sg13g2_nor2_1 _4658_ (.A(_1664_),
    .B(_1665_),
    .Y(_0172_));
 sg13g2_a21oi_1 _4659_ (.A1(net8),
    .A2(net677),
    .Y(_1666_),
    .B1(_1659_));
 sg13g2_o21ai_1 _4660_ (.B1(net801),
    .Y(_1667_),
    .A1(net562),
    .A2(_1658_));
 sg13g2_nor2_1 _4661_ (.A(_1666_),
    .B(_1667_),
    .Y(_0173_));
 sg13g2_nand3b_1 _4662_ (.B(_1638_),
    .C(net560),
    .Y(_1668_),
    .A_N(\core.param_idx[1] ));
 sg13g2_nor2_1 _4663_ (.A(_1641_),
    .B(_1668_),
    .Y(_1669_));
 sg13g2_o21ai_1 _4664_ (.B1(net784),
    .Y(_1670_),
    .A1(net481),
    .A2(net654));
 sg13g2_a21oi_1 _4665_ (.A1(_1861_),
    .A2(net654),
    .Y(_0174_),
    .B1(_1670_));
 sg13g2_o21ai_1 _4666_ (.B1(net800),
    .Y(_1671_),
    .A1(net601),
    .A2(net655));
 sg13g2_a21oi_1 _4667_ (.A1(_1860_),
    .A2(_1669_),
    .Y(_0175_),
    .B1(_1671_));
 sg13g2_o21ai_1 _4668_ (.B1(net785),
    .Y(_1672_),
    .A1(net419),
    .A2(net654));
 sg13g2_a21oi_1 _4669_ (.A1(_1858_),
    .A2(net654),
    .Y(_0176_),
    .B1(_1672_));
 sg13g2_o21ai_1 _4670_ (.B1(net787),
    .Y(_1673_),
    .A1(net359),
    .A2(net654));
 sg13g2_a21oi_1 _4671_ (.A1(_1857_),
    .A2(net654),
    .Y(_0177_),
    .B1(_1673_));
 sg13g2_o21ai_1 _4672_ (.B1(net786),
    .Y(_1674_),
    .A1(net361),
    .A2(net654));
 sg13g2_a21oi_1 _4673_ (.A1(_1856_),
    .A2(net655),
    .Y(_0178_),
    .B1(_1674_));
 sg13g2_o21ai_1 _4674_ (.B1(net786),
    .Y(_1675_),
    .A1(net349),
    .A2(net654));
 sg13g2_a21oi_1 _4675_ (.A1(_1855_),
    .A2(net655),
    .Y(_0179_),
    .B1(_1675_));
 sg13g2_o21ai_1 _4676_ (.B1(net800),
    .Y(_1676_),
    .A1(net479),
    .A2(net655));
 sg13g2_a21oi_1 _4677_ (.A1(_1853_),
    .A2(net655),
    .Y(_0180_),
    .B1(_1676_));
 sg13g2_o21ai_1 _4678_ (.B1(net800),
    .Y(_1677_),
    .A1(net549),
    .A2(net655));
 sg13g2_a21oi_1 _4679_ (.A1(_1851_),
    .A2(net655),
    .Y(_0181_),
    .B1(_1677_));
 sg13g2_o21ai_1 _4680_ (.B1(net785),
    .Y(_1678_),
    .A1(net448),
    .A2(net658));
 sg13g2_a21oi_1 _4681_ (.A1(_1861_),
    .A2(net658),
    .Y(_0182_),
    .B1(_1678_));
 sg13g2_o21ai_1 _4682_ (.B1(net800),
    .Y(_1679_),
    .A1(net599),
    .A2(_1644_));
 sg13g2_a21oi_1 _4683_ (.A1(_1860_),
    .A2(net659),
    .Y(_0183_),
    .B1(_1679_));
 sg13g2_o21ai_1 _4684_ (.B1(net786),
    .Y(_1680_),
    .A1(net451),
    .A2(net658));
 sg13g2_a21oi_1 _4685_ (.A1(_1858_),
    .A2(net658),
    .Y(_0184_),
    .B1(_1680_));
 sg13g2_o21ai_1 _4686_ (.B1(net786),
    .Y(_1681_),
    .A1(net546),
    .A2(net659));
 sg13g2_a21oi_1 _4687_ (.A1(_1857_),
    .A2(net659),
    .Y(_0185_),
    .B1(_1681_));
 sg13g2_o21ai_1 _4688_ (.B1(net786),
    .Y(_1682_),
    .A1(net484),
    .A2(net659));
 sg13g2_a21oi_1 _4689_ (.A1(_1856_),
    .A2(net658),
    .Y(_0186_),
    .B1(_1682_));
 sg13g2_o21ai_1 _4690_ (.B1(net786),
    .Y(_1683_),
    .A1(net535),
    .A2(net658));
 sg13g2_a21oi_1 _4691_ (.A1(_1855_),
    .A2(net659),
    .Y(_0187_),
    .B1(_1683_));
 sg13g2_o21ai_1 _4692_ (.B1(net800),
    .Y(_1684_),
    .A1(net461),
    .A2(net659));
 sg13g2_a21oi_1 _4693_ (.A1(_1853_),
    .A2(net659),
    .Y(_0188_),
    .B1(_1684_));
 sg13g2_o21ai_1 _4694_ (.B1(net786),
    .Y(_1685_),
    .A1(net434),
    .A2(net658));
 sg13g2_a21oi_1 _4695_ (.A1(_1851_),
    .A2(net658),
    .Y(_0189_),
    .B1(_1685_));
 sg13g2_o21ai_1 _4696_ (.B1(net806),
    .Y(_1686_),
    .A1(\core.p_TauW[0] ),
    .A2(net668));
 sg13g2_a21oi_1 _4697_ (.A1(_1880_),
    .A2(net668),
    .Y(_0190_),
    .B1(_1686_));
 sg13g2_o21ai_1 _4698_ (.B1(net805),
    .Y(_1687_),
    .A1(net369),
    .A2(net666));
 sg13g2_a21oi_1 _4699_ (.A1(_1879_),
    .A2(net665),
    .Y(_0191_),
    .B1(_1687_));
 sg13g2_nor2_1 _4700_ (.A(net582),
    .B(_1634_),
    .Y(_1688_));
 sg13g2_o21ai_1 _4701_ (.B1(net806),
    .Y(_1689_),
    .A1(\core.p_TauW[2] ),
    .A2(net668));
 sg13g2_nor2_1 _4702_ (.A(_1688_),
    .B(_1689_),
    .Y(_0192_));
 sg13g2_o21ai_1 _4703_ (.B1(net805),
    .Y(_1690_),
    .A1(\core.p_TauW[3] ),
    .A2(net668));
 sg13g2_a21oi_1 _4704_ (.A1(_1878_),
    .A2(net668),
    .Y(_0193_),
    .B1(_1690_));
 sg13g2_o21ai_1 _4705_ (.B1(net805),
    .Y(_1691_),
    .A1(\core.p_TauW[4] ),
    .A2(net669));
 sg13g2_a21oi_1 _4706_ (.A1(_1877_),
    .A2(net669),
    .Y(_0194_),
    .B1(_1691_));
 sg13g2_nor2_1 _4707_ (.A(net610),
    .B(_1634_),
    .Y(_1692_));
 sg13g2_o21ai_1 _4708_ (.B1(net806),
    .Y(_1693_),
    .A1(net813),
    .A2(net669));
 sg13g2_nor2_1 _4709_ (.A(_1692_),
    .B(_1693_),
    .Y(_0195_));
 sg13g2_nor2_1 _4710_ (.A(net452),
    .B(net676),
    .Y(_1694_));
 sg13g2_o21ai_1 _4711_ (.B1(net806),
    .Y(_1695_),
    .A1(\core.p_TauW[6] ),
    .A2(net669));
 sg13g2_nor2_1 _4712_ (.A(_1694_),
    .B(_1695_),
    .Y(_0196_));
 sg13g2_o21ai_1 _4713_ (.B1(net805),
    .Y(_1696_),
    .A1(\core.p_TauW[7] ),
    .A2(net668));
 sg13g2_a21oi_1 _4714_ (.A1(_1876_),
    .A2(net668),
    .Y(_0197_),
    .B1(_1696_));
 sg13g2_o21ai_1 _4715_ (.B1(net790),
    .Y(_1697_),
    .A1(\core.p_a[0] ),
    .A2(net664));
 sg13g2_a21oi_1 _4716_ (.A1(_1875_),
    .A2(net664),
    .Y(_0198_),
    .B1(_1697_));
 sg13g2_nor2_1 _4717_ (.A(net438),
    .B(net675),
    .Y(_1698_));
 sg13g2_o21ai_1 _4718_ (.B1(net789),
    .Y(_1699_),
    .A1(\core.p_a[1] ),
    .A2(net665));
 sg13g2_nor2_1 _4719_ (.A(_1698_),
    .B(_1699_),
    .Y(_0199_));
 sg13g2_o21ai_1 _4720_ (.B1(net790),
    .Y(_1700_),
    .A1(\core.p_a[2] ),
    .A2(net664));
 sg13g2_a21oi_1 _4721_ (.A1(_1874_),
    .A2(net664),
    .Y(_0200_),
    .B1(_1700_));
 sg13g2_o21ai_1 _4722_ (.B1(net788),
    .Y(_1701_),
    .A1(\core.p_a[3] ),
    .A2(net664));
 sg13g2_a21oi_1 _4723_ (.A1(_1873_),
    .A2(net664),
    .Y(_0201_),
    .B1(_1701_));
 sg13g2_o21ai_1 _4724_ (.B1(net788),
    .Y(_1702_),
    .A1(\core.p_a[4] ),
    .A2(net664));
 sg13g2_a21oi_1 _4725_ (.A1(_1872_),
    .A2(net667),
    .Y(_0202_),
    .B1(_1702_));
 sg13g2_o21ai_1 _4726_ (.B1(net788),
    .Y(_1703_),
    .A1(\core.p_a[5] ),
    .A2(net664));
 sg13g2_a21oi_1 _4727_ (.A1(_1871_),
    .A2(net667),
    .Y(_0203_),
    .B1(_1703_));
 sg13g2_o21ai_1 _4728_ (.B1(net789),
    .Y(_1704_),
    .A1(\core.p_a[6] ),
    .A2(net665));
 sg13g2_a21oi_1 _4729_ (.A1(_1870_),
    .A2(net665),
    .Y(_0204_),
    .B1(_1704_));
 sg13g2_o21ai_1 _4730_ (.B1(net793),
    .Y(_1705_),
    .A1(net351),
    .A2(net666));
 sg13g2_a21oi_1 _4731_ (.A1(_1869_),
    .A2(net666),
    .Y(_0205_),
    .B1(_1705_));
 sg13g2_o21ai_1 _4732_ (.B1(net808),
    .Y(_1706_),
    .A1(net388),
    .A2(net672));
 sg13g2_a21oi_1 _4733_ (.A1(_1868_),
    .A2(net671),
    .Y(_0206_),
    .B1(_1706_));
 sg13g2_o21ai_1 _4734_ (.B1(net807),
    .Y(_1707_),
    .A1(\core.p_b[1] ),
    .A2(net671));
 sg13g2_a21oi_1 _4735_ (.A1(_1867_),
    .A2(net671),
    .Y(_0207_),
    .B1(_1707_));
 sg13g2_o21ai_1 _4736_ (.B1(net807),
    .Y(_1708_),
    .A1(\core.p_b[2] ),
    .A2(net671));
 sg13g2_a21oi_1 _4737_ (.A1(_1866_),
    .A2(net671),
    .Y(_0208_),
    .B1(_1708_));
 sg13g2_o21ai_1 _4738_ (.B1(net807),
    .Y(_1709_),
    .A1(\core.p_b[3] ),
    .A2(net671));
 sg13g2_a21oi_1 _4739_ (.A1(_1865_),
    .A2(net671),
    .Y(_0209_),
    .B1(_1709_));
 sg13g2_o21ai_1 _4740_ (.B1(net802),
    .Y(_1710_),
    .A1(\core.p_b[4] ),
    .A2(net671));
 sg13g2_a21oi_1 _4741_ (.A1(_1864_),
    .A2(net673),
    .Y(_0210_),
    .B1(_1710_));
 sg13g2_nor2_1 _4742_ (.A(net594),
    .B(net676),
    .Y(_1711_));
 sg13g2_o21ai_1 _4743_ (.B1(net809),
    .Y(_1712_),
    .A1(net600),
    .A2(net672));
 sg13g2_nor2_1 _4744_ (.A(_1711_),
    .B(_1712_),
    .Y(_0211_));
 sg13g2_o21ai_1 _4745_ (.B1(net801),
    .Y(_1713_),
    .A1(\core.p_b[6] ),
    .A2(net672));
 sg13g2_a21oi_1 _4746_ (.A1(_1863_),
    .A2(net673),
    .Y(_0212_),
    .B1(_1713_));
 sg13g2_o21ai_1 _4747_ (.B1(net801),
    .Y(_1714_),
    .A1(\core.p_b[7] ),
    .A2(net672));
 sg13g2_a21oi_1 _4748_ (.A1(_1862_),
    .A2(net673),
    .Y(_0213_),
    .B1(_1714_));
 sg13g2_nor2_1 _4749_ (.A(net523),
    .B(net676),
    .Y(_1715_));
 sg13g2_o21ai_1 _4750_ (.B1(net796),
    .Y(_1716_),
    .A1(\core.p_Vreset[0] ),
    .A2(net665));
 sg13g2_nor2_1 _4751_ (.A(_1715_),
    .B(_1716_),
    .Y(_0214_));
 sg13g2_o21ai_1 _4752_ (.B1(net796),
    .Y(_1717_),
    .A1(\core.p_Vreset[1] ),
    .A2(net665));
 sg13g2_a21oi_1 _4753_ (.A1(_1859_),
    .A2(net665),
    .Y(_0215_),
    .B1(_1717_));
 sg13g2_nor2_1 _4754_ (.A(net555),
    .B(net676),
    .Y(_1718_));
 sg13g2_o21ai_1 _4755_ (.B1(net806),
    .Y(_1719_),
    .A1(net527),
    .A2(net668));
 sg13g2_nor2_1 _4756_ (.A(_1718_),
    .B(_1719_),
    .Y(_0216_));
 sg13g2_nor2_1 _4757_ (.A(net579),
    .B(net675),
    .Y(_1720_));
 sg13g2_o21ai_1 _4758_ (.B1(net805),
    .Y(_1721_),
    .A1(\core.p_Vreset[3] ),
    .A2(net666));
 sg13g2_nor2_1 _4759_ (.A(_1720_),
    .B(_1721_),
    .Y(_0217_));
 sg13g2_nor2_1 _4760_ (.A(net449),
    .B(net676),
    .Y(_1722_));
 sg13g2_o21ai_1 _4761_ (.B1(net796),
    .Y(_1723_),
    .A1(\core.p_Vreset[4] ),
    .A2(net670));
 sg13g2_nor2_1 _4762_ (.A(_1722_),
    .B(_1723_),
    .Y(_0218_));
 sg13g2_o21ai_1 _4763_ (.B1(net796),
    .Y(_1724_),
    .A1(\core.p_Vreset[5] ),
    .A2(net670));
 sg13g2_a21oi_1 _4764_ (.A1(_1854_),
    .A2(net670),
    .Y(_0219_),
    .B1(_1724_));
 sg13g2_o21ai_1 _4765_ (.B1(net798),
    .Y(_1725_),
    .A1(\core.p_Vreset[6] ),
    .A2(net670));
 sg13g2_a21oi_1 _4766_ (.A1(_1852_),
    .A2(net670),
    .Y(_0220_),
    .B1(_1725_));
 sg13g2_nor2_1 _4767_ (.A(\core.s_Vreset[7] ),
    .B(net675),
    .Y(_1726_));
 sg13g2_o21ai_1 _4768_ (.B1(net795),
    .Y(_1727_),
    .A1(net519),
    .A2(net665));
 sg13g2_nor2_1 _4769_ (.A(_1726_),
    .B(_1727_),
    .Y(_0221_));
 sg13g2_o21ai_1 _4770_ (.B1(net785),
    .Y(_1728_),
    .A1(net404),
    .A2(net662));
 sg13g2_a21oi_1 _4771_ (.A1(_1899_),
    .A2(net662),
    .Y(_0222_),
    .B1(_1728_));
 sg13g2_nor2_1 _4772_ (.A(net601),
    .B(net675),
    .Y(_1729_));
 sg13g2_o21ai_1 _4773_ (.B1(net789),
    .Y(_1730_),
    .A1(\core.p_VT[1] ),
    .A2(net663));
 sg13g2_nor2_1 _4774_ (.A(_1729_),
    .B(_1730_),
    .Y(_0223_));
 sg13g2_o21ai_1 _4775_ (.B1(net788),
    .Y(_1731_),
    .A1(\core.p_VT[2] ),
    .A2(net662));
 sg13g2_a21oi_1 _4776_ (.A1(_1897_),
    .A2(net662),
    .Y(_0224_),
    .B1(_1731_));
 sg13g2_o21ai_1 _4777_ (.B1(net784),
    .Y(_1732_),
    .A1(\core.p_VT[3] ),
    .A2(net662));
 sg13g2_a21oi_1 _4778_ (.A1(_1896_),
    .A2(net662),
    .Y(_0225_),
    .B1(_1732_));
 sg13g2_o21ai_1 _4779_ (.B1(net787),
    .Y(_1733_),
    .A1(\core.p_VT[4] ),
    .A2(net662));
 sg13g2_a21oi_1 _4780_ (.A1(_1895_),
    .A2(net663),
    .Y(_0226_),
    .B1(_1733_));
 sg13g2_o21ai_1 _4781_ (.B1(net787),
    .Y(_1734_),
    .A1(\core.p_VT[5] ),
    .A2(net663));
 sg13g2_a21oi_1 _4782_ (.A1(_1893_),
    .A2(net663),
    .Y(_0227_),
    .B1(_1734_));
 sg13g2_nor2_1 _4783_ (.A(net479),
    .B(net675),
    .Y(_1735_));
 sg13g2_o21ai_1 _4784_ (.B1(net795),
    .Y(_1736_),
    .A1(\core.p_VT[6] ),
    .A2(net663));
 sg13g2_nor2_1 _4785_ (.A(_1735_),
    .B(_1736_),
    .Y(_0228_));
 sg13g2_nor2_1 _4786_ (.A(\core.s_VT[7] ),
    .B(net675),
    .Y(_1737_));
 sg13g2_o21ai_1 _4787_ (.B1(net789),
    .Y(_1738_),
    .A1(net543),
    .A2(net663));
 sg13g2_nor2_1 _4788_ (.A(_1737_),
    .B(_1738_),
    .Y(_0229_));
 sg13g2_o21ai_1 _4789_ (.B1(net785),
    .Y(_1739_),
    .A1(net429),
    .A2(net661));
 sg13g2_a21oi_1 _4790_ (.A1(_1891_),
    .A2(net661),
    .Y(_0230_),
    .B1(_1739_));
 sg13g2_o21ai_1 _4791_ (.B1(net784),
    .Y(_1740_),
    .A1(net409),
    .A2(net661));
 sg13g2_a21oi_1 _4792_ (.A1(_1889_),
    .A2(net660),
    .Y(_0231_),
    .B1(_1740_));
 sg13g2_o21ai_1 _4793_ (.B1(net784),
    .Y(_1741_),
    .A1(net423),
    .A2(net661));
 sg13g2_a21oi_1 _4794_ (.A1(_1887_),
    .A2(net660),
    .Y(_0232_),
    .B1(_1741_));
 sg13g2_nor2_1 _4795_ (.A(net546),
    .B(net675),
    .Y(_1742_));
 sg13g2_o21ai_1 _4796_ (.B1(net784),
    .Y(_1743_),
    .A1(net576),
    .A2(net661));
 sg13g2_nor2_1 _4797_ (.A(_1742_),
    .B(_1743_),
    .Y(_0233_));
 sg13g2_o21ai_1 _4798_ (.B1(net784),
    .Y(_1744_),
    .A1(net456),
    .A2(net660));
 sg13g2_a21oi_1 _4799_ (.A1(_1885_),
    .A2(net660),
    .Y(_0234_),
    .B1(_1744_));
 sg13g2_o21ai_1 _4800_ (.B1(net784),
    .Y(_1745_),
    .A1(net445),
    .A2(net660));
 sg13g2_a21oi_1 _4801_ (.A1(_1883_),
    .A2(net660),
    .Y(_0235_),
    .B1(_1745_));
 sg13g2_nor2_1 _4802_ (.A(net461),
    .B(net675),
    .Y(_1746_));
 sg13g2_o21ai_1 _4803_ (.B1(net786),
    .Y(_1747_),
    .A1(\core.p_C[6] ),
    .A2(net663));
 sg13g2_nor2_1 _4804_ (.A(_1746_),
    .B(_1747_),
    .Y(_0236_));
 sg13g2_o21ai_1 _4805_ (.B1(net784),
    .Y(_1748_),
    .A1(\core.p_C[7] ),
    .A2(net660));
 sg13g2_a21oi_1 _4806_ (.A1(_1881_),
    .A2(net660),
    .Y(_0237_),
    .B1(_1748_));
 sg13g2_nand2_1 _4807_ (.Y(_1749_),
    .A(net706),
    .B(_2160_));
 sg13g2_a21oi_1 _4808_ (.A1(net676),
    .A2(_1749_),
    .Y(_0238_),
    .B1(net777));
 sg13g2_a22oi_1 _4809_ (.Y(_1750_),
    .B1(_1646_),
    .B2(net406),
    .A2(_2168_),
    .A1(net4));
 sg13g2_nand3b_1 _4810_ (.B(_0016_),
    .C(_1652_),
    .Y(_1751_),
    .A_N(net707));
 sg13g2_o21ai_1 _4811_ (.B1(_1751_),
    .Y(_1752_),
    .A1(_0017_),
    .A2(_2167_));
 sg13g2_nor3_1 _4812_ (.A(net774),
    .B(net407),
    .C(_1752_),
    .Y(_0239_));
 sg13g2_o21ai_1 _4813_ (.B1(_1652_),
    .Y(_1753_),
    .A1(_2158_),
    .A2(net677));
 sg13g2_nand2_1 _4814_ (.Y(_1754_),
    .A(_1646_),
    .B(_1753_));
 sg13g2_o21ai_1 _4815_ (.B1(_1754_),
    .Y(_1755_),
    .A1(_1645_),
    .A2(_1647_));
 sg13g2_inv_1 _4816_ (.Y(_1756_),
    .A(_1755_));
 sg13g2_nand2_1 _4817_ (.Y(_1757_),
    .A(\core.param_idx[0] ),
    .B(_1755_));
 sg13g2_nand3_1 _4818_ (.B(_1638_),
    .C(_1642_),
    .A(net346),
    .Y(_1758_));
 sg13g2_a21oi_1 _4819_ (.A1(_1757_),
    .A2(net347),
    .Y(_0240_),
    .B1(net777));
 sg13g2_nand3b_1 _4820_ (.B(net563),
    .C(_1638_),
    .Y(_1759_),
    .A_N(net825));
 sg13g2_nand2_1 _4821_ (.Y(_1760_),
    .A(net564),
    .B(_1759_));
 sg13g2_a21oi_1 _4822_ (.A1(net563),
    .A2(_1755_),
    .Y(_1761_),
    .B1(_1760_));
 sg13g2_nor2_1 _4823_ (.A(net777),
    .B(_1761_),
    .Y(_0241_));
 sg13g2_nand2_1 _4824_ (.Y(_1762_),
    .A(_1638_),
    .B(_1640_));
 sg13g2_o21ai_1 _4825_ (.B1(net800),
    .Y(_1763_),
    .A1(net554),
    .A2(_1643_));
 sg13g2_a21oi_1 _4826_ (.A1(_1756_),
    .A2(_1762_),
    .Y(_0242_),
    .B1(_1763_));
 sg13g2_nand2_1 _4827_ (.Y(_1764_),
    .A(net374),
    .B(net800));
 sg13g2_a21oi_1 _4828_ (.A1(_1754_),
    .A2(_1762_),
    .Y(_0243_),
    .B1(_1764_));
 sg13g2_nand2_1 _4829_ (.Y(_1765_),
    .A(net804),
    .B(_2167_));
 sg13g2_nand2_1 _4830_ (.Y(_1766_),
    .A(net852),
    .B(_2160_));
 sg13g2_o21ai_1 _4831_ (.B1(_1766_),
    .Y(_1767_),
    .A1(net852),
    .A2(net642));
 sg13g2_nor2_1 _4832_ (.A(net640),
    .B(_1767_),
    .Y(_0244_));
 sg13g2_nand2b_2 _4833_ (.Y(_1768_),
    .B(_1646_),
    .A_N(net639));
 sg13g2_nand2_1 _4834_ (.Y(_1769_),
    .A(\core.watchdog_cnt[0] ),
    .B(\core.watchdog_cnt[1] ));
 sg13g2_xor2_1 _4835_ (.B(_1766_),
    .A(net831),
    .X(_1770_));
 sg13g2_nor2_1 _4836_ (.A(_1768_),
    .B(net832),
    .Y(_0245_));
 sg13g2_xor2_1 _4837_ (.B(_1769_),
    .A(_0009_),
    .X(_1771_));
 sg13g2_a22oi_1 _4838_ (.Y(_1772_),
    .B1(net642),
    .B2(_1771_),
    .A2(net680),
    .A1(net517));
 sg13g2_nor2_1 _4839_ (.A(net639),
    .B(net518),
    .Y(_0246_));
 sg13g2_nand4_1 _4840_ (.B(\core.watchdog_cnt[1] ),
    .C(net517),
    .A(\core.watchdog_cnt[0] ),
    .Y(_1773_),
    .D(_2160_));
 sg13g2_nand4_1 _4841_ (.B(\core.watchdog_cnt[1] ),
    .C(net517),
    .A(\core.watchdog_cnt[0] ),
    .Y(_1774_),
    .D(\core.watchdog_cnt[3] ));
 sg13g2_inv_1 _4842_ (.Y(_1775_),
    .A(_1774_));
 sg13g2_xor2_1 _4843_ (.B(_1773_),
    .A(net595),
    .X(_1776_));
 sg13g2_nor2_1 _4844_ (.A(_1768_),
    .B(net596),
    .Y(_0247_));
 sg13g2_xor2_1 _4845_ (.B(_1774_),
    .A(_0010_),
    .X(_1777_));
 sg13g2_a22oi_1 _4846_ (.Y(_1778_),
    .B1(net641),
    .B2(_1777_),
    .A2(net680),
    .A1(net525));
 sg13g2_nor2_1 _4847_ (.A(net639),
    .B(net526),
    .Y(_0248_));
 sg13g2_nand3_1 _4848_ (.B(\core.watchdog_cnt[5] ),
    .C(_1775_),
    .A(\core.watchdog_cnt[4] ),
    .Y(_1779_));
 sg13g2_nor2_1 _4849_ (.A(net679),
    .B(_1779_),
    .Y(_1780_));
 sg13g2_a21oi_1 _4850_ (.A1(_2160_),
    .A2(_1775_),
    .Y(_1781_),
    .B1(net400));
 sg13g2_nor4_1 _4851_ (.A(_1623_),
    .B(_1768_),
    .C(_1780_),
    .D(net401),
    .Y(_0249_));
 sg13g2_nor2_1 _4852_ (.A(_0011_),
    .B(_1779_),
    .Y(_1782_));
 sg13g2_xor2_1 _4853_ (.B(_1779_),
    .A(_0011_),
    .X(_1783_));
 sg13g2_a22oi_1 _4854_ (.Y(_1784_),
    .B1(net642),
    .B2(_1783_),
    .A2(net679),
    .A1(net586));
 sg13g2_nor2_1 _4855_ (.A(net640),
    .B(net587),
    .Y(_0250_));
 sg13g2_xnor2_1 _4856_ (.Y(_1785_),
    .A(_0019_),
    .B(_1782_));
 sg13g2_a22oi_1 _4857_ (.Y(_1786_),
    .B1(net642),
    .B2(_1785_),
    .A2(net679),
    .A1(net540));
 sg13g2_nor2_1 _4858_ (.A(net640),
    .B(net541),
    .Y(_0251_));
 sg13g2_nand3_1 _4859_ (.B(net586),
    .C(_1780_),
    .A(net540),
    .Y(_1787_));
 sg13g2_nand3_1 _4860_ (.B(\core.watchdog_cnt[7] ),
    .C(\core.watchdog_cnt[6] ),
    .A(\core.watchdog_cnt[8] ),
    .Y(_1788_));
 sg13g2_nor2_1 _4861_ (.A(_1779_),
    .B(_1788_),
    .Y(_1789_));
 sg13g2_xor2_1 _4862_ (.B(_1787_),
    .A(net816),
    .X(_1790_));
 sg13g2_o21ai_1 _4863_ (.B1(_2160_),
    .Y(_1791_),
    .A1(_1629_),
    .A2(_1789_));
 sg13g2_nor2_1 _4864_ (.A(_1768_),
    .B(_1790_),
    .Y(_0252_));
 sg13g2_a21oi_1 _4865_ (.A1(net641),
    .A2(_1789_),
    .Y(_1792_),
    .B1(net477));
 sg13g2_nor2_1 _4866_ (.A(_1960_),
    .B(_1791_),
    .Y(_1793_));
 sg13g2_nor3_1 _4867_ (.A(net639),
    .B(net478),
    .C(_1793_),
    .Y(_0253_));
 sg13g2_nor3_2 _4868_ (.A(_1960_),
    .B(_1779_),
    .C(_1788_),
    .Y(_1794_));
 sg13g2_xnor2_1 _4869_ (.Y(_1795_),
    .A(net571),
    .B(_1794_));
 sg13g2_a22oi_1 _4870_ (.Y(_1796_),
    .B1(net641),
    .B2(_1795_),
    .A2(net679),
    .A1(\core.watchdog_cnt[10] ));
 sg13g2_nor2_1 _4871_ (.A(net639),
    .B(net572),
    .Y(_0254_));
 sg13g2_and3_1 _4872_ (.X(_1797_),
    .A(\core.watchdog_cnt[11] ),
    .B(\core.watchdog_cnt[10] ),
    .C(_1794_));
 sg13g2_nand3_1 _4873_ (.B(\core.watchdog_cnt[10] ),
    .C(_1794_),
    .A(\core.watchdog_cnt[11] ),
    .Y(_1798_));
 sg13g2_a21oi_1 _4874_ (.A1(\core.watchdog_cnt[10] ),
    .A2(_1794_),
    .Y(_1799_),
    .B1(net814));
 sg13g2_nor2_1 _4875_ (.A(_1797_),
    .B(_1799_),
    .Y(_1800_));
 sg13g2_a22oi_1 _4876_ (.Y(_1801_),
    .B1(net641),
    .B2(_1800_),
    .A2(net679),
    .A1(net814));
 sg13g2_nor2_1 _4877_ (.A(net639),
    .B(net815),
    .Y(_0255_));
 sg13g2_o21ai_1 _4878_ (.B1(net641),
    .Y(_1802_),
    .A1(net565),
    .A2(_1798_));
 sg13g2_a21oi_1 _4879_ (.A1(net565),
    .A2(_1798_),
    .Y(_1803_),
    .B1(_1802_));
 sg13g2_a21oi_1 _4880_ (.A1(\core.watchdog_cnt[12] ),
    .A2(net679),
    .Y(_1804_),
    .B1(net566));
 sg13g2_nor2_1 _4881_ (.A(net639),
    .B(net567),
    .Y(_0256_));
 sg13g2_a21oi_1 _4882_ (.A1(\core.watchdog_cnt[12] ),
    .A2(_1797_),
    .Y(_1805_),
    .B1(net608));
 sg13g2_nor2b_1 _4883_ (.A(_1805_),
    .B_N(net641),
    .Y(_1806_));
 sg13g2_nand3_1 _4884_ (.B(\core.watchdog_cnt[12] ),
    .C(_1797_),
    .A(\core.watchdog_cnt[13] ),
    .Y(_1807_));
 sg13g2_a22oi_1 _4885_ (.Y(_1808_),
    .B1(_1806_),
    .B2(_1807_),
    .A2(net679),
    .A1(net608));
 sg13g2_nor2_1 _4886_ (.A(net639),
    .B(net609),
    .Y(_0257_));
 sg13g2_o21ai_1 _4887_ (.B1(net641),
    .Y(_1809_),
    .A1(net506),
    .A2(_1807_));
 sg13g2_a21oi_1 _4888_ (.A1(net506),
    .A2(_1807_),
    .Y(_1810_),
    .B1(_1809_));
 sg13g2_a21oi_1 _4889_ (.A1(\core.watchdog_cnt[14] ),
    .A2(net680),
    .Y(_1811_),
    .B1(_1810_));
 sg13g2_nor2_1 _4890_ (.A(net640),
    .B(net507),
    .Y(_0258_));
 sg13g2_nor3_1 _4891_ (.A(_1959_),
    .B(net680),
    .C(_1807_),
    .Y(_1812_));
 sg13g2_nor2_1 _4892_ (.A(net459),
    .B(_1812_),
    .Y(_1813_));
 sg13g2_nor2_1 _4893_ (.A(_1768_),
    .B(net460),
    .Y(_0259_));
 sg13g2_nor2_1 _4894_ (.A(\core.param_idx[3] ),
    .B(\core.param_idx[2] ),
    .Y(_1814_));
 sg13g2_nor2b_1 _4895_ (.A(_1668_),
    .B_N(_1814_),
    .Y(_1815_));
 sg13g2_o21ai_1 _4896_ (.B1(net797),
    .Y(_1816_),
    .A1(net427),
    .A2(net652));
 sg13g2_a21oi_1 _4897_ (.A1(_1861_),
    .A2(net652),
    .Y(_0260_),
    .B1(_1816_));
 sg13g2_o21ai_1 _4898_ (.B1(net796),
    .Y(_1817_),
    .A1(net373),
    .A2(net653));
 sg13g2_a21oi_1 _4899_ (.A1(_1860_),
    .A2(net653),
    .Y(_0261_),
    .B1(_1817_));
 sg13g2_o21ai_1 _4900_ (.B1(net797),
    .Y(_1818_),
    .A1(net582),
    .A2(net651));
 sg13g2_a21oi_1 _4901_ (.A1(_1858_),
    .A2(net651),
    .Y(_0262_),
    .B1(_1818_));
 sg13g2_o21ai_1 _4902_ (.B1(net798),
    .Y(_1819_),
    .A1(net415),
    .A2(net653));
 sg13g2_a21oi_1 _4903_ (.A1(_1857_),
    .A2(net653),
    .Y(_0263_),
    .B1(_1819_));
 sg13g2_o21ai_1 _4904_ (.B1(net798),
    .Y(_1820_),
    .A1(net396),
    .A2(net652));
 sg13g2_a21oi_1 _4905_ (.A1(_1856_),
    .A2(net651),
    .Y(_0264_),
    .B1(_1820_));
 sg13g2_o21ai_1 _4906_ (.B1(net797),
    .Y(_1821_),
    .A1(net610),
    .A2(net651));
 sg13g2_a21oi_1 _4907_ (.A1(_1855_),
    .A2(net651),
    .Y(_0265_),
    .B1(_1821_));
 sg13g2_o21ai_1 _4908_ (.B1(net797),
    .Y(_1822_),
    .A1(net452),
    .A2(net651));
 sg13g2_a21oi_1 _4909_ (.A1(_1853_),
    .A2(net651),
    .Y(_0266_),
    .B1(_1822_));
 sg13g2_o21ai_1 _4910_ (.B1(net798),
    .Y(_1823_),
    .A1(net398),
    .A2(net651));
 sg13g2_a21oi_1 _4911_ (.A1(_1851_),
    .A2(net652),
    .Y(_0267_),
    .B1(_1823_));
 sg13g2_nor2b_1 _4912_ (.A(_1759_),
    .B_N(_1814_),
    .Y(_1824_));
 sg13g2_o21ai_1 _4913_ (.B1(net788),
    .Y(_1825_),
    .A1(net386),
    .A2(net649));
 sg13g2_a21oi_1 _4914_ (.A1(_1861_),
    .A2(net649),
    .Y(_0268_),
    .B1(_1825_));
 sg13g2_o21ai_1 _4915_ (.B1(net795),
    .Y(_1826_),
    .A1(net438),
    .A2(net650));
 sg13g2_a21oi_1 _4916_ (.A1(_1860_),
    .A2(net650),
    .Y(_0269_),
    .B1(_1826_));
 sg13g2_o21ai_1 _4917_ (.B1(net788),
    .Y(_1827_),
    .A1(net357),
    .A2(net649));
 sg13g2_a21oi_1 _4918_ (.A1(_1858_),
    .A2(net649),
    .Y(_0270_),
    .B1(_1827_));
 sg13g2_o21ai_1 _4919_ (.B1(net789),
    .Y(_1828_),
    .A1(net367),
    .A2(net649));
 sg13g2_a21oi_1 _4920_ (.A1(_1857_),
    .A2(net649),
    .Y(_0271_),
    .B1(_1828_));
 sg13g2_o21ai_1 _4921_ (.B1(net789),
    .Y(_1829_),
    .A1(net353),
    .A2(net650));
 sg13g2_a21oi_1 _4922_ (.A1(_1856_),
    .A2(net650),
    .Y(_0272_),
    .B1(_1829_));
 sg13g2_o21ai_1 _4923_ (.B1(net789),
    .Y(_1830_),
    .A1(net380),
    .A2(net649));
 sg13g2_a21oi_1 _4924_ (.A1(_1855_),
    .A2(net649),
    .Y(_0273_),
    .B1(_1830_));
 sg13g2_o21ai_1 _4925_ (.B1(net795),
    .Y(_1831_),
    .A1(net355),
    .A2(net650));
 sg13g2_a21oi_1 _4926_ (.A1(_1853_),
    .A2(net650),
    .Y(_0274_),
    .B1(_1831_));
 sg13g2_o21ai_1 _4927_ (.B1(net789),
    .Y(_1832_),
    .A1(net352),
    .A2(_1824_));
 sg13g2_a21oi_1 _4928_ (.A1(_1851_),
    .A2(net650),
    .Y(_0275_),
    .B1(_1832_));
 sg13g2_and2_1 _4929_ (.A(_1643_),
    .B(_1814_),
    .X(_1833_));
 sg13g2_o21ai_1 _4930_ (.B1(net803),
    .Y(_1834_),
    .A1(net403),
    .A2(net648));
 sg13g2_a21oi_1 _4931_ (.A1(_1861_),
    .A2(_1833_),
    .Y(_0276_),
    .B1(_1834_));
 sg13g2_o21ai_1 _4932_ (.B1(net802),
    .Y(_1835_),
    .A1(net363),
    .A2(net647));
 sg13g2_a21oi_1 _4933_ (.A1(_1860_),
    .A2(net647),
    .Y(_0277_),
    .B1(_1835_));
 sg13g2_o21ai_1 _4934_ (.B1(net802),
    .Y(_1836_),
    .A1(net425),
    .A2(net647));
 sg13g2_a21oi_1 _4935_ (.A1(_1858_),
    .A2(net647),
    .Y(_0278_),
    .B1(_1836_));
 sg13g2_o21ai_1 _4936_ (.B1(net803),
    .Y(_1837_),
    .A1(net496),
    .A2(net647));
 sg13g2_a21oi_1 _4937_ (.A1(_1857_),
    .A2(net647),
    .Y(_0279_),
    .B1(_1837_));
 sg13g2_o21ai_1 _4938_ (.B1(net802),
    .Y(_1838_),
    .A1(net376),
    .A2(net647));
 sg13g2_a21oi_1 _4939_ (.A1(_1856_),
    .A2(net647),
    .Y(_0280_),
    .B1(_1838_));
 sg13g2_o21ai_1 _4940_ (.B1(net801),
    .Y(_1839_),
    .A1(net594),
    .A2(net648));
 sg13g2_a21oi_1 _4941_ (.A1(_1855_),
    .A2(net648),
    .Y(_0281_),
    .B1(_1839_));
 sg13g2_o21ai_1 _4942_ (.B1(net801),
    .Y(_1840_),
    .A1(net390),
    .A2(net648));
 sg13g2_a21oi_1 _4943_ (.A1(_1853_),
    .A2(net648),
    .Y(_0282_),
    .B1(_1840_));
 sg13g2_o21ai_1 _4944_ (.B1(net803),
    .Y(_1841_),
    .A1(net392),
    .A2(net648));
 sg13g2_a21oi_1 _4945_ (.A1(_1851_),
    .A2(net648),
    .Y(_0283_),
    .B1(_1841_));
 sg13g2_nor4_1 _4946_ (.A(\core.param_idx[0] ),
    .B(\core.param_idx[1] ),
    .C(_1639_),
    .D(_1641_),
    .Y(_1842_));
 sg13g2_o21ai_1 _4947_ (.B1(net795),
    .Y(_1843_),
    .A1(net523),
    .A2(net656));
 sg13g2_a21oi_1 _4948_ (.A1(_1861_),
    .A2(net656),
    .Y(_0284_),
    .B1(_1843_));
 sg13g2_o21ai_1 _4949_ (.B1(net795),
    .Y(_1844_),
    .A1(net378),
    .A2(net656));
 sg13g2_a21oi_1 _4950_ (.A1(_1860_),
    .A2(net656),
    .Y(_0285_),
    .B1(_1844_));
 sg13g2_o21ai_1 _4951_ (.B1(net797),
    .Y(_1845_),
    .A1(net555),
    .A2(net657));
 sg13g2_a21oi_1 _4952_ (.A1(_1858_),
    .A2(net657),
    .Y(_0286_),
    .B1(_1845_));
 sg13g2_o21ai_1 _4953_ (.B1(net795),
    .Y(_1846_),
    .A1(net579),
    .A2(net656));
 sg13g2_a21oi_1 _4954_ (.A1(_1857_),
    .A2(net656),
    .Y(_0287_),
    .B1(_1846_));
 sg13g2_o21ai_1 _4955_ (.B1(net797),
    .Y(_1847_),
    .A1(net449),
    .A2(net657));
 sg13g2_a21oi_1 _4956_ (.A1(_1856_),
    .A2(net657),
    .Y(_0288_),
    .B1(_1847_));
 sg13g2_o21ai_1 _4957_ (.B1(net797),
    .Y(_1848_),
    .A1(net371),
    .A2(net657));
 sg13g2_a21oi_1 _4958_ (.A1(_1855_),
    .A2(net657),
    .Y(_0289_),
    .B1(_1848_));
 sg13g2_o21ai_1 _4959_ (.B1(net797),
    .Y(_1849_),
    .A1(net365),
    .A2(net657));
 sg13g2_a21oi_1 _4960_ (.A1(_1853_),
    .A2(net657),
    .Y(_0290_),
    .B1(_1849_));
 sg13g2_o21ai_1 _4961_ (.B1(net795),
    .Y(_1850_),
    .A1(net590),
    .A2(net656));
 sg13g2_a21oi_1 _4962_ (.A1(_1851_),
    .A2(net656),
    .Y(_0291_),
    .B1(_1850_));
 sg13g2_dfrbp_1 _4963_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net45),
    .D(_0036_),
    .Q_N(_2479_),
    .Q(\core.w[4] ));
 sg13g2_dfrbp_1 _4964_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net196),
    .D(_0037_),
    .Q_N(_2478_),
    .Q(\core.w[5] ));
 sg13g2_dfrbp_1 _4965_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net194),
    .D(_0038_),
    .Q_N(_2477_),
    .Q(\core.w[6] ));
 sg13g2_dfrbp_1 _4966_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net192),
    .D(_0039_),
    .Q_N(_2476_),
    .Q(\core.w[7] ));
 sg13g2_dfrbp_1 _4967_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net190),
    .D(_0040_),
    .Q_N(_2475_),
    .Q(\core.w[8] ));
 sg13g2_dfrbp_1 _4968_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net188),
    .D(_0041_),
    .Q_N(_2474_),
    .Q(\core.w[9] ));
 sg13g2_dfrbp_1 _4969_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net186),
    .D(_0042_),
    .Q_N(_2473_),
    .Q(\core.w[10] ));
 sg13g2_dfrbp_1 _4970_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net184),
    .D(_0043_),
    .Q_N(_2472_),
    .Q(\core.w[11] ));
 sg13g2_dfrbp_1 _4971_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net182),
    .D(_0044_),
    .Q_N(_2471_),
    .Q(\core.w[12] ));
 sg13g2_dfrbp_1 _4972_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net180),
    .D(_0045_),
    .Q_N(_2470_),
    .Q(\core.w[13] ));
 sg13g2_dfrbp_1 _4973_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net178),
    .D(_0046_),
    .Q_N(_2469_),
    .Q(\core.w[14] ));
 sg13g2_dfrbp_1 _4974_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net176),
    .D(net822),
    .Q_N(_0035_),
    .Q(\core.w[15] ));
 sg13g2_dfrbp_1 _4975_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net174),
    .D(_0048_),
    .Q_N(_2468_),
    .Q(\core.load_prev ));
 sg13g2_dfrbp_1 _4976_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net173),
    .D(_0049_),
    .Q_N(_2467_),
    .Q(\core.byte_acc[0] ));
 sg13g2_dfrbp_1 _4977_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net171),
    .D(_0050_),
    .Q_N(_2466_),
    .Q(\core.byte_acc[1] ));
 sg13g2_dfrbp_1 _4978_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net169),
    .D(_0051_),
    .Q_N(_2465_),
    .Q(\core.byte_acc[2] ));
 sg13g2_dfrbp_1 _4979_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net167),
    .D(_0052_),
    .Q_N(_2464_),
    .Q(\core.byte_acc[3] ));
 sg13g2_dfrbp_1 _4980_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net165),
    .D(net604),
    .Q_N(_0021_),
    .Q(\core.drive[0] ));
 sg13g2_dfrbp_1 _4981_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net164),
    .D(_0054_),
    .Q_N(_0024_),
    .Q(\core.drive[1] ));
 sg13g2_dfrbp_1 _4982_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net163),
    .D(_0055_),
    .Q_N(_0023_),
    .Q(\core.drive[2] ));
 sg13g2_dfrbp_1 _4983_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net162),
    .D(_0056_),
    .Q_N(_2463_),
    .Q(\core.drive[3] ));
 sg13g2_dfrbp_1 _4984_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net161),
    .D(net441),
    .Q_N(_2462_),
    .Q(\core.w8_reg[2] ));
 sg13g2_dfrbp_1 _4985_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net160),
    .D(net486),
    .Q_N(_2461_),
    .Q(\core.w8_reg[3] ));
 sg13g2_dfrbp_1 _4986_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net159),
    .D(net412),
    .Q_N(_2460_),
    .Q(\core.w8_reg[7] ));
 sg13g2_dfrbp_1 _4987_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net158),
    .D(net422),
    .Q_N(_2459_),
    .Q(\core.vm8_reg[2] ));
 sg13g2_dfrbp_1 _4988_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net157),
    .D(net418),
    .Q_N(_2458_),
    .Q(\core.vm8_reg[3] ));
 sg13g2_dfrbp_1 _4989_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net156),
    .D(net383),
    .Q_N(_2457_),
    .Q(\core.vm8_reg[7] ));
 sg13g2_dfrbp_1 _4990_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net155),
    .D(_0063_),
    .Q_N(_2456_),
    .Q(\core.dw[0] ));
 sg13g2_dfrbp_1 _4991_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net153),
    .D(_0064_),
    .Q_N(_2455_),
    .Q(\core.dw[1] ));
 sg13g2_dfrbp_1 _4992_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net151),
    .D(_0065_),
    .Q_N(_2454_),
    .Q(\core.dw[2] ));
 sg13g2_dfrbp_1 _4993_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net149),
    .D(_0066_),
    .Q_N(_2453_),
    .Q(\core.dw[3] ));
 sg13g2_dfrbp_1 _4994_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net147),
    .D(_0067_),
    .Q_N(_2452_),
    .Q(\core.dw[4] ));
 sg13g2_dfrbp_1 _4995_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net145),
    .D(_0068_),
    .Q_N(_2451_),
    .Q(\core.dw[5] ));
 sg13g2_dfrbp_1 _4996_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net143),
    .D(_0069_),
    .Q_N(_2450_),
    .Q(\core.dw[6] ));
 sg13g2_dfrbp_1 _4997_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net141),
    .D(_0070_),
    .Q_N(_2449_),
    .Q(\core.dw[7] ));
 sg13g2_dfrbp_1 _4998_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net139),
    .D(_0071_),
    .Q_N(_2448_),
    .Q(\core.dw[8] ));
 sg13g2_dfrbp_1 _4999_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net137),
    .D(_0072_),
    .Q_N(_2447_),
    .Q(\core.dw[9] ));
 sg13g2_dfrbp_1 _5000_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net135),
    .D(_0073_),
    .Q_N(_2446_),
    .Q(\core.dw[10] ));
 sg13g2_dfrbp_1 _5001_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net133),
    .D(_0074_),
    .Q_N(_2445_),
    .Q(\core.dw[11] ));
 sg13g2_dfrbp_1 _5002_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net131),
    .D(_0075_),
    .Q_N(_2444_),
    .Q(\core.dw[12] ));
 sg13g2_dfrbp_1 _5003_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net129),
    .D(_0076_),
    .Q_N(_2443_),
    .Q(\core.dw[13] ));
 sg13g2_dfrbp_1 _5004_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net127),
    .D(_0077_),
    .Q_N(_2442_),
    .Q(\core.dw[14] ));
 sg13g2_dfrbp_1 _5005_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net125),
    .D(_0078_),
    .Q_N(_2441_),
    .Q(\core.dw[15] ));
 sg13g2_dfrbp_1 _5006_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net123),
    .D(_0079_),
    .Q_N(_2440_),
    .Q(\core.dV[0] ));
 sg13g2_dfrbp_1 _5007_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net121),
    .D(net476),
    .Q_N(_2439_),
    .Q(\core.dV[1] ));
 sg13g2_dfrbp_1 _5008_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net119),
    .D(_0081_),
    .Q_N(_2438_),
    .Q(\core.dV[2] ));
 sg13g2_dfrbp_1 _5009_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net117),
    .D(_0082_),
    .Q_N(_2437_),
    .Q(\core.dV[3] ));
 sg13g2_dfrbp_1 _5010_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net115),
    .D(_0083_),
    .Q_N(_2436_),
    .Q(\core.dV[4] ));
 sg13g2_dfrbp_1 _5011_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net113),
    .D(_0084_),
    .Q_N(_2435_),
    .Q(\core.dV[5] ));
 sg13g2_dfrbp_1 _5012_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net111),
    .D(_0085_),
    .Q_N(_2434_),
    .Q(\core.dV[6] ));
 sg13g2_dfrbp_1 _5013_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net109),
    .D(_0086_),
    .Q_N(_2433_),
    .Q(\core.dV[7] ));
 sg13g2_dfrbp_1 _5014_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net107),
    .D(_0087_),
    .Q_N(_2432_),
    .Q(\core.dV[8] ));
 sg13g2_dfrbp_1 _5015_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net105),
    .D(_0088_),
    .Q_N(_2431_),
    .Q(\core.dV[9] ));
 sg13g2_dfrbp_1 _5016_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net103),
    .D(_0089_),
    .Q_N(_2430_),
    .Q(\core.dV[10] ));
 sg13g2_dfrbp_1 _5017_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net101),
    .D(_0090_),
    .Q_N(_2429_),
    .Q(\core.dV[11] ));
 sg13g2_dfrbp_1 _5018_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net99),
    .D(_0091_),
    .Q_N(_2428_),
    .Q(\core.dV[12] ));
 sg13g2_dfrbp_1 _5019_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net97),
    .D(_0092_),
    .Q_N(_2427_),
    .Q(\core.dV[13] ));
 sg13g2_dfrbp_1 _5020_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net95),
    .D(_0093_),
    .Q_N(_2426_),
    .Q(\core.dV[14] ));
 sg13g2_dfrbp_1 _5021_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net93),
    .D(_0094_),
    .Q_N(_2425_),
    .Q(\core.dV[15] ));
 sg13g2_dfrbp_1 _5022_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net91),
    .D(net819),
    .Q_N(_2424_),
    .Q(\core.leak[1] ));
 sg13g2_dfrbp_1 _5023_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net90),
    .D(net500),
    .Q_N(_2423_),
    .Q(\core.leak[2] ));
 sg13g2_dfrbp_1 _5024_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net89),
    .D(_0097_),
    .Q_N(_2422_),
    .Q(\core.leak[10] ));
 sg13g2_dfrbp_1 _5025_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net88),
    .D(net430),
    .Q_N(_0026_),
    .Q(\core.C_q[4] ));
 sg13g2_dfrbp_1 _5026_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net86),
    .D(net410),
    .Q_N(_0027_),
    .Q(\core.C_q[5] ));
 sg13g2_dfrbp_1 _5027_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net84),
    .D(net424),
    .Q_N(_0028_),
    .Q(\core.C_q[6] ));
 sg13g2_dfrbp_1 _5028_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net82),
    .D(_0101_),
    .Q_N(_0022_),
    .Q(\core.C_q[7] ));
 sg13g2_dfrbp_1 _5029_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net80),
    .D(net457),
    .Q_N(_0029_),
    .Q(\core.C_q[8] ));
 sg13g2_dfrbp_1 _5030_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net78),
    .D(net446),
    .Q_N(_0030_),
    .Q(\core.C_q[9] ));
 sg13g2_dfrbp_1 _5031_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net76),
    .D(_0104_),
    .Q_N(_0031_),
    .Q(\core.C_q[10] ));
 sg13g2_dfrbp_1 _5032_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net74),
    .D(net827),
    .Q_N(_0025_),
    .Q(\core.C_q[11] ));
 sg13g2_dfrbp_1 _5033_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net72),
    .D(net405),
    .Q_N(_2421_),
    .Q(\core.VT_q[4] ));
 sg13g2_dfrbp_1 _5034_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net70),
    .D(net516),
    .Q_N(_2420_),
    .Q(\core.VT_q[5] ));
 sg13g2_dfrbp_1 _5035_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net68),
    .D(net495),
    .Q_N(_2419_),
    .Q(\core.VT_q[6] ));
 sg13g2_dfrbp_1 _5036_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net66),
    .D(net532),
    .Q_N(_2418_),
    .Q(\core.VT_q[7] ));
 sg13g2_dfrbp_1 _5037_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net64),
    .D(net385),
    .Q_N(_2417_),
    .Q(\core.VT_q[8] ));
 sg13g2_dfrbp_1 _5038_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net62),
    .D(net530),
    .Q_N(_2416_),
    .Q(\core.VT_q[9] ));
 sg13g2_dfrbp_1 _5039_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net60),
    .D(net483),
    .Q_N(_2415_),
    .Q(\core.VT_q[10] ));
 sg13g2_dfrbp_1 _5040_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net58),
    .D(net468),
    .Q_N(_2414_),
    .Q(\core.VT_q[11] ));
 sg13g2_dfrbp_1 _5041_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net56),
    .D(net493),
    .Q_N(_2413_),
    .Q(\core.Vreset_q[4] ));
 sg13g2_dfrbp_1 _5042_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net54),
    .D(net491),
    .Q_N(_2412_),
    .Q(\core.Vreset_q[5] ));
 sg13g2_dfrbp_1 _5043_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net52),
    .D(net528),
    .Q_N(_2411_),
    .Q(\core.Vreset_q[6] ));
 sg13g2_dfrbp_1 _5044_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net50),
    .D(net534),
    .Q_N(_2410_),
    .Q(\core.Vreset_q[7] ));
 sg13g2_dfrbp_1 _5045_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net48),
    .D(net474),
    .Q_N(_2409_),
    .Q(\core.Vreset_q[8] ));
 sg13g2_dfrbp_1 _5046_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net46),
    .D(net513),
    .Q_N(_2408_),
    .Q(\core.Vreset_q[9] ));
 sg13g2_dfrbp_1 _5047_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net44),
    .D(net538),
    .Q_N(_2407_),
    .Q(\core.Vreset_q[10] ));
 sg13g2_dfrbp_1 _5048_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net42),
    .D(net414),
    .Q_N(_0008_),
    .Q(\core.Vreset_q[11] ));
 sg13g2_dfrbp_1 _5049_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net40),
    .D(net389),
    .Q_N(_2406_),
    .Q(\core.b_q[4] ));
 sg13g2_dfrbp_1 _5050_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net38),
    .D(net488),
    .Q_N(_2405_),
    .Q(\core.b_q[5] ));
 sg13g2_dfrbp_1 _5051_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net36),
    .D(net502),
    .Q_N(_2404_),
    .Q(\core.b_q[6] ));
 sg13g2_dfrbp_1 _5052_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net34),
    .D(net598),
    .Q_N(_2403_),
    .Q(\core.b_q[7] ));
 sg13g2_dfrbp_1 _5053_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net32),
    .D(net471),
    .Q_N(_2402_),
    .Q(\core.b_q[8] ));
 sg13g2_dfrbp_1 _5054_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net30),
    .D(net574),
    .Q_N(_2401_),
    .Q(\core.b_q[9] ));
 sg13g2_dfrbp_1 _5055_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net28),
    .D(net433),
    .Q_N(_2400_),
    .Q(\core.b_q[10] ));
 sg13g2_dfrbp_1 _5056_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net26),
    .D(net443),
    .Q_N(_2399_),
    .Q(\core.b_q[11] ));
 sg13g2_dfrbp_1 _5057_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net280),
    .D(net395),
    .Q_N(_2398_),
    .Q(\core.a_q[4] ));
 sg13g2_dfrbp_1 _5058_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net278),
    .D(net844),
    .Q_N(_2397_),
    .Q(\core.a_q[5] ));
 sg13g2_dfrbp_1 _5059_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net276),
    .D(net466),
    .Q_N(_2396_),
    .Q(\core.a_q[6] ));
 sg13g2_dfrbp_1 _5060_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net274),
    .D(net509),
    .Q_N(_2395_),
    .Q(\core.a_q[7] ));
 sg13g2_dfrbp_1 _5061_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net272),
    .D(net829),
    .Q_N(_2394_),
    .Q(\core.a_q[8] ));
 sg13g2_dfrbp_1 _5062_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net270),
    .D(net838),
    .Q_N(_2393_),
    .Q(\core.a_q[9] ));
 sg13g2_dfrbp_1 _5063_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net268),
    .D(net589),
    .Q_N(_2392_),
    .Q(\core.a_q[10] ));
 sg13g2_dfrbp_1 _5064_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net266),
    .D(_0137_),
    .Q_N(_2391_),
    .Q(\core.a_q[11] ));
 sg13g2_dfrbp_1 _5065_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net264),
    .D(net585),
    .Q_N(_0001_),
    .Q(\core.TauW_q[4] ));
 sg13g2_dfrbp_1 _5066_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net262),
    .D(net370),
    .Q_N(_0002_),
    .Q(\core.TauW_q[5] ));
 sg13g2_dfrbp_1 _5067_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net260),
    .D(_0140_),
    .Q_N(_0003_),
    .Q(\core.TauW_q[6] ));
 sg13g2_dfrbp_1 _5068_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net258),
    .D(net437),
    .Q_N(_0004_),
    .Q(\core.TauW_q[7] ));
 sg13g2_dfrbp_1 _5069_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net256),
    .D(_0142_),
    .Q_N(_0005_),
    .Q(\core.TauW_q[8] ));
 sg13g2_dfrbp_1 _5070_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net254),
    .D(_0143_),
    .Q_N(_0006_),
    .Q(\core.TauW_q[9] ));
 sg13g2_dfrbp_1 _5071_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net252),
    .D(_0144_),
    .Q_N(_0007_),
    .Q(\core.TauW_q[10] ));
 sg13g2_dfrbp_1 _5072_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net250),
    .D(net612),
    .Q_N(_0000_),
    .Q(\core.TauW_q[11] ));
 sg13g2_dfrbp_1 _5073_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net248),
    .D(_0146_),
    .Q_N(_2390_),
    .Q(\core.spike_reg ));
 sg13g2_dfrbp_1 _5074_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net246),
    .D(_0147_),
    .Q_N(_2389_),
    .Q(\core.V[0] ));
 sg13g2_dfrbp_1 _5075_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net244),
    .D(_0148_),
    .Q_N(_2388_),
    .Q(\core.V[1] ));
 sg13g2_dfrbp_1 _5076_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net242),
    .D(_0149_),
    .Q_N(_2387_),
    .Q(\core.V[2] ));
 sg13g2_dfrbp_1 _5077_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net240),
    .D(_0150_),
    .Q_N(_2386_),
    .Q(\core.V[3] ));
 sg13g2_dfrbp_1 _5078_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net238),
    .D(_0151_),
    .Q_N(_2385_),
    .Q(\core.V[4] ));
 sg13g2_dfrbp_1 _5079_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net236),
    .D(_0152_),
    .Q_N(_2384_),
    .Q(\core.V[5] ));
 sg13g2_dfrbp_1 _5080_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net234),
    .D(net841),
    .Q_N(_2383_),
    .Q(\core.V[6] ));
 sg13g2_dfrbp_1 _5081_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net232),
    .D(_0154_),
    .Q_N(_2382_),
    .Q(\core.V[7] ));
 sg13g2_dfrbp_1 _5082_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net230),
    .D(net866),
    .Q_N(_2381_),
    .Q(\core.V[8] ));
 sg13g2_dfrbp_1 _5083_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net228),
    .D(_0156_),
    .Q_N(_2380_),
    .Q(\core.V[9] ));
 sg13g2_dfrbp_1 _5084_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net226),
    .D(_0157_),
    .Q_N(_2379_),
    .Q(\core.V[10] ));
 sg13g2_dfrbp_1 _5085_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net224),
    .D(_0158_),
    .Q_N(_2378_),
    .Q(\core.V[11] ));
 sg13g2_dfrbp_1 _5086_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net222),
    .D(_0159_),
    .Q_N(_2377_),
    .Q(\core.V[12] ));
 sg13g2_dfrbp_1 _5087_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net220),
    .D(net864),
    .Q_N(_2376_),
    .Q(\core.V[13] ));
 sg13g2_dfrbp_1 _5088_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net218),
    .D(net859),
    .Q_N(_2375_),
    .Q(\core.V[14] ));
 sg13g2_dfrbp_1 _5089_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net216),
    .D(net869),
    .Q_N(_0034_),
    .Q(\core.V[15] ));
 sg13g2_dfrbp_1 _5090_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net214),
    .D(_0163_),
    .Q_N(_2374_),
    .Q(\core.w[0] ));
 sg13g2_dfrbp_1 _5091_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net212),
    .D(_0164_),
    .Q_N(_2373_),
    .Q(\core.w[1] ));
 sg13g2_dfrbp_1 _5092_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net210),
    .D(_0165_),
    .Q_N(_2372_),
    .Q(\core.w[2] ));
 sg13g2_dfrbp_1 _5093_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net208),
    .D(_0166_),
    .Q_N(_2371_),
    .Q(\core.w[3] ));
 sg13g2_dfrbp_1 _5094_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net206),
    .D(net851),
    .Q_N(_0016_),
    .Q(\core.lstate[2] ));
 sg13g2_dfrbp_1 _5095_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net205),
    .D(net854),
    .Q_N(_0020_),
    .Q(\core.lstate[1] ));
 sg13g2_dfrbp_1 _5096_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net204),
    .D(net522),
    .Q_N(_0018_),
    .Q(\core.lstate[0] ));
 sg13g2_dfrbp_1 _5097_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net203),
    .D(_0170_),
    .Q_N(_2370_),
    .Q(\core.byte_acc[4] ));
 sg13g2_dfrbp_1 _5098_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net201),
    .D(_0171_),
    .Q_N(_2369_),
    .Q(\core.byte_acc[5] ));
 sg13g2_dfrbp_1 _5099_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net199),
    .D(_0172_),
    .Q_N(_2368_),
    .Q(\core.byte_acc[6] ));
 sg13g2_dfrbp_1 _5100_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net197),
    .D(_0173_),
    .Q_N(_2367_),
    .Q(\core.byte_acc[7] ));
 sg13g2_dfrbp_1 _5101_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net193),
    .D(_0174_),
    .Q_N(_2366_),
    .Q(\core.s_VT[0] ));
 sg13g2_dfrbp_1 _5102_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net189),
    .D(_0175_),
    .Q_N(_2365_),
    .Q(\core.s_VT[1] ));
 sg13g2_dfrbp_1 _5103_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net185),
    .D(_0176_),
    .Q_N(_2364_),
    .Q(\core.s_VT[2] ));
 sg13g2_dfrbp_1 _5104_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net181),
    .D(_0177_),
    .Q_N(_2363_),
    .Q(\core.s_VT[3] ));
 sg13g2_dfrbp_1 _5105_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net177),
    .D(_0178_),
    .Q_N(_2362_),
    .Q(\core.s_VT[4] ));
 sg13g2_dfrbp_1 _5106_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net172),
    .D(_0179_),
    .Q_N(_2361_),
    .Q(\core.s_VT[5] ));
 sg13g2_dfrbp_1 _5107_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net168),
    .D(_0180_),
    .Q_N(_2360_),
    .Q(\core.s_VT[6] ));
 sg13g2_dfrbp_1 _5108_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net154),
    .D(net550),
    .Q_N(_2359_),
    .Q(\core.s_VT[7] ));
 sg13g2_dfrbp_1 _5109_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net150),
    .D(_0182_),
    .Q_N(_2358_),
    .Q(\core.s_C[0] ));
 sg13g2_dfrbp_1 _5110_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net146),
    .D(_0183_),
    .Q_N(_2357_),
    .Q(\core.s_C[1] ));
 sg13g2_dfrbp_1 _5111_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net142),
    .D(_0184_),
    .Q_N(_2356_),
    .Q(\core.s_C[2] ));
 sg13g2_dfrbp_1 _5112_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net138),
    .D(net547),
    .Q_N(_2355_),
    .Q(\core.s_C[3] ));
 sg13g2_dfrbp_1 _5113_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net134),
    .D(_0186_),
    .Q_N(_2354_),
    .Q(\core.s_C[4] ));
 sg13g2_dfrbp_1 _5114_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net130),
    .D(_0187_),
    .Q_N(_2353_),
    .Q(\core.s_C[5] ));
 sg13g2_dfrbp_1 _5115_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net126),
    .D(_0188_),
    .Q_N(_2352_),
    .Q(\core.s_C[6] ));
 sg13g2_dfrbp_1 _5116_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net122),
    .D(_0189_),
    .Q_N(_2351_),
    .Q(\core.s_C[7] ));
 sg13g2_dfrbp_1 _5117_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net118),
    .D(net428),
    .Q_N(_2350_),
    .Q(\core.p_TauW[0] ));
 sg13g2_dfrbp_1 _5118_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net114),
    .D(_0191_),
    .Q_N(_2349_),
    .Q(\core.p_TauW[1] ));
 sg13g2_dfrbp_1 _5119_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net110),
    .D(net583),
    .Q_N(_2348_),
    .Q(\core.p_TauW[2] ));
 sg13g2_dfrbp_1 _5120_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net106),
    .D(net416),
    .Q_N(_2347_),
    .Q(\core.p_TauW[3] ));
 sg13g2_dfrbp_1 _5121_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net102),
    .D(net397),
    .Q_N(_2346_),
    .Q(\core.p_TauW[4] ));
 sg13g2_dfrbp_1 _5122_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net98),
    .D(_0195_),
    .Q_N(_2345_),
    .Q(\core.p_TauW[5] ));
 sg13g2_dfrbp_1 _5123_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net94),
    .D(net453),
    .Q_N(_2344_),
    .Q(\core.p_TauW[6] ));
 sg13g2_dfrbp_1 _5124_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net87),
    .D(net399),
    .Q_N(_2343_),
    .Q(\core.p_TauW[7] ));
 sg13g2_dfrbp_1 _5125_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net83),
    .D(net387),
    .Q_N(_2342_),
    .Q(\core.p_a[0] ));
 sg13g2_dfrbp_1 _5126_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net79),
    .D(net439),
    .Q_N(_2341_),
    .Q(\core.p_a[1] ));
 sg13g2_dfrbp_1 _5127_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net75),
    .D(net358),
    .Q_N(_2340_),
    .Q(\core.p_a[2] ));
 sg13g2_dfrbp_1 _5128_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net71),
    .D(net368),
    .Q_N(_2339_),
    .Q(\core.p_a[3] ));
 sg13g2_dfrbp_1 _5129_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net67),
    .D(net354),
    .Q_N(_2338_),
    .Q(\core.p_a[4] ));
 sg13g2_dfrbp_1 _5130_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net63),
    .D(net381),
    .Q_N(_2337_),
    .Q(\core.p_a[5] ));
 sg13g2_dfrbp_1 _5131_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net59),
    .D(net356),
    .Q_N(_2336_),
    .Q(\core.p_a[6] ));
 sg13g2_dfrbp_1 _5132_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net55),
    .D(_0205_),
    .Q_N(_2335_),
    .Q(\core.p_a[7] ));
 sg13g2_dfrbp_1 _5133_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net51),
    .D(_0206_),
    .Q_N(_2334_),
    .Q(\core.p_b[0] ));
 sg13g2_dfrbp_1 _5134_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net47),
    .D(net364),
    .Q_N(_2333_),
    .Q(\core.p_b[1] ));
 sg13g2_dfrbp_1 _5135_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net43),
    .D(net426),
    .Q_N(_2332_),
    .Q(\core.p_b[2] ));
 sg13g2_dfrbp_1 _5136_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net39),
    .D(net497),
    .Q_N(_2331_),
    .Q(\core.p_b[3] ));
 sg13g2_dfrbp_1 _5137_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net35),
    .D(net377),
    .Q_N(_2330_),
    .Q(\core.p_b[4] ));
 sg13g2_dfrbp_1 _5138_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net31),
    .D(_0211_),
    .Q_N(_2329_),
    .Q(\core.p_b[5] ));
 sg13g2_dfrbp_1 _5139_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net27),
    .D(net391),
    .Q_N(_2328_),
    .Q(\core.p_b[6] ));
 sg13g2_dfrbp_1 _5140_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net279),
    .D(net393),
    .Q_N(_2327_),
    .Q(\core.p_b[7] ));
 sg13g2_dfrbp_1 _5141_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net275),
    .D(net524),
    .Q_N(_2326_),
    .Q(\core.p_Vreset[0] ));
 sg13g2_dfrbp_1 _5142_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net271),
    .D(net379),
    .Q_N(_2325_),
    .Q(\core.p_Vreset[1] ));
 sg13g2_dfrbp_1 _5143_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net267),
    .D(_0216_),
    .Q_N(_2324_),
    .Q(\core.p_Vreset[2] ));
 sg13g2_dfrbp_1 _5144_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net263),
    .D(net580),
    .Q_N(_2323_),
    .Q(\core.p_Vreset[3] ));
 sg13g2_dfrbp_1 _5145_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net259),
    .D(net450),
    .Q_N(_2322_),
    .Q(\core.p_Vreset[4] ));
 sg13g2_dfrbp_1 _5146_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net255),
    .D(net372),
    .Q_N(_2321_),
    .Q(\core.p_Vreset[5] ));
 sg13g2_dfrbp_1 _5147_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net251),
    .D(net366),
    .Q_N(_2320_),
    .Q(\core.p_Vreset[6] ));
 sg13g2_dfrbp_1 _5148_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net247),
    .D(net520),
    .Q_N(_0033_),
    .Q(\core.p_Vreset[7] ));
 sg13g2_dfrbp_1 _5149_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net243),
    .D(_0222_),
    .Q_N(_2319_),
    .Q(\core.p_VT[0] ));
 sg13g2_dfrbp_1 _5150_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net239),
    .D(net602),
    .Q_N(_2318_),
    .Q(\core.p_VT[1] ));
 sg13g2_dfrbp_1 _5151_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net235),
    .D(net420),
    .Q_N(_2317_),
    .Q(\core.p_VT[2] ));
 sg13g2_dfrbp_1 _5152_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net231),
    .D(net360),
    .Q_N(_2316_),
    .Q(\core.p_VT[3] ));
 sg13g2_dfrbp_1 _5153_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net227),
    .D(net362),
    .Q_N(_2315_),
    .Q(\core.p_VT[4] ));
 sg13g2_dfrbp_1 _5154_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net223),
    .D(net350),
    .Q_N(_2314_),
    .Q(\core.p_VT[5] ));
 sg13g2_dfrbp_1 _5155_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net219),
    .D(net480),
    .Q_N(_2313_),
    .Q(\core.p_VT[6] ));
 sg13g2_dfrbp_1 _5156_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net215),
    .D(net544),
    .Q_N(_0032_),
    .Q(\core.p_VT[7] ));
 sg13g2_dfrbp_1 _5157_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net211),
    .D(_0230_),
    .Q_N(_2312_),
    .Q(\core.p_C[0] ));
 sg13g2_dfrbp_1 _5158_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net207),
    .D(_0231_),
    .Q_N(_2311_),
    .Q(\core.p_C[1] ));
 sg13g2_dfrbp_1 _5159_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net200),
    .D(_0232_),
    .Q_N(_2310_),
    .Q(\core.p_C[2] ));
 sg13g2_dfrbp_1 _5160_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net195),
    .D(_0233_),
    .Q_N(_2309_),
    .Q(\core.p_C[3] ));
 sg13g2_dfrbp_1 _5161_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net187),
    .D(_0234_),
    .Q_N(_2308_),
    .Q(\core.p_C[4] ));
 sg13g2_dfrbp_1 _5162_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net179),
    .D(_0235_),
    .Q_N(_2307_),
    .Q(\core.p_C[5] ));
 sg13g2_dfrbp_1 _5163_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net170),
    .D(net462),
    .Q_N(_2306_),
    .Q(\core.p_C[6] ));
 sg13g2_dfrbp_1 _5164_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net152),
    .D(net435),
    .Q_N(_2305_),
    .Q(\core.p_C[7] ));
 sg13g2_dfrbp_1 _5165_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net144),
    .D(_0238_),
    .Q_N(_2304_),
    .Q(\core.params_ready ));
 sg13g2_dfrbp_1 _5166_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net136),
    .D(net408),
    .Q_N(_0017_),
    .Q(\core.nibble_cnt ));
 sg13g2_dfrbp_1 _5167_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net132),
    .D(net348),
    .Q_N(_0015_),
    .Q(\core.param_idx[0] ));
 sg13g2_dfrbp_1 _5168_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net128),
    .D(_0241_),
    .Q_N(_2303_),
    .Q(\core.param_idx[1] ));
 sg13g2_dfrbp_1 _5169_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net124),
    .D(_0242_),
    .Q_N(_2302_),
    .Q(\core.param_idx[2] ));
 sg13g2_dfrbp_1 _5170_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net120),
    .D(net375),
    .Q_N(_2301_),
    .Q(\core.param_idx[3] ));
 sg13g2_dfrbp_1 _5171_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net116),
    .D(_0244_),
    .Q_N(_2300_),
    .Q(\core.watchdog_cnt[0] ));
 sg13g2_dfrbp_1 _5172_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net112),
    .D(_0245_),
    .Q_N(_2299_),
    .Q(\core.watchdog_cnt[1] ));
 sg13g2_dfrbp_1 _5173_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net108),
    .D(_0246_),
    .Q_N(_0009_),
    .Q(\core.watchdog_cnt[2] ));
 sg13g2_dfrbp_1 _5174_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net104),
    .D(_0247_),
    .Q_N(_2298_),
    .Q(\core.watchdog_cnt[3] ));
 sg13g2_dfrbp_1 _5175_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net100),
    .D(_0248_),
    .Q_N(_0010_),
    .Q(\core.watchdog_cnt[4] ));
 sg13g2_dfrbp_1 _5176_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net96),
    .D(net402),
    .Q_N(_2297_),
    .Q(\core.watchdog_cnt[5] ));
 sg13g2_dfrbp_1 _5177_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net92),
    .D(_0250_),
    .Q_N(_0011_),
    .Q(\core.watchdog_cnt[6] ));
 sg13g2_dfrbp_1 _5178_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net85),
    .D(_0251_),
    .Q_N(_0019_),
    .Q(\core.watchdog_cnt[7] ));
 sg13g2_dfrbp_1 _5179_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net81),
    .D(_0252_),
    .Q_N(_2296_),
    .Q(\core.watchdog_cnt[8] ));
 sg13g2_dfrbp_1 _5180_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net77),
    .D(_0253_),
    .Q_N(_2295_),
    .Q(\core.watchdog_cnt[9] ));
 sg13g2_dfrbp_1 _5181_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net73),
    .D(_0254_),
    .Q_N(_0012_),
    .Q(\core.watchdog_cnt[10] ));
 sg13g2_dfrbp_1 _5182_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net69),
    .D(_0255_),
    .Q_N(_2294_),
    .Q(\core.watchdog_cnt[11] ));
 sg13g2_dfrbp_1 _5183_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net65),
    .D(_0256_),
    .Q_N(_0013_),
    .Q(\core.watchdog_cnt[12] ));
 sg13g2_dfrbp_1 _5184_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net61),
    .D(_0257_),
    .Q_N(_2293_),
    .Q(\core.watchdog_cnt[13] ));
 sg13g2_dfrbp_1 _5185_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net57),
    .D(_0258_),
    .Q_N(_0014_),
    .Q(\core.watchdog_cnt[14] ));
 sg13g2_dfrbp_1 _5186_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net53),
    .D(_0259_),
    .Q_N(_2292_),
    .Q(\core.watchdog_cnt[15] ));
 sg13g2_dfrbp_1 _5187_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net49),
    .D(_0260_),
    .Q_N(_2291_),
    .Q(\core.s_TauW[0] ));
 sg13g2_dfrbp_1 _5188_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net41),
    .D(_0261_),
    .Q_N(_2290_),
    .Q(\core.s_TauW[1] ));
 sg13g2_dfrbp_1 _5189_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net33),
    .D(_0262_),
    .Q_N(_2289_),
    .Q(\core.s_TauW[2] ));
 sg13g2_dfrbp_1 _5190_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net281),
    .D(_0263_),
    .Q_N(_2288_),
    .Q(\core.s_TauW[3] ));
 sg13g2_dfrbp_1 _5191_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net273),
    .D(_0264_),
    .Q_N(_2287_),
    .Q(\core.s_TauW[4] ));
 sg13g2_dfrbp_1 _5192_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net265),
    .D(_0265_),
    .Q_N(_2286_),
    .Q(\core.s_TauW[5] ));
 sg13g2_dfrbp_1 _5193_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net257),
    .D(_0266_),
    .Q_N(_2285_),
    .Q(\core.s_TauW[6] ));
 sg13g2_dfrbp_1 _5194_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net249),
    .D(_0267_),
    .Q_N(_2284_),
    .Q(\core.s_TauW[7] ));
 sg13g2_dfrbp_1 _5195_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net241),
    .D(_0268_),
    .Q_N(_2283_),
    .Q(\core.s_a[0] ));
 sg13g2_dfrbp_1 _5196_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net233),
    .D(_0269_),
    .Q_N(_2282_),
    .Q(\core.s_a[1] ));
 sg13g2_dfrbp_1 _5197_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net225),
    .D(_0270_),
    .Q_N(_2281_),
    .Q(\core.s_a[2] ));
 sg13g2_dfrbp_1 _5198_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net217),
    .D(_0271_),
    .Q_N(_2280_),
    .Q(\core.s_a[3] ));
 sg13g2_dfrbp_1 _5199_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net209),
    .D(_0272_),
    .Q_N(_2279_),
    .Q(\core.s_a[4] ));
 sg13g2_dfrbp_1 _5200_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net198),
    .D(_0273_),
    .Q_N(_2278_),
    .Q(\core.s_a[5] ));
 sg13g2_dfrbp_1 _5201_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net183),
    .D(_0274_),
    .Q_N(_2277_),
    .Q(\core.s_a[6] ));
 sg13g2_dfrbp_1 _5202_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net166),
    .D(_0275_),
    .Q_N(_2276_),
    .Q(\core.s_a[7] ));
 sg13g2_dfrbp_1 _5203_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net140),
    .D(_0276_),
    .Q_N(_2275_),
    .Q(\core.s_b[0] ));
 sg13g2_dfrbp_1 _5204_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net37),
    .D(_0277_),
    .Q_N(_2274_),
    .Q(\core.s_b[1] ));
 sg13g2_dfrbp_1 _5205_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net277),
    .D(_0278_),
    .Q_N(_2273_),
    .Q(\core.s_b[2] ));
 sg13g2_dfrbp_1 _5206_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net261),
    .D(_0279_),
    .Q_N(_2272_),
    .Q(\core.s_b[3] ));
 sg13g2_dfrbp_1 _5207_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net245),
    .D(_0280_),
    .Q_N(_2271_),
    .Q(\core.s_b[4] ));
 sg13g2_dfrbp_1 _5208_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net229),
    .D(_0281_),
    .Q_N(_2270_),
    .Q(\core.s_b[5] ));
 sg13g2_dfrbp_1 _5209_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net213),
    .D(_0282_),
    .Q_N(_2269_),
    .Q(\core.s_b[6] ));
 sg13g2_dfrbp_1 _5210_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net191),
    .D(_0283_),
    .Q_N(_2268_),
    .Q(\core.s_b[7] ));
 sg13g2_dfrbp_1 _5211_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net148),
    .D(_0284_),
    .Q_N(_2267_),
    .Q(\core.s_Vreset[0] ));
 sg13g2_dfrbp_1 _5212_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net29),
    .D(_0285_),
    .Q_N(_2266_),
    .Q(\core.s_Vreset[1] ));
 sg13g2_dfrbp_1 _5213_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net253),
    .D(_0286_),
    .Q_N(_2265_),
    .Q(\core.s_Vreset[2] ));
 sg13g2_dfrbp_1 _5214_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net221),
    .D(_0287_),
    .Q_N(_2264_),
    .Q(\core.s_Vreset[3] ));
 sg13g2_dfrbp_1 _5215_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net175),
    .D(_0288_),
    .Q_N(_2263_),
    .Q(\core.s_Vreset[4] ));
 sg13g2_dfrbp_1 _5216_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net269),
    .D(_0289_),
    .Q_N(_2262_),
    .Q(\core.s_Vreset[5] ));
 sg13g2_dfrbp_1 _5217_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net202),
    .D(_0290_),
    .Q_N(_2261_),
    .Q(\core.s_Vreset[6] ));
 sg13g2_dfrbp_1 _5218_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net237),
    .D(_0291_),
    .Q_N(_2260_),
    .Q(\core.s_Vreset[7] ));
 sg13g2_tiehi _5139__27 (.L_HI(net27));
 sg13g2_tiehi _5055__28 (.L_HI(net28));
 sg13g2_tiehi _5212__29 (.L_HI(net29));
 sg13g2_tiehi _5054__30 (.L_HI(net30));
 sg13g2_tiehi _5138__31 (.L_HI(net31));
 sg13g2_tiehi _5053__32 (.L_HI(net32));
 sg13g2_tiehi _5189__33 (.L_HI(net33));
 sg13g2_tiehi _5052__34 (.L_HI(net34));
 sg13g2_tiehi _5137__35 (.L_HI(net35));
 sg13g2_tiehi _5051__36 (.L_HI(net36));
 sg13g2_tiehi _5204__37 (.L_HI(net37));
 sg13g2_tiehi _5050__38 (.L_HI(net38));
 sg13g2_tiehi _5136__39 (.L_HI(net39));
 sg13g2_tiehi _5049__40 (.L_HI(net40));
 sg13g2_tiehi _5188__41 (.L_HI(net41));
 sg13g2_tiehi _5048__42 (.L_HI(net42));
 sg13g2_tiehi _5135__43 (.L_HI(net43));
 sg13g2_tiehi _5047__44 (.L_HI(net44));
 sg13g2_tiehi _4963__45 (.L_HI(net45));
 sg13g2_tiehi _5046__46 (.L_HI(net46));
 sg13g2_tiehi _5134__47 (.L_HI(net47));
 sg13g2_tiehi _5045__48 (.L_HI(net48));
 sg13g2_tiehi _5187__49 (.L_HI(net49));
 sg13g2_tiehi _5044__50 (.L_HI(net50));
 sg13g2_tiehi _5133__51 (.L_HI(net51));
 sg13g2_tiehi _5043__52 (.L_HI(net52));
 sg13g2_tiehi _5186__53 (.L_HI(net53));
 sg13g2_tiehi _5042__54 (.L_HI(net54));
 sg13g2_tiehi _5132__55 (.L_HI(net55));
 sg13g2_tiehi _5041__56 (.L_HI(net56));
 sg13g2_tiehi _5185__57 (.L_HI(net57));
 sg13g2_tiehi _5040__58 (.L_HI(net58));
 sg13g2_tiehi _5131__59 (.L_HI(net59));
 sg13g2_tiehi _5039__60 (.L_HI(net60));
 sg13g2_tiehi _5184__61 (.L_HI(net61));
 sg13g2_tiehi _5038__62 (.L_HI(net62));
 sg13g2_tiehi _5130__63 (.L_HI(net63));
 sg13g2_tiehi _5037__64 (.L_HI(net64));
 sg13g2_tiehi _5183__65 (.L_HI(net65));
 sg13g2_tiehi _5036__66 (.L_HI(net66));
 sg13g2_tiehi _5129__67 (.L_HI(net67));
 sg13g2_tiehi _5035__68 (.L_HI(net68));
 sg13g2_tiehi _5182__69 (.L_HI(net69));
 sg13g2_tiehi _5034__70 (.L_HI(net70));
 sg13g2_tiehi _5128__71 (.L_HI(net71));
 sg13g2_tiehi _5033__72 (.L_HI(net72));
 sg13g2_tiehi _5181__73 (.L_HI(net73));
 sg13g2_tiehi _5032__74 (.L_HI(net74));
 sg13g2_tiehi _5127__75 (.L_HI(net75));
 sg13g2_tiehi _5031__76 (.L_HI(net76));
 sg13g2_tiehi _5180__77 (.L_HI(net77));
 sg13g2_tiehi _5030__78 (.L_HI(net78));
 sg13g2_tiehi _5126__79 (.L_HI(net79));
 sg13g2_tiehi _5029__80 (.L_HI(net80));
 sg13g2_tiehi _5179__81 (.L_HI(net81));
 sg13g2_tiehi _5028__82 (.L_HI(net82));
 sg13g2_tiehi _5125__83 (.L_HI(net83));
 sg13g2_tiehi _5027__84 (.L_HI(net84));
 sg13g2_tiehi _5178__85 (.L_HI(net85));
 sg13g2_tiehi _5026__86 (.L_HI(net86));
 sg13g2_tiehi _5124__87 (.L_HI(net87));
 sg13g2_tiehi _5025__88 (.L_HI(net88));
 sg13g2_tiehi _5024__89 (.L_HI(net89));
 sg13g2_tiehi _5023__90 (.L_HI(net90));
 sg13g2_tiehi _5022__91 (.L_HI(net91));
 sg13g2_tiehi _5177__92 (.L_HI(net92));
 sg13g2_tiehi _5021__93 (.L_HI(net93));
 sg13g2_tiehi _5123__94 (.L_HI(net94));
 sg13g2_tiehi _5020__95 (.L_HI(net95));
 sg13g2_tiehi _5176__96 (.L_HI(net96));
 sg13g2_tiehi _5019__97 (.L_HI(net97));
 sg13g2_tiehi _5122__98 (.L_HI(net98));
 sg13g2_tiehi _5018__99 (.L_HI(net99));
 sg13g2_tiehi _5175__100 (.L_HI(net100));
 sg13g2_tiehi _5017__101 (.L_HI(net101));
 sg13g2_tiehi _5121__102 (.L_HI(net102));
 sg13g2_tiehi _5016__103 (.L_HI(net103));
 sg13g2_tiehi _5174__104 (.L_HI(net104));
 sg13g2_tiehi _5015__105 (.L_HI(net105));
 sg13g2_tiehi _5120__106 (.L_HI(net106));
 sg13g2_tiehi _5014__107 (.L_HI(net107));
 sg13g2_tiehi _5173__108 (.L_HI(net108));
 sg13g2_tiehi _5013__109 (.L_HI(net109));
 sg13g2_tiehi _5119__110 (.L_HI(net110));
 sg13g2_tiehi _5012__111 (.L_HI(net111));
 sg13g2_tiehi _5172__112 (.L_HI(net112));
 sg13g2_tiehi _5011__113 (.L_HI(net113));
 sg13g2_tiehi _5118__114 (.L_HI(net114));
 sg13g2_tiehi _5010__115 (.L_HI(net115));
 sg13g2_tiehi _5171__116 (.L_HI(net116));
 sg13g2_tiehi _5009__117 (.L_HI(net117));
 sg13g2_tiehi _5117__118 (.L_HI(net118));
 sg13g2_tiehi _5008__119 (.L_HI(net119));
 sg13g2_tiehi _5170__120 (.L_HI(net120));
 sg13g2_tiehi _5007__121 (.L_HI(net121));
 sg13g2_tiehi _5116__122 (.L_HI(net122));
 sg13g2_tiehi _5006__123 (.L_HI(net123));
 sg13g2_tiehi _5169__124 (.L_HI(net124));
 sg13g2_tiehi _5005__125 (.L_HI(net125));
 sg13g2_tiehi _5115__126 (.L_HI(net126));
 sg13g2_tiehi _5004__127 (.L_HI(net127));
 sg13g2_tiehi _5168__128 (.L_HI(net128));
 sg13g2_tiehi _5003__129 (.L_HI(net129));
 sg13g2_tiehi _5114__130 (.L_HI(net130));
 sg13g2_tiehi _5002__131 (.L_HI(net131));
 sg13g2_tiehi _5167__132 (.L_HI(net132));
 sg13g2_tiehi _5001__133 (.L_HI(net133));
 sg13g2_tiehi _5113__134 (.L_HI(net134));
 sg13g2_tiehi _5000__135 (.L_HI(net135));
 sg13g2_tiehi _5166__136 (.L_HI(net136));
 sg13g2_tiehi _4999__137 (.L_HI(net137));
 sg13g2_tiehi _5112__138 (.L_HI(net138));
 sg13g2_tiehi _4998__139 (.L_HI(net139));
 sg13g2_tiehi _5203__140 (.L_HI(net140));
 sg13g2_tiehi _4997__141 (.L_HI(net141));
 sg13g2_tiehi _5111__142 (.L_HI(net142));
 sg13g2_tiehi _4996__143 (.L_HI(net143));
 sg13g2_tiehi _5165__144 (.L_HI(net144));
 sg13g2_tiehi _4995__145 (.L_HI(net145));
 sg13g2_tiehi _5110__146 (.L_HI(net146));
 sg13g2_tiehi _4994__147 (.L_HI(net147));
 sg13g2_tiehi _5211__148 (.L_HI(net148));
 sg13g2_tiehi _4993__149 (.L_HI(net149));
 sg13g2_tiehi _5109__150 (.L_HI(net150));
 sg13g2_tiehi _4992__151 (.L_HI(net151));
 sg13g2_tiehi _5164__152 (.L_HI(net152));
 sg13g2_tiehi _4991__153 (.L_HI(net153));
 sg13g2_tiehi _5108__154 (.L_HI(net154));
 sg13g2_tiehi _4990__155 (.L_HI(net155));
 sg13g2_tiehi _4989__156 (.L_HI(net156));
 sg13g2_tiehi _4988__157 (.L_HI(net157));
 sg13g2_tiehi _4987__158 (.L_HI(net158));
 sg13g2_tiehi _4986__159 (.L_HI(net159));
 sg13g2_tiehi _4985__160 (.L_HI(net160));
 sg13g2_tiehi _4984__161 (.L_HI(net161));
 sg13g2_tiehi _4983__162 (.L_HI(net162));
 sg13g2_tiehi _4982__163 (.L_HI(net163));
 sg13g2_tiehi _4981__164 (.L_HI(net164));
 sg13g2_tiehi _4980__165 (.L_HI(net165));
 sg13g2_tiehi _5202__166 (.L_HI(net166));
 sg13g2_tiehi _4979__167 (.L_HI(net167));
 sg13g2_tiehi _5107__168 (.L_HI(net168));
 sg13g2_tiehi _4978__169 (.L_HI(net169));
 sg13g2_tiehi _5163__170 (.L_HI(net170));
 sg13g2_tiehi _4977__171 (.L_HI(net171));
 sg13g2_tiehi _5106__172 (.L_HI(net172));
 sg13g2_tiehi _4976__173 (.L_HI(net173));
 sg13g2_tiehi _4975__174 (.L_HI(net174));
 sg13g2_tiehi _5215__175 (.L_HI(net175));
 sg13g2_tiehi _4974__176 (.L_HI(net176));
 sg13g2_tiehi _5105__177 (.L_HI(net177));
 sg13g2_tiehi _4973__178 (.L_HI(net178));
 sg13g2_tiehi _5162__179 (.L_HI(net179));
 sg13g2_tiehi _4972__180 (.L_HI(net180));
 sg13g2_tiehi _5104__181 (.L_HI(net181));
 sg13g2_tiehi _4971__182 (.L_HI(net182));
 sg13g2_tiehi _5201__183 (.L_HI(net183));
 sg13g2_tiehi _4970__184 (.L_HI(net184));
 sg13g2_tiehi _5103__185 (.L_HI(net185));
 sg13g2_tiehi _4969__186 (.L_HI(net186));
 sg13g2_tiehi _5161__187 (.L_HI(net187));
 sg13g2_tiehi _4968__188 (.L_HI(net188));
 sg13g2_tiehi _5102__189 (.L_HI(net189));
 sg13g2_tiehi _4967__190 (.L_HI(net190));
 sg13g2_tiehi _5210__191 (.L_HI(net191));
 sg13g2_tiehi _4966__192 (.L_HI(net192));
 sg13g2_tiehi _5101__193 (.L_HI(net193));
 sg13g2_tiehi _4965__194 (.L_HI(net194));
 sg13g2_tiehi _5160__195 (.L_HI(net195));
 sg13g2_tiehi _4964__196 (.L_HI(net196));
 sg13g2_tiehi _5100__197 (.L_HI(net197));
 sg13g2_tiehi _5200__198 (.L_HI(net198));
 sg13g2_tiehi _5099__199 (.L_HI(net199));
 sg13g2_tiehi _5159__200 (.L_HI(net200));
 sg13g2_tiehi _5098__201 (.L_HI(net201));
 sg13g2_tiehi _5217__202 (.L_HI(net202));
 sg13g2_tiehi _5097__203 (.L_HI(net203));
 sg13g2_tiehi _5096__204 (.L_HI(net204));
 sg13g2_tiehi _5095__205 (.L_HI(net205));
 sg13g2_tiehi _5094__206 (.L_HI(net206));
 sg13g2_tiehi _5158__207 (.L_HI(net207));
 sg13g2_tiehi _5093__208 (.L_HI(net208));
 sg13g2_tiehi _5199__209 (.L_HI(net209));
 sg13g2_tiehi _5092__210 (.L_HI(net210));
 sg13g2_tiehi _5157__211 (.L_HI(net211));
 sg13g2_tiehi _5091__212 (.L_HI(net212));
 sg13g2_tiehi _5209__213 (.L_HI(net213));
 sg13g2_tiehi _5090__214 (.L_HI(net214));
 sg13g2_tiehi _5156__215 (.L_HI(net215));
 sg13g2_tiehi _5089__216 (.L_HI(net216));
 sg13g2_tiehi _5198__217 (.L_HI(net217));
 sg13g2_tiehi _5088__218 (.L_HI(net218));
 sg13g2_tiehi _5155__219 (.L_HI(net219));
 sg13g2_tiehi _5087__220 (.L_HI(net220));
 sg13g2_tiehi _5214__221 (.L_HI(net221));
 sg13g2_tiehi _5086__222 (.L_HI(net222));
 sg13g2_tiehi _5154__223 (.L_HI(net223));
 sg13g2_tiehi _5085__224 (.L_HI(net224));
 sg13g2_tiehi _5197__225 (.L_HI(net225));
 sg13g2_tiehi _5084__226 (.L_HI(net226));
 sg13g2_tiehi _5153__227 (.L_HI(net227));
 sg13g2_tiehi _5083__228 (.L_HI(net228));
 sg13g2_tiehi _5208__229 (.L_HI(net229));
 sg13g2_tiehi _5082__230 (.L_HI(net230));
 sg13g2_tiehi _5152__231 (.L_HI(net231));
 sg13g2_tiehi _5081__232 (.L_HI(net232));
 sg13g2_tiehi _5196__233 (.L_HI(net233));
 sg13g2_tiehi _5080__234 (.L_HI(net234));
 sg13g2_tiehi _5151__235 (.L_HI(net235));
 sg13g2_tiehi _5079__236 (.L_HI(net236));
 sg13g2_tiehi _5218__237 (.L_HI(net237));
 sg13g2_tiehi _5078__238 (.L_HI(net238));
 sg13g2_tiehi _5150__239 (.L_HI(net239));
 sg13g2_tiehi _5077__240 (.L_HI(net240));
 sg13g2_tiehi _5195__241 (.L_HI(net241));
 sg13g2_tiehi _5076__242 (.L_HI(net242));
 sg13g2_tiehi _5149__243 (.L_HI(net243));
 sg13g2_tiehi _5075__244 (.L_HI(net244));
 sg13g2_tiehi _5207__245 (.L_HI(net245));
 sg13g2_tiehi _5074__246 (.L_HI(net246));
 sg13g2_tiehi _5148__247 (.L_HI(net247));
 sg13g2_tiehi _5073__248 (.L_HI(net248));
 sg13g2_tiehi _5194__249 (.L_HI(net249));
 sg13g2_tiehi _5072__250 (.L_HI(net250));
 sg13g2_tiehi _5147__251 (.L_HI(net251));
 sg13g2_tiehi _5071__252 (.L_HI(net252));
 sg13g2_tiehi _5213__253 (.L_HI(net253));
 sg13g2_tiehi _5070__254 (.L_HI(net254));
 sg13g2_tiehi _5146__255 (.L_HI(net255));
 sg13g2_tiehi _5069__256 (.L_HI(net256));
 sg13g2_tiehi _5193__257 (.L_HI(net257));
 sg13g2_tiehi _5068__258 (.L_HI(net258));
 sg13g2_tiehi _5145__259 (.L_HI(net259));
 sg13g2_tiehi _5067__260 (.L_HI(net260));
 sg13g2_tiehi _5206__261 (.L_HI(net261));
 sg13g2_tiehi _5066__262 (.L_HI(net262));
 sg13g2_tiehi _5144__263 (.L_HI(net263));
 sg13g2_tiehi _5065__264 (.L_HI(net264));
 sg13g2_tiehi _5192__265 (.L_HI(net265));
 sg13g2_tiehi _5064__266 (.L_HI(net266));
 sg13g2_tiehi _5143__267 (.L_HI(net267));
 sg13g2_tiehi _5063__268 (.L_HI(net268));
 sg13g2_tiehi _5216__269 (.L_HI(net269));
 sg13g2_tiehi _5062__270 (.L_HI(net270));
 sg13g2_tiehi _5142__271 (.L_HI(net271));
 sg13g2_tiehi _5061__272 (.L_HI(net272));
 sg13g2_tiehi _5191__273 (.L_HI(net273));
 sg13g2_tiehi _5060__274 (.L_HI(net274));
 sg13g2_tiehi _5141__275 (.L_HI(net275));
 sg13g2_tiehi _5059__276 (.L_HI(net276));
 sg13g2_tiehi _5205__277 (.L_HI(net277));
 sg13g2_tiehi _5058__278 (.L_HI(net278));
 sg13g2_tiehi _5140__279 (.L_HI(net279));
 sg13g2_tiehi _5057__280 (.L_HI(net280));
 sg13g2_tiehi _5190__281 (.L_HI(net281));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_dpi_adexp_10 (.L_LO(net10));
 sg13g2_tielo tt_um_dpi_adexp_11 (.L_LO(net11));
 sg13g2_tielo tt_um_dpi_adexp_12 (.L_LO(net12));
 sg13g2_tielo tt_um_dpi_adexp_13 (.L_LO(net13));
 sg13g2_tielo tt_um_dpi_adexp_14 (.L_LO(net14));
 sg13g2_tielo tt_um_dpi_adexp_15 (.L_LO(net15));
 sg13g2_tielo tt_um_dpi_adexp_16 (.L_LO(net16));
 sg13g2_tielo tt_um_dpi_adexp_17 (.L_LO(net17));
 sg13g2_tielo tt_um_dpi_adexp_18 (.L_LO(net18));
 sg13g2_tielo tt_um_dpi_adexp_19 (.L_LO(net19));
 sg13g2_tielo tt_um_dpi_adexp_20 (.L_LO(net20));
 sg13g2_tielo tt_um_dpi_adexp_21 (.L_LO(net21));
 sg13g2_tielo tt_um_dpi_adexp_22 (.L_LO(net22));
 sg13g2_tielo tt_um_dpi_adexp_23 (.L_LO(net23));
 sg13g2_tielo tt_um_dpi_adexp_24 (.L_LO(net24));
 sg13g2_tielo tt_um_dpi_adexp_25 (.L_LO(net25));
 sg13g2_tiehi _5056__26 (.L_HI(net26));
 sg13g2_buf_1 _5492_ (.A(\core.spike_reg ),
    .X(uo_out[0]));
 sg13g2_buf_2 _5493_ (.A(uo_out[5]),
    .X(uo_out[2]));
 sg13g2_buf_2 _5494_ (.A(uo_out[5]),
    .X(uo_out[3]));
 sg13g2_buf_2 _5495_ (.A(uo_out[5]),
    .X(uo_out[4]));
 sg13g2_buf_2 fanout613 (.A(_1327_),
    .X(net613));
 sg13g2_buf_16 fanout614 (.X(net614),
    .A(net615));
 sg13g2_buf_8 fanout615 (.A(_0841_),
    .X(net615));
 sg13g2_buf_2 fanout616 (.A(net617),
    .X(net616));
 sg13g2_buf_2 fanout617 (.A(_1276_),
    .X(net617));
 sg13g2_buf_8 fanout618 (.A(_0709_),
    .X(net618));
 sg13g2_buf_8 fanout619 (.A(_1224_),
    .X(net619));
 sg13g2_buf_2 fanout620 (.A(_0671_),
    .X(net620));
 sg13g2_buf_16 fanout621 (.X(net621),
    .A(net622));
 sg13g2_buf_8 fanout622 (.A(_0665_),
    .X(net622));
 sg13g2_buf_2 fanout623 (.A(net624),
    .X(net623));
 sg13g2_buf_8 fanout624 (.A(_1180_),
    .X(net624));
 sg13g2_buf_8 fanout625 (.A(_1144_),
    .X(net625));
 sg13g2_buf_8 fanout626 (.A(_0585_),
    .X(net626));
 sg13g2_buf_8 fanout627 (.A(_0495_),
    .X(net627));
 sg13g2_buf_8 fanout628 (.A(_0494_),
    .X(net628));
 sg13g2_buf_4 fanout629 (.X(net629),
    .A(net630));
 sg13g2_buf_2 fanout630 (.A(net631),
    .X(net630));
 sg13g2_buf_4 fanout631 (.X(net631),
    .A(_2014_));
 sg13g2_buf_2 fanout632 (.A(net633),
    .X(net632));
 sg13g2_buf_1 fanout633 (.A(_2013_),
    .X(net633));
 sg13g2_buf_2 fanout634 (.A(net636),
    .X(net634));
 sg13g2_buf_2 fanout635 (.A(net636),
    .X(net635));
 sg13g2_buf_2 fanout636 (.A(_2013_),
    .X(net636));
 sg13g2_buf_2 fanout637 (.A(net638),
    .X(net637));
 sg13g2_buf_2 fanout638 (.A(_1991_),
    .X(net638));
 sg13g2_buf_2 fanout639 (.A(_1765_),
    .X(net639));
 sg13g2_buf_2 fanout640 (.A(_1765_),
    .X(net640));
 sg13g2_buf_4 fanout641 (.X(net641),
    .A(_1630_));
 sg13g2_buf_2 fanout642 (.A(_1630_),
    .X(net642));
 sg13g2_buf_2 fanout643 (.A(_1382_),
    .X(net643));
 sg13g2_buf_2 fanout644 (.A(_1382_),
    .X(net644));
 sg13g2_buf_2 fanout645 (.A(net646),
    .X(net645));
 sg13g2_buf_4 fanout646 (.X(net646),
    .A(_0946_));
 sg13g2_buf_2 fanout647 (.A(net648),
    .X(net647));
 sg13g2_buf_2 fanout648 (.A(_1833_),
    .X(net648));
 sg13g2_buf_2 fanout649 (.A(net650),
    .X(net649));
 sg13g2_buf_2 fanout650 (.A(_1824_),
    .X(net650));
 sg13g2_buf_2 fanout651 (.A(net653),
    .X(net651));
 sg13g2_buf_1 fanout652 (.A(net653),
    .X(net652));
 sg13g2_buf_2 fanout653 (.A(_1815_),
    .X(net653));
 sg13g2_buf_2 fanout654 (.A(net655),
    .X(net654));
 sg13g2_buf_2 fanout655 (.A(_1669_),
    .X(net655));
 sg13g2_buf_2 fanout656 (.A(_1842_),
    .X(net656));
 sg13g2_buf_2 fanout657 (.A(_1842_),
    .X(net657));
 sg13g2_buf_2 fanout658 (.A(net659),
    .X(net658));
 sg13g2_buf_2 fanout659 (.A(_1644_),
    .X(net659));
 sg13g2_buf_2 fanout660 (.A(net661),
    .X(net660));
 sg13g2_buf_2 fanout661 (.A(net662),
    .X(net661));
 sg13g2_buf_2 fanout662 (.A(net663),
    .X(net662));
 sg13g2_buf_2 fanout663 (.A(net674),
    .X(net663));
 sg13g2_buf_2 fanout664 (.A(net667),
    .X(net664));
 sg13g2_buf_2 fanout665 (.A(net667),
    .X(net665));
 sg13g2_buf_1 fanout666 (.A(net667),
    .X(net666));
 sg13g2_buf_2 fanout667 (.A(net674),
    .X(net667));
 sg13g2_buf_2 fanout668 (.A(net670),
    .X(net668));
 sg13g2_buf_1 fanout669 (.A(net670),
    .X(net669));
 sg13g2_buf_2 fanout670 (.A(net674),
    .X(net670));
 sg13g2_buf_2 fanout671 (.A(net672),
    .X(net671));
 sg13g2_buf_2 fanout672 (.A(net673),
    .X(net672));
 sg13g2_buf_1 fanout673 (.A(net674),
    .X(net673));
 sg13g2_buf_2 fanout674 (.A(_1637_),
    .X(net674));
 sg13g2_buf_2 fanout675 (.A(net676),
    .X(net675));
 sg13g2_buf_4 fanout676 (.X(net676),
    .A(_1634_));
 sg13g2_buf_2 fanout677 (.A(_2166_),
    .X(net677));
 sg13g2_buf_1 fanout678 (.A(_2166_),
    .X(net678));
 sg13g2_buf_2 fanout679 (.A(net680),
    .X(net679));
 sg13g2_buf_2 fanout680 (.A(_2159_),
    .X(net680));
 sg13g2_buf_8 fanout681 (.A(_2139_),
    .X(net681));
 sg13g2_buf_4 fanout682 (.X(net682),
    .A(_1965_));
 sg13g2_buf_4 fanout683 (.X(net683),
    .A(_1931_));
 sg13g2_buf_4 fanout684 (.X(net684),
    .A(_1930_));
 sg13g2_buf_4 fanout685 (.X(net685),
    .A(_1929_));
 sg13g2_buf_1 fanout686 (.A(_1929_),
    .X(net686));
 sg13g2_buf_4 fanout687 (.X(net687),
    .A(_1928_));
 sg13g2_buf_2 fanout688 (.A(net689),
    .X(net688));
 sg13g2_buf_1 fanout689 (.A(net693),
    .X(net689));
 sg13g2_buf_2 fanout690 (.A(net691),
    .X(net690));
 sg13g2_buf_2 fanout691 (.A(net692),
    .X(net691));
 sg13g2_buf_2 fanout692 (.A(net693),
    .X(net692));
 sg13g2_buf_2 fanout693 (.A(\core.params_ready ),
    .X(net693));
 sg13g2_buf_2 fanout694 (.A(net695),
    .X(net694));
 sg13g2_buf_1 fanout695 (.A(net696),
    .X(net695));
 sg13g2_buf_2 fanout696 (.A(net698),
    .X(net696));
 sg13g2_buf_2 fanout697 (.A(net698),
    .X(net697));
 sg13g2_buf_1 fanout698 (.A(\core.params_ready ),
    .X(net698));
 sg13g2_buf_2 fanout699 (.A(net700),
    .X(net699));
 sg13g2_buf_1 fanout700 (.A(net706),
    .X(net700));
 sg13g2_buf_2 fanout701 (.A(net702),
    .X(net701));
 sg13g2_buf_2 fanout702 (.A(net706),
    .X(net702));
 sg13g2_buf_2 fanout703 (.A(net705),
    .X(net703));
 sg13g2_buf_1 fanout704 (.A(net705),
    .X(net704));
 sg13g2_buf_2 fanout705 (.A(net706),
    .X(net705));
 sg13g2_buf_2 fanout706 (.A(\core.params_ready ),
    .X(net706));
 sg13g2_buf_2 fanout707 (.A(\core.lstate[1] ),
    .X(net707));
 sg13g2_buf_4 fanout708 (.X(net708),
    .A(net830));
 sg13g2_buf_4 fanout709 (.X(net709),
    .A(\core.V[8] ));
 sg13g2_buf_4 fanout710 (.X(net710),
    .A(\core.V[7] ));
 sg13g2_buf_4 fanout711 (.X(net711),
    .A(\core.V[6] ));
 sg13g2_buf_1 fanout712 (.A(\core.V[6] ),
    .X(net712));
 sg13g2_buf_8 fanout713 (.A(net714),
    .X(net713));
 sg13g2_buf_8 fanout714 (.A(\core.V[5] ),
    .X(net714));
 sg13g2_buf_16 fanout715 (.X(net715),
    .A(net716));
 sg13g2_buf_16 fanout716 (.X(net716),
    .A(net717));
 sg13g2_buf_8 fanout717 (.A(\core.V[4] ),
    .X(net717));
 sg13g2_buf_8 fanout718 (.A(net719),
    .X(net718));
 sg13g2_buf_8 fanout719 (.A(\core.V[3] ),
    .X(net719));
 sg13g2_buf_8 fanout720 (.A(net721),
    .X(net720));
 sg13g2_buf_8 fanout721 (.A(net722),
    .X(net721));
 sg13g2_buf_8 fanout722 (.A(\core.V[2] ),
    .X(net722));
 sg13g2_buf_8 fanout723 (.A(net724),
    .X(net723));
 sg13g2_buf_8 fanout724 (.A(net725),
    .X(net724));
 sg13g2_buf_8 fanout725 (.A(\core.V[1] ),
    .X(net725));
 sg13g2_buf_4 fanout726 (.X(net726),
    .A(net728));
 sg13g2_buf_2 fanout727 (.A(net728),
    .X(net727));
 sg13g2_buf_2 fanout728 (.A(\core.V[0] ),
    .X(net728));
 sg13g2_buf_4 fanout729 (.X(net729),
    .A(net730));
 sg13g2_buf_4 fanout730 (.X(net730),
    .A(\core.TauW_q[8] ));
 sg13g2_buf_4 fanout731 (.X(net731),
    .A(\core.TauW_q[7] ));
 sg13g2_buf_4 fanout732 (.X(net732),
    .A(\core.TauW_q[6] ));
 sg13g2_buf_4 fanout733 (.X(net733),
    .A(_0002_));
 sg13g2_buf_2 fanout734 (.A(net735),
    .X(net734));
 sg13g2_buf_4 fanout735 (.X(net735),
    .A(_0001_));
 sg13g2_buf_4 fanout736 (.X(net736),
    .A(net737));
 sg13g2_buf_2 fanout737 (.A(\core.TauW_q[4] ),
    .X(net737));
 sg13g2_buf_4 fanout738 (.X(net738),
    .A(\core.a_q[10] ));
 sg13g2_buf_2 fanout739 (.A(\core.a_q[9] ),
    .X(net739));
 sg13g2_buf_8 fanout740 (.A(\core.a_q[8] ),
    .X(net740));
 sg13g2_buf_2 fanout741 (.A(\core.a_q[7] ),
    .X(net741));
 sg13g2_buf_16 fanout742 (.X(net742),
    .A(net743));
 sg13g2_buf_16 fanout743 (.X(net743),
    .A(net744));
 sg13g2_buf_8 fanout744 (.A(\core.a_q[6] ),
    .X(net744));
 sg13g2_buf_4 fanout745 (.X(net745),
    .A(net746));
 sg13g2_buf_16 fanout746 (.X(net746),
    .A(net747));
 sg13g2_buf_8 fanout747 (.A(\core.a_q[5] ),
    .X(net747));
 sg13g2_buf_4 fanout748 (.X(net748),
    .A(\core.a_q[4] ));
 sg13g2_buf_1 fanout749 (.A(\core.a_q[4] ),
    .X(net749));
 sg13g2_buf_4 fanout750 (.X(net750),
    .A(_0030_));
 sg13g2_buf_4 fanout751 (.X(net751),
    .A(_0029_));
 sg13g2_buf_4 fanout752 (.X(net752),
    .A(_0028_));
 sg13g2_buf_4 fanout753 (.X(net753),
    .A(_0027_));
 sg13g2_buf_1 fanout754 (.A(_0027_),
    .X(net754));
 sg13g2_buf_4 fanout755 (.X(net755),
    .A(\core.C_q[5] ));
 sg13g2_buf_2 fanout756 (.A(\core.C_q[5] ),
    .X(net756));
 sg13g2_buf_4 fanout757 (.X(net757),
    .A(_0026_));
 sg13g2_buf_4 fanout758 (.X(net758),
    .A(\core.C_q[4] ));
 sg13g2_buf_2 fanout759 (.A(\core.C_q[4] ),
    .X(net759));
 sg13g2_buf_16 fanout760 (.X(net760),
    .A(net761));
 sg13g2_buf_16 fanout761 (.X(net761),
    .A(net762));
 sg13g2_buf_8 fanout762 (.A(\core.drive[3] ),
    .X(net762));
 sg13g2_buf_2 fanout763 (.A(net882),
    .X(net763));
 sg13g2_buf_2 fanout764 (.A(net765),
    .X(net764));
 sg13g2_buf_2 fanout765 (.A(net766),
    .X(net765));
 sg13g2_buf_2 fanout766 (.A(net770),
    .X(net766));
 sg13g2_buf_2 fanout767 (.A(net770),
    .X(net767));
 sg13g2_buf_2 fanout768 (.A(net769),
    .X(net768));
 sg13g2_buf_2 fanout769 (.A(net770),
    .X(net769));
 sg13g2_buf_2 fanout770 (.A(_2140_),
    .X(net770));
 sg13g2_buf_4 fanout771 (.X(net771),
    .A(_1958_));
 sg13g2_buf_2 fanout772 (.A(net773),
    .X(net772));
 sg13g2_buf_4 fanout773 (.X(net773),
    .A(_1958_));
 sg13g2_buf_4 fanout774 (.X(net774),
    .A(net777));
 sg13g2_buf_4 fanout775 (.X(net775),
    .A(net776));
 sg13g2_buf_4 fanout776 (.X(net776),
    .A(net777));
 sg13g2_buf_2 fanout777 (.A(_1958_),
    .X(net777));
 sg13g2_buf_2 fanout778 (.A(net779),
    .X(net778));
 sg13g2_buf_2 fanout779 (.A(net780),
    .X(net779));
 sg13g2_buf_4 fanout780 (.X(net780),
    .A(_1921_));
 sg13g2_buf_2 fanout781 (.A(net782),
    .X(net781));
 sg13g2_buf_2 fanout782 (.A(_1921_),
    .X(net782));
 sg13g2_buf_4 fanout783 (.X(net783),
    .A(net2));
 sg13g2_buf_2 fanout784 (.A(net787),
    .X(net784));
 sg13g2_buf_1 fanout785 (.A(net787),
    .X(net785));
 sg13g2_buf_2 fanout786 (.A(net787),
    .X(net786));
 sg13g2_buf_2 fanout787 (.A(net794),
    .X(net787));
 sg13g2_buf_2 fanout788 (.A(net794),
    .X(net788));
 sg13g2_buf_2 fanout789 (.A(net794),
    .X(net789));
 sg13g2_buf_4 fanout790 (.X(net790),
    .A(net794));
 sg13g2_buf_2 fanout791 (.A(net792),
    .X(net791));
 sg13g2_buf_2 fanout792 (.A(net793),
    .X(net792));
 sg13g2_buf_4 fanout793 (.X(net793),
    .A(net794));
 sg13g2_buf_2 fanout794 (.A(net812),
    .X(net794));
 sg13g2_buf_2 fanout795 (.A(net799),
    .X(net795));
 sg13g2_buf_2 fanout796 (.A(net799),
    .X(net796));
 sg13g2_buf_2 fanout797 (.A(net799),
    .X(net797));
 sg13g2_buf_1 fanout798 (.A(net799),
    .X(net798));
 sg13g2_buf_1 fanout799 (.A(net800),
    .X(net799));
 sg13g2_buf_2 fanout800 (.A(net812),
    .X(net800));
 sg13g2_buf_2 fanout801 (.A(net803),
    .X(net801));
 sg13g2_buf_2 fanout802 (.A(net803),
    .X(net802));
 sg13g2_buf_2 fanout803 (.A(net804),
    .X(net803));
 sg13g2_buf_2 fanout804 (.A(net812),
    .X(net804));
 sg13g2_buf_4 fanout805 (.X(net805),
    .A(net811));
 sg13g2_buf_2 fanout806 (.A(net811),
    .X(net806));
 sg13g2_buf_2 fanout807 (.A(net808),
    .X(net807));
 sg13g2_buf_2 fanout808 (.A(net809),
    .X(net808));
 sg13g2_buf_2 fanout809 (.A(net810),
    .X(net809));
 sg13g2_buf_4 fanout810 (.X(net810),
    .A(net811));
 sg13g2_buf_2 fanout811 (.A(net812),
    .X(net811));
 sg13g2_buf_2 fanout812 (.A(rst_n),
    .X(net812));
 sg13g2_buf_2 input1 (.A(ui_in[1]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[2]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[3]),
    .X(net3));
 sg13g2_buf_4 input4 (.X(net4),
    .A(ui_in[4]));
 sg13g2_buf_2 input5 (.A(uio_in[0]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(uio_in[1]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(uio_in[2]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(uio_in[3]),
    .X(net8));
 sg13g2_tielo tt_um_dpi_adexp_9 (.L_LO(net9));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_3_0__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_3_1__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkload3 (.A(clknet_3_4__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_1 clkload5 (.A(clknet_3_6__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_leaf_6_clk));
 sg13g2_inv_4 clkload8 (.A(clknet_leaf_35_clk));
 sg13g2_inv_8 clkload9 (.A(clknet_leaf_29_clk));
 sg13g2_inv_2 clkload10 (.A(clknet_leaf_30_clk));
 sg13g2_inv_2 clkload11 (.A(clknet_leaf_27_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_leaf_14_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_leaf_10_clk));
 sg13g2_inv_2 clkload14 (.A(clknet_leaf_22_clk));
 sg13g2_inv_4 clkload15 (.A(clknet_leaf_25_clk));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_21_clk));
 sg13g2_inv_4 clkload17 (.A(clknet_leaf_23_clk));
 sg13g2_dlygate4sd1_1 rebuffer1 (.A(_0494_),
    .X(net282));
 sg13g2_buf_1 rebuffer2 (.A(net282),
    .X(net283));
 sg13g2_dlygate4sd1_1 rebuffer3 (.A(_0495_),
    .X(net284));
 sg13g2_dlygate4sd1_1 rebuffer4 (.A(_0529_),
    .X(net285));
 sg13g2_dlygate4sd1_1 rebuffer5 (.A(_0503_),
    .X(net286));
 sg13g2_dlygate4sd1_1 rebuffer6 (.A(net286),
    .X(net287));
 sg13g2_dlygate4sd1_1 rebuffer7 (.A(_2251_),
    .X(net288));
 sg13g2_buf_1 rebuffer8 (.A(_0297_),
    .X(net289));
 sg13g2_dlygate4sd1_1 rebuffer9 (.A(_0709_),
    .X(net290));
 sg13g2_dlygate4sd1_1 rebuffer10 (.A(_2249_),
    .X(net291));
 sg13g2_dlygate4sd1_1 rebuffer11 (.A(_0345_),
    .X(net292));
 sg13g2_buf_2 rebuffer12 (.A(_0366_),
    .X(net293));
 sg13g2_buf_1 rebuffer13 (.A(_2214_),
    .X(net294));
 sg13g2_dlygate4sd1_1 rebuffer14 (.A(_0343_),
    .X(net295));
 sg13g2_buf_1 rebuffer15 (.A(_2248_),
    .X(net296));
 sg13g2_dlygate4sd1_1 rebuffer16 (.A(_2232_),
    .X(net297));
 sg13g2_dlygate4sd1_1 rebuffer17 (.A(_2231_),
    .X(net298));
 sg13g2_dlygate4sd1_1 rebuffer18 (.A(_2204_),
    .X(net299));
 sg13g2_dlygate4sd1_1 rebuffer19 (.A(_0371_),
    .X(net300));
 sg13g2_dlygate4sd1_1 rebuffer20 (.A(_2234_),
    .X(net301));
 sg13g2_dlygate4sd1_1 rebuffer21 (.A(_0378_),
    .X(net302));
 sg13g2_dlygate4sd1_1 rebuffer22 (.A(net305),
    .X(net303));
 sg13g2_dlygate4sd1_1 rebuffer23 (.A(_0348_),
    .X(net304));
 sg13g2_dlygate4sd1_1 rebuffer24 (.A(_0342_),
    .X(net305));
 sg13g2_dlygate4sd1_1 rebuffer25 (.A(_2216_),
    .X(net306));
 sg13g2_dlygate4sd1_1 rebuffer26 (.A(_2258_),
    .X(net307));
 sg13g2_dlygate4sd1_1 rebuffer27 (.A(\core.V[7] ),
    .X(net308));
 sg13g2_dlygate4sd1_1 rebuffer28 (.A(\core.a_q[11] ),
    .X(net309));
 sg13g2_dlygate4sd1_1 rebuffer29 (.A(\core.a_q[11] ),
    .X(net310));
 sg13g2_dlygate4sd1_1 rebuffer30 (.A(\core.a_q[11] ),
    .X(net311));
 sg13g2_dlygate4sd1_1 rebuffer31 (.A(\core.a_q[11] ),
    .X(net312));
 sg13g2_dlygate4sd1_1 rebuffer32 (.A(net717),
    .X(net313));
 sg13g2_dlygate4sd1_1 rebuffer33 (.A(net714),
    .X(net314));
 sg13g2_dlygate4sd1_1 rebuffer34 (.A(net747),
    .X(net315));
 sg13g2_dlygate4sd1_1 rebuffer35 (.A(net315),
    .X(net316));
 sg13g2_buf_1 rebuffer36 (.A(_2198_),
    .X(net317));
 sg13g2_buf_1 rebuffer37 (.A(_2242_),
    .X(net318));
 sg13g2_dlygate4sd1_1 rebuffer38 (.A(net725),
    .X(net319));
 sg13g2_dlygate4sd1_1 rebuffer39 (.A(_2245_),
    .X(net320));
 sg13g2_dlygate4sd1_1 rebuffer40 (.A(_2220_),
    .X(net321));
 sg13g2_dlygate4sd1_1 rebuffer41 (.A(_2259_),
    .X(net322));
 sg13g2_dlygate4sd1_1 rebuffer42 (.A(_0332_),
    .X(net323));
 sg13g2_dlygate4sd1_1 rebuffer43 (.A(_2238_),
    .X(net324));
 sg13g2_dlygate4sd1_1 rebuffer44 (.A(net324),
    .X(net325));
 sg13g2_dlygate4sd1_1 rebuffer45 (.A(net719),
    .X(net326));
 sg13g2_dlygate4sd1_1 rebuffer46 (.A(net326),
    .X(net327));
 sg13g2_dlygate4sd1_1 rebuffer47 (.A(net326),
    .X(net328));
 sg13g2_dlygate4sd1_1 rebuffer48 (.A(net715),
    .X(net329));
 sg13g2_buf_1 rebuffer49 (.A(net742),
    .X(net330));
 sg13g2_dlygate4sd1_1 rebuffer50 (.A(net714),
    .X(net331));
 sg13g2_dlygate4sd1_1 rebuffer51 (.A(_1040_),
    .X(net332));
 sg13g2_dlygate4sd1_1 rebuffer52 (.A(_1039_),
    .X(net333));
 sg13g2_buf_2 rebuffer53 (.A(_1007_),
    .X(net334));
 sg13g2_dlygate4sd1_1 rebuffer54 (.A(_1011_),
    .X(net335));
 sg13g2_dlygate4sd1_1 rebuffer55 (.A(\core.C_q[7] ),
    .X(net336));
 sg13g2_dlygate4sd1_1 rebuffer56 (.A(\core.C_q[7] ),
    .X(net337));
 sg13g2_dlygate4sd1_1 rebuffer57 (.A(net337),
    .X(net338));
 sg13g2_buf_1 rebuffer58 (.A(net338),
    .X(net339));
 sg13g2_dlygate4sd1_1 rebuffer59 (.A(net338),
    .X(net340));
 sg13g2_dlygate4sd1_1 rebuffer60 (.A(\core.C_q[10] ),
    .X(net341));
 sg13g2_dlygate4sd1_1 rebuffer61 (.A(\core.C_q[10] ),
    .X(net342));
 sg13g2_dlygate4sd1_1 rebuffer62 (.A(\core.drive[0] ),
    .X(net343));
 sg13g2_dlygate4sd1_1 rebuffer63 (.A(net343),
    .X(net344));
 sg13g2_dlygate4sd1_1 rebuffer64 (.A(\core.drive[0] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0015_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold66 (.A(_1758_),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0240_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold68 (.A(\core.s_VT[5] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0227_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold70 (.A(\core.p_a[7] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold71 (.A(\core.s_a[7] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold72 (.A(\core.s_a[4] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0202_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold74 (.A(\core.s_a[6] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0204_),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold76 (.A(\core.s_a[2] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0200_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold78 (.A(\core.s_VT[3] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0225_),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold80 (.A(\core.s_VT[4] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0226_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold82 (.A(\core.s_b[1] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0207_),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold84 (.A(\core.s_Vreset[6] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0220_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold86 (.A(\core.s_a[3] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0201_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold88 (.A(\core.p_TauW[1] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0139_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold90 (.A(\core.s_Vreset[5] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0219_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold92 (.A(\core.s_TauW[1] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold93 (.A(\core.param_idx[3] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0243_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold95 (.A(\core.s_b[4] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0210_),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold97 (.A(\core.s_Vreset[1] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0215_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold99 (.A(\core.s_a[5] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0203_),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold101 (.A(\core.vm8_reg[7] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0062_),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold103 (.A(\core.p_VT[4] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0110_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold105 (.A(\core.s_a[0] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0198_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold107 (.A(\core.p_b[0] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0122_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold109 (.A(\core.s_b[6] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0212_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold111 (.A(\core.s_b[7] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0213_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold113 (.A(\core.p_a[0] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0130_),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold115 (.A(\core.s_TauW[4] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0194_),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold117 (.A(\core.s_TauW[7] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0197_),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold119 (.A(\core.watchdog_cnt[5] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold120 (.A(_1781_),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0249_),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold122 (.A(\core.s_b[0] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold123 (.A(\core.p_VT[0] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0106_),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold125 (.A(\core.nibble_cnt ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold126 (.A(_1750_),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0239_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold128 (.A(\core.p_C[1] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0099_),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold130 (.A(\core.w8_reg[7] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0059_),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0033_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0121_),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold134 (.A(\core.s_TauW[3] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0193_),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold136 (.A(\core.vm8_reg[3] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0061_),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold138 (.A(\core.s_VT[2] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0224_),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold140 (.A(\core.vm8_reg[2] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0060_),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold142 (.A(\core.p_C[2] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0100_),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold144 (.A(\core.s_b[2] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0208_),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold146 (.A(\core.s_TauW[0] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0190_),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold148 (.A(\core.p_C[0] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0098_),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold150 (.A(\core.leak[10] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold151 (.A(\core.p_b[6] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0128_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold153 (.A(\core.s_C[7] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0237_),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold155 (.A(\core.p_TauW[3] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0141_),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold157 (.A(\core.s_a[1] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0199_),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold159 (.A(\core.w8_reg[2] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0057_),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold161 (.A(\core.p_b[7] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0129_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold163 (.A(\core.dV[4] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold164 (.A(\core.p_C[5] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0103_),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold166 (.A(\core.dV[2] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold167 (.A(\core.s_C[0] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold168 (.A(\core.s_Vreset[4] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0218_),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold170 (.A(\core.s_C[2] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold171 (.A(\core.s_TauW[6] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0196_),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold173 (.A(\core.dV[7] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold174 (.A(\core.dV[3] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold175 (.A(\core.p_C[4] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0102_),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold177 (.A(\core.drive[2] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold178 (.A(\core.watchdog_cnt[15] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold179 (.A(_1813_),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold180 (.A(\core.s_C[6] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0236_),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold182 (.A(\core.p_TauW[4] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold183 (.A(\core.dV[6] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold184 (.A(\core.p_a[2] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0132_),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0032_),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0113_),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold188 (.A(\core.dw[11] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold189 (.A(\core.p_b[4] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0126_),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold191 (.A(\core.dw[0] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold192 (.A(\core.p_Vreset[4] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0118_),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold194 (.A(\core.dV[1] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0080_),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold196 (.A(\core.watchdog_cnt[9] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold197 (.A(_1792_),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold198 (.A(\core.s_VT[6] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0228_),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold200 (.A(\core.s_VT[0] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold201 (.A(\core.VT_q[10] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold202 (.A(_0112_),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold203 (.A(\core.s_C[4] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold204 (.A(\core.w8_reg[3] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0058_),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold206 (.A(\core.p_b[1] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0123_),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold208 (.A(\core.drive[1] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold209 (.A(\core.Vreset_q[5] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold210 (.A(_0115_),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold211 (.A(\core.Vreset_q[4] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0114_),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold213 (.A(\core.VT_q[6] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0108_),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold215 (.A(\core.s_b[3] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold216 (.A(_0209_),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold217 (.A(\core.dw[1] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold218 (.A(\core.leak[2] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0096_),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold220 (.A(\core.p_b[2] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold221 (.A(_0124_),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold222 (.A(\core.dV[9] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold223 (.A(\core.dV[10] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold224 (.A(\core.dw[4] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold225 (.A(_0014_),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold226 (.A(_1811_),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold227 (.A(\core.p_a[3] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold228 (.A(_0133_),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold229 (.A(\core.spike_reg ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold230 (.A(\core.dV[5] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold231 (.A(\core.Vreset_q[9] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold232 (.A(_0119_),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold233 (.A(\core.dw[10] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold234 (.A(\core.VT_q[5] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold235 (.A(_0107_),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold236 (.A(\core.watchdog_cnt[2] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold237 (.A(_1772_),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold238 (.A(\core.p_Vreset[7] ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold239 (.A(_0221_),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0018_),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold241 (.A(_0169_),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold242 (.A(\core.s_Vreset[0] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold243 (.A(_0214_),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold244 (.A(\core.watchdog_cnt[4] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold245 (.A(_1778_),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold246 (.A(\core.p_Vreset[2] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold247 (.A(_0116_),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold248 (.A(\core.p_VT[5] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold249 (.A(_0111_),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold250 (.A(\core.VT_q[7] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0109_),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold252 (.A(\core.Vreset_q[7] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold253 (.A(_0117_),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold254 (.A(\core.s_C[5] ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold255 (.A(\core.dV[8] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold256 (.A(\core.p_Vreset[6] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold257 (.A(_0120_),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold258 (.A(\core.dw[6] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold259 (.A(\core.watchdog_cnt[7] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold260 (.A(_1786_),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold261 (.A(\core.dw[2] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold262 (.A(\core.p_VT[7] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold263 (.A(_0229_),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold264 (.A(\core.byte_acc[4] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold265 (.A(\core.s_C[3] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold266 (.A(_0185_),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold267 (.A(\core.byte_acc[0] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold268 (.A(\core.s_VT[7] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold269 (.A(_0181_),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold270 (.A(\core.dV[15] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold271 (.A(\core.dV[11] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold272 (.A(\core.dw[15] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold273 (.A(\core.param_idx[2] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold274 (.A(\core.s_Vreset[2] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold275 (.A(\core.dw[7] ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold276 (.A(\core.byte_acc[6] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold277 (.A(\core.dV[12] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold278 (.A(\core.dw[3] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold279 (.A(\core.param_idx[0] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold280 (.A(\core.dV[13] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold281 (.A(\core.byte_acc[7] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold282 (.A(\core.param_idx[1] ),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold283 (.A(_1668_),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold284 (.A(_0013_),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold285 (.A(_1803_),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold286 (.A(_1804_),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold287 (.A(\core.byte_acc[1] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold288 (.A(\core.dV[0] ),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold289 (.A(\core.byte_acc[2] ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold290 (.A(_0012_),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold291 (.A(_1796_),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold292 (.A(\core.b_q[9] ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold293 (.A(_0127_),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold294 (.A(\core.byte_acc[3] ),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold295 (.A(\core.p_C[3] ),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold296 (.A(\core.byte_acc[5] ),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold297 (.A(\core.dw[14] ),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold298 (.A(\core.s_Vreset[3] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold299 (.A(_0217_),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold300 (.A(\core.dw[8] ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold301 (.A(\core.s_TauW[2] ),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold302 (.A(_0192_),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold303 (.A(\core.p_TauW[0] ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold304 (.A(_0138_),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold305 (.A(\core.watchdog_cnt[6] ),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold306 (.A(_1784_),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold307 (.A(\core.a_q[10] ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold308 (.A(_0136_),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold309 (.A(\core.s_Vreset[7] ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold310 (.A(\core.param_idx[3] ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold311 (.A(\core.param_idx[1] ),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold312 (.A(\core.dw[5] ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold313 (.A(\core.s_b[5] ),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold314 (.A(\core.watchdog_cnt[3] ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold315 (.A(_1776_),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold316 (.A(\core.b_q[7] ),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold317 (.A(_0125_),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold318 (.A(\core.s_C[1] ),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold319 (.A(\core.p_b[5] ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold320 (.A(\core.s_VT[1] ),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold321 (.A(_0223_),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold322 (.A(\core.drive[0] ),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold323 (.A(_0053_),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold324 (.A(\core.dw[9] ),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold325 (.A(\core.dV[14] ),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold326 (.A(\core.lstate[0] ),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold327 (.A(\core.watchdog_cnt[13] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold328 (.A(_1808_),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold329 (.A(\core.s_TauW[5] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold330 (.A(\core.p_TauW[7] ),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold331 (.A(_0145_),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold332 (.A(\core.p_TauW[5] ),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold333 (.A(\core.watchdog_cnt[11] ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold334 (.A(_1801_),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold335 (.A(\core.watchdog_cnt[8] ),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold336 (.A(\core.dw[12] ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold337 (.A(\core.leak[1] ),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold338 (.A(_0095_),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold339 (.A(\core.w[15] ),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold340 (.A(_1989_),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold341 (.A(_0047_),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold342 (.A(\core.dw[13] ),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold343 (.A(_1953_),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold344 (.A(\core.param_idx[0] ),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold345 (.A(\core.C_q[11] ),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold346 (.A(_0105_),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold347 (.A(\core.p_a[4] ),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold348 (.A(_0134_),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold349 (.A(\core.w[0] ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold350 (.A(\core.watchdog_cnt[1] ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold351 (.A(_1770_),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold352 (.A(\core.w[10] ),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold353 (.A(\core.w[4] ),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold354 (.A(\core.p_TauW[6] ),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold355 (.A(\core.w[11] ),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold356 (.A(\core.p_a[5] ),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold357 (.A(_0135_),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold358 (.A(\core.p_TauW[2] ),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold359 (.A(\core.Vreset_q[6] ),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold360 (.A(_0153_),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold361 (.A(\core.w[8] ),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold362 (.A(\core.p_a[1] ),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold363 (.A(_0131_),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold364 (.A(net710),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold365 (.A(\core.V[12] ),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold366 (.A(_1588_),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold367 (.A(net717),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold368 (.A(\core.w[5] ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold369 (.A(\core.lstate[2] ),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold370 (.A(_0167_),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold371 (.A(\core.watchdog_cnt[0] ),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold372 (.A(_0020_),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold373 (.A(_0168_),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold374 (.A(\core.p_C[6] ),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold375 (.A(net722),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold376 (.A(_1510_),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold377 (.A(\core.Vreset_q[11] ),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold378 (.A(_0161_),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold379 (.A(net762),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold380 (.A(\core.V[10] ),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold381 (.A(_1574_),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold382 (.A(\core.V[13] ),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold383 (.A(_0160_),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold384 (.A(\core.Vreset_q[8] ),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold385 (.A(_0155_),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold386 (.A(\core.w[1] ),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold387 (.A(_0034_),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold388 (.A(_0162_),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold389 (.A(\core.w[2] ),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold390 (.A(_1617_),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold391 (.A(\core.V[9] ),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold392 (.A(_1567_),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold393 (.A(net724),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold394 (.A(\core.V[11] ),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold395 (.A(_1581_),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold396 (.A(\core.w[6] ),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold397 (.A(\core.w[3] ),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold398 (.A(net714),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold399 (.A(\core.w[13] ),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold400 (.A(\core.w[7] ),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold401 (.A(\core.w[14] ),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold402 (.A(\core.w[12] ),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold403 (.A(\core.dV[2] ),
    .X(net884));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_4 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_71 ();
 sg13g2_decap_8 FILLER_0_82 ();
 sg13g2_decap_8 FILLER_0_89 ();
 sg13g2_decap_8 FILLER_0_96 ();
 sg13g2_decap_8 FILLER_0_103 ();
 sg13g2_decap_4 FILLER_0_110 ();
 sg13g2_fill_1 FILLER_0_114 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_fill_2 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_302 ();
 sg13g2_decap_8 FILLER_0_309 ();
 sg13g2_decap_8 FILLER_0_316 ();
 sg13g2_decap_8 FILLER_0_323 ();
 sg13g2_decap_8 FILLER_0_330 ();
 sg13g2_decap_8 FILLER_0_337 ();
 sg13g2_decap_8 FILLER_0_344 ();
 sg13g2_decap_8 FILLER_0_351 ();
 sg13g2_decap_8 FILLER_0_358 ();
 sg13g2_decap_8 FILLER_0_365 ();
 sg13g2_decap_8 FILLER_0_372 ();
 sg13g2_decap_8 FILLER_0_379 ();
 sg13g2_decap_8 FILLER_0_386 ();
 sg13g2_decap_8 FILLER_0_393 ();
 sg13g2_decap_8 FILLER_0_400 ();
 sg13g2_fill_2 FILLER_0_407 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_4 FILLER_1_56 ();
 sg13g2_fill_2 FILLER_1_60 ();
 sg13g2_fill_2 FILLER_1_68 ();
 sg13g2_fill_2 FILLER_1_75 ();
 sg13g2_fill_1 FILLER_1_77 ();
 sg13g2_fill_2 FILLER_1_99 ();
 sg13g2_fill_1 FILLER_1_101 ();
 sg13g2_fill_2 FILLER_1_118 ();
 sg13g2_fill_1 FILLER_1_120 ();
 sg13g2_decap_8 FILLER_1_130 ();
 sg13g2_decap_8 FILLER_1_137 ();
 sg13g2_decap_8 FILLER_1_144 ();
 sg13g2_decap_8 FILLER_1_151 ();
 sg13g2_decap_8 FILLER_1_158 ();
 sg13g2_decap_8 FILLER_1_165 ();
 sg13g2_decap_8 FILLER_1_172 ();
 sg13g2_decap_8 FILLER_1_179 ();
 sg13g2_decap_8 FILLER_1_186 ();
 sg13g2_decap_8 FILLER_1_193 ();
 sg13g2_decap_8 FILLER_1_200 ();
 sg13g2_decap_8 FILLER_1_207 ();
 sg13g2_decap_8 FILLER_1_214 ();
 sg13g2_decap_8 FILLER_1_221 ();
 sg13g2_decap_8 FILLER_1_228 ();
 sg13g2_decap_8 FILLER_1_235 ();
 sg13g2_decap_8 FILLER_1_242 ();
 sg13g2_decap_8 FILLER_1_249 ();
 sg13g2_decap_8 FILLER_1_256 ();
 sg13g2_decap_8 FILLER_1_316 ();
 sg13g2_decap_8 FILLER_1_323 ();
 sg13g2_decap_8 FILLER_1_330 ();
 sg13g2_decap_8 FILLER_1_337 ();
 sg13g2_decap_8 FILLER_1_344 ();
 sg13g2_decap_8 FILLER_1_351 ();
 sg13g2_decap_8 FILLER_1_358 ();
 sg13g2_decap_8 FILLER_1_365 ();
 sg13g2_decap_8 FILLER_1_372 ();
 sg13g2_decap_8 FILLER_1_379 ();
 sg13g2_decap_8 FILLER_1_386 ();
 sg13g2_decap_8 FILLER_1_393 ();
 sg13g2_decap_8 FILLER_1_400 ();
 sg13g2_fill_2 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_4 FILLER_2_49 ();
 sg13g2_fill_2 FILLER_2_53 ();
 sg13g2_fill_1 FILLER_2_71 ();
 sg13g2_fill_2 FILLER_2_96 ();
 sg13g2_fill_1 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_136 ();
 sg13g2_decap_8 FILLER_2_143 ();
 sg13g2_decap_8 FILLER_2_150 ();
 sg13g2_decap_8 FILLER_2_157 ();
 sg13g2_decap_8 FILLER_2_164 ();
 sg13g2_decap_8 FILLER_2_171 ();
 sg13g2_decap_8 FILLER_2_178 ();
 sg13g2_decap_8 FILLER_2_185 ();
 sg13g2_decap_8 FILLER_2_192 ();
 sg13g2_decap_8 FILLER_2_199 ();
 sg13g2_decap_8 FILLER_2_206 ();
 sg13g2_decap_8 FILLER_2_213 ();
 sg13g2_decap_8 FILLER_2_220 ();
 sg13g2_decap_8 FILLER_2_227 ();
 sg13g2_decap_8 FILLER_2_234 ();
 sg13g2_decap_8 FILLER_2_241 ();
 sg13g2_decap_4 FILLER_2_248 ();
 sg13g2_fill_2 FILLER_2_252 ();
 sg13g2_fill_1 FILLER_2_268 ();
 sg13g2_fill_1 FILLER_2_276 ();
 sg13g2_fill_2 FILLER_2_322 ();
 sg13g2_fill_1 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_334 ();
 sg13g2_decap_8 FILLER_2_341 ();
 sg13g2_decap_8 FILLER_2_348 ();
 sg13g2_decap_8 FILLER_2_355 ();
 sg13g2_decap_8 FILLER_2_362 ();
 sg13g2_decap_8 FILLER_2_369 ();
 sg13g2_decap_8 FILLER_2_376 ();
 sg13g2_decap_8 FILLER_2_383 ();
 sg13g2_decap_8 FILLER_2_390 ();
 sg13g2_decap_8 FILLER_2_397 ();
 sg13g2_decap_4 FILLER_2_404 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_fill_2 FILLER_3_49 ();
 sg13g2_fill_2 FILLER_3_86 ();
 sg13g2_fill_1 FILLER_3_88 ();
 sg13g2_fill_1 FILLER_3_98 ();
 sg13g2_decap_4 FILLER_3_111 ();
 sg13g2_decap_8 FILLER_3_144 ();
 sg13g2_decap_8 FILLER_3_151 ();
 sg13g2_decap_8 FILLER_3_158 ();
 sg13g2_decap_8 FILLER_3_165 ();
 sg13g2_decap_8 FILLER_3_172 ();
 sg13g2_decap_8 FILLER_3_179 ();
 sg13g2_decap_8 FILLER_3_186 ();
 sg13g2_decap_8 FILLER_3_193 ();
 sg13g2_decap_8 FILLER_3_200 ();
 sg13g2_decap_8 FILLER_3_207 ();
 sg13g2_decap_8 FILLER_3_214 ();
 sg13g2_decap_8 FILLER_3_221 ();
 sg13g2_decap_8 FILLER_3_228 ();
 sg13g2_decap_4 FILLER_3_235 ();
 sg13g2_fill_1 FILLER_3_326 ();
 sg13g2_fill_1 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_363 ();
 sg13g2_decap_8 FILLER_3_370 ();
 sg13g2_decap_8 FILLER_3_377 ();
 sg13g2_decap_8 FILLER_3_384 ();
 sg13g2_decap_8 FILLER_3_391 ();
 sg13g2_decap_8 FILLER_3_398 ();
 sg13g2_decap_4 FILLER_3_405 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_fill_2 FILLER_4_42 ();
 sg13g2_fill_1 FILLER_4_69 ();
 sg13g2_fill_1 FILLER_4_93 ();
 sg13g2_decap_8 FILLER_4_102 ();
 sg13g2_decap_8 FILLER_4_150 ();
 sg13g2_decap_8 FILLER_4_157 ();
 sg13g2_decap_8 FILLER_4_164 ();
 sg13g2_decap_4 FILLER_4_171 ();
 sg13g2_decap_8 FILLER_4_188 ();
 sg13g2_fill_1 FILLER_4_195 ();
 sg13g2_decap_8 FILLER_4_204 ();
 sg13g2_decap_8 FILLER_4_211 ();
 sg13g2_decap_8 FILLER_4_218 ();
 sg13g2_fill_1 FILLER_4_225 ();
 sg13g2_fill_2 FILLER_4_256 ();
 sg13g2_fill_1 FILLER_4_258 ();
 sg13g2_fill_1 FILLER_4_264 ();
 sg13g2_fill_2 FILLER_4_283 ();
 sg13g2_fill_2 FILLER_4_295 ();
 sg13g2_fill_2 FILLER_4_304 ();
 sg13g2_fill_2 FILLER_4_319 ();
 sg13g2_decap_8 FILLER_4_360 ();
 sg13g2_decap_8 FILLER_4_367 ();
 sg13g2_decap_8 FILLER_4_374 ();
 sg13g2_decap_8 FILLER_4_381 ();
 sg13g2_decap_8 FILLER_4_388 ();
 sg13g2_decap_8 FILLER_4_395 ();
 sg13g2_decap_8 FILLER_4_402 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_fill_1 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_83 ();
 sg13g2_decap_4 FILLER_5_111 ();
 sg13g2_fill_1 FILLER_5_115 ();
 sg13g2_fill_1 FILLER_5_120 ();
 sg13g2_decap_4 FILLER_5_126 ();
 sg13g2_fill_1 FILLER_5_130 ();
 sg13g2_decap_8 FILLER_5_142 ();
 sg13g2_decap_8 FILLER_5_149 ();
 sg13g2_decap_8 FILLER_5_156 ();
 sg13g2_decap_8 FILLER_5_163 ();
 sg13g2_decap_4 FILLER_5_170 ();
 sg13g2_fill_1 FILLER_5_174 ();
 sg13g2_decap_8 FILLER_5_212 ();
 sg13g2_fill_2 FILLER_5_219 ();
 sg13g2_fill_2 FILLER_5_231 ();
 sg13g2_fill_1 FILLER_5_233 ();
 sg13g2_fill_2 FILLER_5_247 ();
 sg13g2_fill_1 FILLER_5_249 ();
 sg13g2_decap_8 FILLER_5_363 ();
 sg13g2_decap_8 FILLER_5_370 ();
 sg13g2_decap_8 FILLER_5_377 ();
 sg13g2_decap_8 FILLER_5_384 ();
 sg13g2_decap_8 FILLER_5_391 ();
 sg13g2_decap_8 FILLER_5_398 ();
 sg13g2_decap_4 FILLER_5_405 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_4 FILLER_6_28 ();
 sg13g2_fill_1 FILLER_6_53 ();
 sg13g2_fill_2 FILLER_6_71 ();
 sg13g2_fill_1 FILLER_6_73 ();
 sg13g2_fill_1 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_150 ();
 sg13g2_fill_1 FILLER_6_157 ();
 sg13g2_fill_2 FILLER_6_283 ();
 sg13g2_fill_1 FILLER_6_285 ();
 sg13g2_fill_1 FILLER_6_294 ();
 sg13g2_fill_1 FILLER_6_321 ();
 sg13g2_decap_8 FILLER_6_362 ();
 sg13g2_decap_8 FILLER_6_369 ();
 sg13g2_decap_8 FILLER_6_376 ();
 sg13g2_decap_8 FILLER_6_383 ();
 sg13g2_decap_8 FILLER_6_390 ();
 sg13g2_decap_8 FILLER_6_397 ();
 sg13g2_decap_4 FILLER_6_404 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_4 FILLER_7_35 ();
 sg13g2_fill_1 FILLER_7_39 ();
 sg13g2_fill_1 FILLER_7_51 ();
 sg13g2_fill_2 FILLER_7_59 ();
 sg13g2_fill_2 FILLER_7_93 ();
 sg13g2_fill_2 FILLER_7_100 ();
 sg13g2_fill_2 FILLER_7_107 ();
 sg13g2_fill_1 FILLER_7_146 ();
 sg13g2_fill_2 FILLER_7_220 ();
 sg13g2_fill_2 FILLER_7_275 ();
 sg13g2_fill_1 FILLER_7_277 ();
 sg13g2_fill_1 FILLER_7_294 ();
 sg13g2_fill_1 FILLER_7_326 ();
 sg13g2_decap_8 FILLER_7_370 ();
 sg13g2_decap_8 FILLER_7_377 ();
 sg13g2_decap_8 FILLER_7_384 ();
 sg13g2_decap_8 FILLER_7_391 ();
 sg13g2_decap_8 FILLER_7_398 ();
 sg13g2_decap_4 FILLER_7_405 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_fill_2 FILLER_8_49 ();
 sg13g2_fill_1 FILLER_8_51 ();
 sg13g2_decap_4 FILLER_8_56 ();
 sg13g2_decap_4 FILLER_8_69 ();
 sg13g2_fill_2 FILLER_8_79 ();
 sg13g2_fill_1 FILLER_8_121 ();
 sg13g2_decap_8 FILLER_8_158 ();
 sg13g2_fill_2 FILLER_8_165 ();
 sg13g2_fill_1 FILLER_8_167 ();
 sg13g2_fill_2 FILLER_8_185 ();
 sg13g2_fill_2 FILLER_8_230 ();
 sg13g2_fill_1 FILLER_8_280 ();
 sg13g2_fill_1 FILLER_8_287 ();
 sg13g2_fill_2 FILLER_8_333 ();
 sg13g2_decap_8 FILLER_8_358 ();
 sg13g2_decap_8 FILLER_8_365 ();
 sg13g2_decap_8 FILLER_8_372 ();
 sg13g2_decap_8 FILLER_8_379 ();
 sg13g2_decap_8 FILLER_8_386 ();
 sg13g2_decap_8 FILLER_8_393 ();
 sg13g2_decap_8 FILLER_8_400 ();
 sg13g2_fill_2 FILLER_8_407 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_fill_1 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_55 ();
 sg13g2_decap_8 FILLER_9_62 ();
 sg13g2_fill_2 FILLER_9_69 ();
 sg13g2_decap_8 FILLER_9_74 ();
 sg13g2_decap_8 FILLER_9_81 ();
 sg13g2_fill_2 FILLER_9_88 ();
 sg13g2_fill_1 FILLER_9_102 ();
 sg13g2_decap_8 FILLER_9_124 ();
 sg13g2_fill_2 FILLER_9_131 ();
 sg13g2_fill_1 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_141 ();
 sg13g2_decap_4 FILLER_9_148 ();
 sg13g2_fill_1 FILLER_9_152 ();
 sg13g2_decap_4 FILLER_9_158 ();
 sg13g2_fill_2 FILLER_9_170 ();
 sg13g2_fill_1 FILLER_9_195 ();
 sg13g2_fill_1 FILLER_9_225 ();
 sg13g2_fill_1 FILLER_9_248 ();
 sg13g2_fill_2 FILLER_9_327 ();
 sg13g2_decap_8 FILLER_9_366 ();
 sg13g2_decap_8 FILLER_9_373 ();
 sg13g2_decap_8 FILLER_9_380 ();
 sg13g2_decap_8 FILLER_9_387 ();
 sg13g2_decap_8 FILLER_9_394 ();
 sg13g2_decap_8 FILLER_9_401 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_4 FILLER_10_35 ();
 sg13g2_fill_1 FILLER_10_39 ();
 sg13g2_fill_2 FILLER_10_62 ();
 sg13g2_fill_1 FILLER_10_64 ();
 sg13g2_fill_2 FILLER_10_69 ();
 sg13g2_fill_1 FILLER_10_71 ();
 sg13g2_decap_8 FILLER_10_82 ();
 sg13g2_decap_4 FILLER_10_89 ();
 sg13g2_fill_2 FILLER_10_93 ();
 sg13g2_decap_4 FILLER_10_99 ();
 sg13g2_fill_1 FILLER_10_103 ();
 sg13g2_decap_8 FILLER_10_130 ();
 sg13g2_decap_4 FILLER_10_137 ();
 sg13g2_fill_2 FILLER_10_209 ();
 sg13g2_fill_2 FILLER_10_249 ();
 sg13g2_fill_1 FILLER_10_278 ();
 sg13g2_fill_2 FILLER_10_333 ();
 sg13g2_decap_8 FILLER_10_365 ();
 sg13g2_decap_8 FILLER_10_372 ();
 sg13g2_decap_8 FILLER_10_379 ();
 sg13g2_decap_8 FILLER_10_386 ();
 sg13g2_decap_8 FILLER_10_393 ();
 sg13g2_decap_8 FILLER_10_400 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_fill_1 FILLER_11_65 ();
 sg13g2_fill_1 FILLER_11_110 ();
 sg13g2_fill_2 FILLER_11_123 ();
 sg13g2_fill_1 FILLER_11_125 ();
 sg13g2_decap_8 FILLER_11_138 ();
 sg13g2_decap_4 FILLER_11_145 ();
 sg13g2_fill_1 FILLER_11_149 ();
 sg13g2_fill_2 FILLER_11_158 ();
 sg13g2_fill_1 FILLER_11_160 ();
 sg13g2_fill_2 FILLER_11_197 ();
 sg13g2_fill_2 FILLER_11_212 ();
 sg13g2_fill_2 FILLER_11_270 ();
 sg13g2_fill_1 FILLER_11_272 ();
 sg13g2_fill_2 FILLER_11_278 ();
 sg13g2_fill_1 FILLER_11_335 ();
 sg13g2_fill_1 FILLER_11_341 ();
 sg13g2_decap_8 FILLER_11_368 ();
 sg13g2_decap_8 FILLER_11_375 ();
 sg13g2_decap_8 FILLER_11_382 ();
 sg13g2_decap_8 FILLER_11_389 ();
 sg13g2_decap_8 FILLER_11_396 ();
 sg13g2_decap_4 FILLER_11_403 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_4 FILLER_12_35 ();
 sg13g2_fill_1 FILLER_12_63 ();
 sg13g2_decap_4 FILLER_12_97 ();
 sg13g2_fill_1 FILLER_12_117 ();
 sg13g2_fill_1 FILLER_12_128 ();
 sg13g2_fill_1 FILLER_12_142 ();
 sg13g2_fill_2 FILLER_12_169 ();
 sg13g2_fill_1 FILLER_12_171 ();
 sg13g2_fill_1 FILLER_12_190 ();
 sg13g2_fill_2 FILLER_12_284 ();
 sg13g2_fill_1 FILLER_12_286 ();
 sg13g2_fill_1 FILLER_12_339 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_4 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_85 ();
 sg13g2_fill_1 FILLER_13_115 ();
 sg13g2_fill_2 FILLER_13_122 ();
 sg13g2_fill_1 FILLER_13_124 ();
 sg13g2_decap_4 FILLER_13_130 ();
 sg13g2_fill_2 FILLER_13_134 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_fill_1 FILLER_13_203 ();
 sg13g2_fill_2 FILLER_13_227 ();
 sg13g2_fill_1 FILLER_13_229 ();
 sg13g2_fill_2 FILLER_13_242 ();
 sg13g2_fill_1 FILLER_13_339 ();
 sg13g2_decap_8 FILLER_13_374 ();
 sg13g2_decap_8 FILLER_13_381 ();
 sg13g2_decap_8 FILLER_13_388 ();
 sg13g2_decap_8 FILLER_13_395 ();
 sg13g2_decap_8 FILLER_13_402 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_4 FILLER_14_91 ();
 sg13g2_fill_2 FILLER_14_95 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_4 FILLER_14_123 ();
 sg13g2_fill_1 FILLER_14_171 ();
 sg13g2_fill_1 FILLER_14_219 ();
 sg13g2_fill_2 FILLER_14_248 ();
 sg13g2_fill_2 FILLER_14_258 ();
 sg13g2_fill_1 FILLER_14_300 ();
 sg13g2_fill_2 FILLER_14_325 ();
 sg13g2_decap_8 FILLER_14_370 ();
 sg13g2_decap_8 FILLER_14_377 ();
 sg13g2_decap_8 FILLER_14_384 ();
 sg13g2_decap_8 FILLER_14_391 ();
 sg13g2_decap_8 FILLER_14_398 ();
 sg13g2_decap_4 FILLER_14_405 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_4 FILLER_15_61 ();
 sg13g2_fill_2 FILLER_15_69 ();
 sg13g2_fill_1 FILLER_15_71 ();
 sg13g2_fill_2 FILLER_15_99 ();
 sg13g2_decap_8 FILLER_15_109 ();
 sg13g2_decap_8 FILLER_15_116 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_fill_2 FILLER_15_224 ();
 sg13g2_fill_1 FILLER_15_226 ();
 sg13g2_fill_1 FILLER_15_269 ();
 sg13g2_fill_1 FILLER_15_300 ();
 sg13g2_decap_8 FILLER_15_379 ();
 sg13g2_decap_8 FILLER_15_386 ();
 sg13g2_decap_8 FILLER_15_393 ();
 sg13g2_decap_8 FILLER_15_400 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_fill_2 FILLER_16_42 ();
 sg13g2_fill_2 FILLER_16_65 ();
 sg13g2_fill_2 FILLER_16_78 ();
 sg13g2_fill_2 FILLER_16_88 ();
 sg13g2_fill_2 FILLER_16_96 ();
 sg13g2_fill_1 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_fill_2 FILLER_16_155 ();
 sg13g2_decap_8 FILLER_16_172 ();
 sg13g2_decap_8 FILLER_16_179 ();
 sg13g2_fill_2 FILLER_16_186 ();
 sg13g2_fill_2 FILLER_16_223 ();
 sg13g2_fill_1 FILLER_16_225 ();
 sg13g2_fill_2 FILLER_16_239 ();
 sg13g2_fill_1 FILLER_16_241 ();
 sg13g2_fill_2 FILLER_16_251 ();
 sg13g2_fill_1 FILLER_16_253 ();
 sg13g2_fill_2 FILLER_16_286 ();
 sg13g2_fill_2 FILLER_16_348 ();
 sg13g2_decap_8 FILLER_16_380 ();
 sg13g2_decap_8 FILLER_16_387 ();
 sg13g2_decap_8 FILLER_16_394 ();
 sg13g2_decap_8 FILLER_16_401 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_fill_2 FILLER_17_52 ();
 sg13g2_fill_1 FILLER_17_88 ();
 sg13g2_decap_4 FILLER_17_116 ();
 sg13g2_decap_4 FILLER_17_156 ();
 sg13g2_fill_1 FILLER_17_160 ();
 sg13g2_decap_4 FILLER_17_177 ();
 sg13g2_fill_1 FILLER_17_181 ();
 sg13g2_fill_2 FILLER_17_320 ();
 sg13g2_fill_1 FILLER_17_332 ();
 sg13g2_fill_1 FILLER_17_338 ();
 sg13g2_fill_2 FILLER_17_348 ();
 sg13g2_fill_1 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_377 ();
 sg13g2_decap_8 FILLER_17_384 ();
 sg13g2_decap_8 FILLER_17_391 ();
 sg13g2_decap_8 FILLER_17_398 ();
 sg13g2_decap_4 FILLER_17_405 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_4 FILLER_18_35 ();
 sg13g2_fill_1 FILLER_18_39 ();
 sg13g2_fill_1 FILLER_18_51 ();
 sg13g2_fill_1 FILLER_18_66 ();
 sg13g2_decap_8 FILLER_18_92 ();
 sg13g2_decap_4 FILLER_18_99 ();
 sg13g2_fill_2 FILLER_18_103 ();
 sg13g2_decap_8 FILLER_18_114 ();
 sg13g2_fill_1 FILLER_18_121 ();
 sg13g2_decap_8 FILLER_18_137 ();
 sg13g2_fill_1 FILLER_18_250 ();
 sg13g2_fill_2 FILLER_18_284 ();
 sg13g2_fill_1 FILLER_18_286 ();
 sg13g2_fill_1 FILLER_18_323 ();
 sg13g2_fill_2 FILLER_18_329 ();
 sg13g2_fill_2 FILLER_18_357 ();
 sg13g2_fill_1 FILLER_18_359 ();
 sg13g2_decap_8 FILLER_18_377 ();
 sg13g2_decap_8 FILLER_18_384 ();
 sg13g2_decap_8 FILLER_18_391 ();
 sg13g2_decap_8 FILLER_18_398 ();
 sg13g2_decap_4 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_fill_1 FILLER_19_49 ();
 sg13g2_fill_2 FILLER_19_55 ();
 sg13g2_fill_1 FILLER_19_57 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_fill_2 FILLER_19_91 ();
 sg13g2_fill_2 FILLER_19_108 ();
 sg13g2_fill_1 FILLER_19_110 ();
 sg13g2_fill_2 FILLER_19_116 ();
 sg13g2_fill_1 FILLER_19_168 ();
 sg13g2_decap_4 FILLER_19_177 ();
 sg13g2_decap_4 FILLER_19_186 ();
 sg13g2_fill_1 FILLER_19_208 ();
 sg13g2_fill_1 FILLER_19_313 ();
 sg13g2_fill_1 FILLER_19_342 ();
 sg13g2_decap_8 FILLER_19_352 ();
 sg13g2_decap_8 FILLER_19_359 ();
 sg13g2_fill_2 FILLER_19_366 ();
 sg13g2_fill_1 FILLER_19_368 ();
 sg13g2_decap_4 FILLER_19_379 ();
 sg13g2_fill_1 FILLER_19_383 ();
 sg13g2_fill_2 FILLER_19_388 ();
 sg13g2_decap_8 FILLER_19_395 ();
 sg13g2_decap_8 FILLER_19_402 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_4 FILLER_20_49 ();
 sg13g2_fill_1 FILLER_20_66 ();
 sg13g2_fill_2 FILLER_20_72 ();
 sg13g2_fill_2 FILLER_20_118 ();
 sg13g2_fill_2 FILLER_20_164 ();
 sg13g2_fill_2 FILLER_20_214 ();
 sg13g2_fill_1 FILLER_20_216 ();
 sg13g2_fill_2 FILLER_20_286 ();
 sg13g2_fill_1 FILLER_20_288 ();
 sg13g2_decap_8 FILLER_20_326 ();
 sg13g2_decap_8 FILLER_20_333 ();
 sg13g2_decap_8 FILLER_20_340 ();
 sg13g2_decap_8 FILLER_20_347 ();
 sg13g2_fill_2 FILLER_20_354 ();
 sg13g2_fill_2 FILLER_20_366 ();
 sg13g2_fill_1 FILLER_20_368 ();
 sg13g2_fill_1 FILLER_20_374 ();
 sg13g2_fill_2 FILLER_20_401 ();
 sg13g2_fill_1 FILLER_20_403 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_4 FILLER_21_42 ();
 sg13g2_fill_1 FILLER_21_55 ();
 sg13g2_fill_2 FILLER_21_64 ();
 sg13g2_fill_1 FILLER_21_82 ();
 sg13g2_fill_2 FILLER_21_161 ();
 sg13g2_fill_2 FILLER_21_178 ();
 sg13g2_fill_2 FILLER_21_189 ();
 sg13g2_fill_1 FILLER_21_191 ();
 sg13g2_fill_2 FILLER_21_201 ();
 sg13g2_fill_1 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_213 ();
 sg13g2_fill_2 FILLER_21_228 ();
 sg13g2_fill_1 FILLER_21_285 ();
 sg13g2_decap_4 FILLER_21_303 ();
 sg13g2_fill_2 FILLER_21_307 ();
 sg13g2_decap_4 FILLER_21_328 ();
 sg13g2_fill_1 FILLER_21_332 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_fill_1 FILLER_22_42 ();
 sg13g2_fill_2 FILLER_22_59 ();
 sg13g2_fill_2 FILLER_22_154 ();
 sg13g2_fill_2 FILLER_22_159 ();
 sg13g2_fill_1 FILLER_22_165 ();
 sg13g2_decap_8 FILLER_22_212 ();
 sg13g2_fill_2 FILLER_22_219 ();
 sg13g2_fill_2 FILLER_22_225 ();
 sg13g2_fill_1 FILLER_22_227 ();
 sg13g2_fill_2 FILLER_22_254 ();
 sg13g2_fill_2 FILLER_22_261 ();
 sg13g2_decap_4 FILLER_22_301 ();
 sg13g2_fill_2 FILLER_22_353 ();
 sg13g2_fill_1 FILLER_22_355 ();
 sg13g2_fill_1 FILLER_22_364 ();
 sg13g2_fill_2 FILLER_22_373 ();
 sg13g2_fill_1 FILLER_22_375 ();
 sg13g2_fill_2 FILLER_22_383 ();
 sg13g2_fill_1 FILLER_22_385 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_4 FILLER_23_42 ();
 sg13g2_fill_2 FILLER_23_46 ();
 sg13g2_fill_2 FILLER_23_65 ();
 sg13g2_fill_2 FILLER_23_80 ();
 sg13g2_fill_1 FILLER_23_82 ();
 sg13g2_fill_2 FILLER_23_88 ();
 sg13g2_fill_1 FILLER_23_90 ();
 sg13g2_fill_2 FILLER_23_96 ();
 sg13g2_decap_8 FILLER_23_107 ();
 sg13g2_fill_2 FILLER_23_114 ();
 sg13g2_fill_1 FILLER_23_116 ();
 sg13g2_fill_2 FILLER_23_141 ();
 sg13g2_fill_1 FILLER_23_143 ();
 sg13g2_fill_1 FILLER_23_149 ();
 sg13g2_decap_8 FILLER_23_162 ();
 sg13g2_decap_4 FILLER_23_169 ();
 sg13g2_fill_2 FILLER_23_173 ();
 sg13g2_fill_2 FILLER_23_183 ();
 sg13g2_fill_1 FILLER_23_185 ();
 sg13g2_decap_4 FILLER_23_226 ();
 sg13g2_fill_2 FILLER_23_256 ();
 sg13g2_decap_4 FILLER_23_284 ();
 sg13g2_fill_2 FILLER_23_288 ();
 sg13g2_decap_4 FILLER_23_303 ();
 sg13g2_fill_2 FILLER_23_344 ();
 sg13g2_fill_1 FILLER_23_363 ();
 sg13g2_fill_1 FILLER_23_379 ();
 sg13g2_fill_1 FILLER_23_404 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_4 FILLER_24_49 ();
 sg13g2_fill_1 FILLER_24_53 ();
 sg13g2_fill_1 FILLER_24_79 ();
 sg13g2_decap_8 FILLER_24_92 ();
 sg13g2_fill_2 FILLER_24_99 ();
 sg13g2_fill_1 FILLER_24_101 ();
 sg13g2_fill_2 FILLER_24_120 ();
 sg13g2_fill_1 FILLER_24_122 ();
 sg13g2_fill_1 FILLER_24_163 ();
 sg13g2_fill_1 FILLER_24_180 ();
 sg13g2_fill_2 FILLER_24_185 ();
 sg13g2_fill_1 FILLER_24_187 ();
 sg13g2_fill_2 FILLER_24_232 ();
 sg13g2_fill_2 FILLER_24_290 ();
 sg13g2_fill_1 FILLER_24_308 ();
 sg13g2_decap_4 FILLER_24_314 ();
 sg13g2_fill_1 FILLER_24_326 ();
 sg13g2_decap_4 FILLER_24_336 ();
 sg13g2_fill_1 FILLER_24_340 ();
 sg13g2_fill_1 FILLER_24_373 ();
 sg13g2_fill_2 FILLER_24_387 ();
 sg13g2_fill_2 FILLER_24_394 ();
 sg13g2_fill_1 FILLER_24_396 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_fill_1 FILLER_25_35 ();
 sg13g2_fill_2 FILLER_25_62 ();
 sg13g2_fill_1 FILLER_25_64 ();
 sg13g2_decap_4 FILLER_25_95 ();
 sg13g2_fill_2 FILLER_25_99 ();
 sg13g2_fill_2 FILLER_25_109 ();
 sg13g2_fill_1 FILLER_25_111 ();
 sg13g2_fill_1 FILLER_25_126 ();
 sg13g2_decap_4 FILLER_25_143 ();
 sg13g2_fill_2 FILLER_25_183 ();
 sg13g2_decap_8 FILLER_25_195 ();
 sg13g2_decap_8 FILLER_25_202 ();
 sg13g2_decap_8 FILLER_25_209 ();
 sg13g2_fill_1 FILLER_25_216 ();
 sg13g2_fill_2 FILLER_25_235 ();
 sg13g2_fill_1 FILLER_25_237 ();
 sg13g2_fill_1 FILLER_25_247 ();
 sg13g2_fill_2 FILLER_25_261 ();
 sg13g2_fill_1 FILLER_25_263 ();
 sg13g2_fill_1 FILLER_25_277 ();
 sg13g2_fill_1 FILLER_25_286 ();
 sg13g2_decap_8 FILLER_25_295 ();
 sg13g2_decap_4 FILLER_25_302 ();
 sg13g2_fill_2 FILLER_25_306 ();
 sg13g2_decap_8 FILLER_25_316 ();
 sg13g2_decap_8 FILLER_25_323 ();
 sg13g2_fill_2 FILLER_25_330 ();
 sg13g2_decap_8 FILLER_25_360 ();
 sg13g2_fill_1 FILLER_25_367 ();
 sg13g2_decap_8 FILLER_25_372 ();
 sg13g2_fill_2 FILLER_25_379 ();
 sg13g2_fill_1 FILLER_25_392 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_4 FILLER_26_42 ();
 sg13g2_fill_1 FILLER_26_46 ();
 sg13g2_decap_4 FILLER_26_51 ();
 sg13g2_fill_1 FILLER_26_72 ();
 sg13g2_fill_2 FILLER_26_122 ();
 sg13g2_fill_1 FILLER_26_124 ();
 sg13g2_fill_2 FILLER_26_132 ();
 sg13g2_fill_1 FILLER_26_142 ();
 sg13g2_fill_1 FILLER_26_219 ();
 sg13g2_decap_8 FILLER_26_277 ();
 sg13g2_fill_1 FILLER_26_297 ();
 sg13g2_decap_8 FILLER_26_306 ();
 sg13g2_fill_1 FILLER_26_313 ();
 sg13g2_fill_1 FILLER_26_333 ();
 sg13g2_fill_1 FILLER_26_362 ();
 sg13g2_decap_4 FILLER_26_375 ();
 sg13g2_fill_2 FILLER_26_379 ();
 sg13g2_fill_2 FILLER_26_400 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_fill_1 FILLER_27_56 ();
 sg13g2_fill_1 FILLER_27_87 ();
 sg13g2_fill_1 FILLER_27_100 ();
 sg13g2_fill_1 FILLER_27_118 ();
 sg13g2_fill_2 FILLER_27_127 ();
 sg13g2_fill_1 FILLER_27_144 ();
 sg13g2_fill_2 FILLER_27_173 ();
 sg13g2_fill_1 FILLER_27_195 ();
 sg13g2_fill_1 FILLER_27_221 ();
 sg13g2_fill_1 FILLER_27_228 ();
 sg13g2_decap_8 FILLER_27_262 ();
 sg13g2_fill_1 FILLER_27_269 ();
 sg13g2_fill_1 FILLER_27_278 ();
 sg13g2_decap_4 FILLER_27_311 ();
 sg13g2_fill_1 FILLER_27_315 ();
 sg13g2_fill_1 FILLER_27_334 ();
 sg13g2_fill_2 FILLER_27_372 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_4 FILLER_28_28 ();
 sg13g2_fill_1 FILLER_28_32 ();
 sg13g2_decap_8 FILLER_28_73 ();
 sg13g2_fill_2 FILLER_28_80 ();
 sg13g2_fill_1 FILLER_28_82 ();
 sg13g2_fill_2 FILLER_28_92 ();
 sg13g2_decap_4 FILLER_28_103 ();
 sg13g2_decap_4 FILLER_28_121 ();
 sg13g2_fill_2 FILLER_28_144 ();
 sg13g2_fill_1 FILLER_28_166 ();
 sg13g2_fill_1 FILLER_28_178 ();
 sg13g2_fill_2 FILLER_28_188 ();
 sg13g2_fill_2 FILLER_28_216 ();
 sg13g2_fill_1 FILLER_28_218 ();
 sg13g2_decap_4 FILLER_28_222 ();
 sg13g2_fill_2 FILLER_28_226 ();
 sg13g2_decap_4 FILLER_28_241 ();
 sg13g2_fill_2 FILLER_28_250 ();
 sg13g2_fill_1 FILLER_28_252 ();
 sg13g2_decap_8 FILLER_28_292 ();
 sg13g2_decap_4 FILLER_28_299 ();
 sg13g2_fill_2 FILLER_28_303 ();
 sg13g2_fill_1 FILLER_28_310 ();
 sg13g2_fill_1 FILLER_28_326 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_fill_2 FILLER_29_28 ();
 sg13g2_fill_2 FILLER_29_65 ();
 sg13g2_decap_4 FILLER_29_132 ();
 sg13g2_fill_1 FILLER_29_141 ();
 sg13g2_decap_8 FILLER_29_146 ();
 sg13g2_fill_1 FILLER_29_153 ();
 sg13g2_decap_4 FILLER_29_163 ();
 sg13g2_decap_4 FILLER_29_172 ();
 sg13g2_fill_2 FILLER_29_179 ();
 sg13g2_fill_1 FILLER_29_211 ();
 sg13g2_fill_2 FILLER_29_231 ();
 sg13g2_fill_1 FILLER_29_233 ();
 sg13g2_decap_8 FILLER_29_264 ();
 sg13g2_decap_8 FILLER_29_271 ();
 sg13g2_fill_2 FILLER_29_278 ();
 sg13g2_fill_2 FILLER_29_298 ();
 sg13g2_fill_2 FILLER_29_345 ();
 sg13g2_fill_1 FILLER_29_347 ();
 sg13g2_fill_2 FILLER_29_374 ();
 sg13g2_decap_8 FILLER_29_380 ();
 sg13g2_fill_2 FILLER_29_387 ();
 sg13g2_fill_1 FILLER_29_389 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_4 FILLER_30_28 ();
 sg13g2_fill_2 FILLER_30_32 ();
 sg13g2_fill_2 FILLER_30_54 ();
 sg13g2_decap_4 FILLER_30_61 ();
 sg13g2_fill_2 FILLER_30_75 ();
 sg13g2_fill_2 FILLER_30_112 ();
 sg13g2_fill_1 FILLER_30_114 ();
 sg13g2_decap_8 FILLER_30_149 ();
 sg13g2_decap_8 FILLER_30_156 ();
 sg13g2_decap_8 FILLER_30_181 ();
 sg13g2_decap_4 FILLER_30_188 ();
 sg13g2_fill_2 FILLER_30_227 ();
 sg13g2_fill_1 FILLER_30_229 ();
 sg13g2_fill_1 FILLER_30_273 ();
 sg13g2_decap_8 FILLER_30_301 ();
 sg13g2_decap_4 FILLER_30_308 ();
 sg13g2_fill_2 FILLER_30_324 ();
 sg13g2_fill_1 FILLER_30_331 ();
 sg13g2_decap_8 FILLER_30_348 ();
 sg13g2_decap_8 FILLER_30_355 ();
 sg13g2_decap_4 FILLER_30_362 ();
 sg13g2_fill_2 FILLER_30_366 ();
 sg13g2_fill_1 FILLER_30_376 ();
 sg13g2_fill_1 FILLER_30_388 ();
 sg13g2_fill_2 FILLER_30_402 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_4 FILLER_31_42 ();
 sg13g2_decap_4 FILLER_31_67 ();
 sg13g2_fill_2 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_134 ();
 sg13g2_decap_4 FILLER_31_141 ();
 sg13g2_fill_1 FILLER_31_145 ();
 sg13g2_decap_4 FILLER_31_150 ();
 sg13g2_fill_1 FILLER_31_154 ();
 sg13g2_fill_2 FILLER_31_186 ();
 sg13g2_fill_2 FILLER_31_226 ();
 sg13g2_fill_1 FILLER_31_228 ();
 sg13g2_fill_1 FILLER_31_273 ();
 sg13g2_fill_2 FILLER_31_282 ();
 sg13g2_decap_8 FILLER_31_303 ();
 sg13g2_decap_4 FILLER_31_310 ();
 sg13g2_fill_2 FILLER_31_337 ();
 sg13g2_fill_2 FILLER_31_349 ();
 sg13g2_fill_1 FILLER_31_351 ();
 sg13g2_decap_8 FILLER_31_356 ();
 sg13g2_fill_1 FILLER_31_363 ();
 sg13g2_fill_1 FILLER_31_381 ();
 sg13g2_decap_4 FILLER_31_389 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_4 FILLER_32_35 ();
 sg13g2_fill_1 FILLER_32_39 ();
 sg13g2_decap_4 FILLER_32_49 ();
 sg13g2_fill_2 FILLER_32_56 ();
 sg13g2_fill_1 FILLER_32_58 ();
 sg13g2_decap_8 FILLER_32_68 ();
 sg13g2_fill_2 FILLER_32_75 ();
 sg13g2_fill_1 FILLER_32_77 ();
 sg13g2_fill_1 FILLER_32_92 ();
 sg13g2_fill_2 FILLER_32_121 ();
 sg13g2_fill_2 FILLER_32_127 ();
 sg13g2_fill_1 FILLER_32_134 ();
 sg13g2_fill_2 FILLER_32_161 ();
 sg13g2_fill_1 FILLER_32_180 ();
 sg13g2_fill_1 FILLER_32_237 ();
 sg13g2_fill_1 FILLER_32_251 ();
 sg13g2_fill_2 FILLER_32_266 ();
 sg13g2_decap_4 FILLER_32_302 ();
 sg13g2_fill_1 FILLER_32_306 ();
 sg13g2_fill_2 FILLER_32_335 ();
 sg13g2_fill_1 FILLER_32_350 ();
 sg13g2_fill_2 FILLER_32_384 ();
 sg13g2_fill_1 FILLER_32_386 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_fill_2 FILLER_33_28 ();
 sg13g2_fill_1 FILLER_33_30 ();
 sg13g2_fill_2 FILLER_33_112 ();
 sg13g2_fill_1 FILLER_33_114 ();
 sg13g2_fill_2 FILLER_33_132 ();
 sg13g2_fill_1 FILLER_33_186 ();
 sg13g2_fill_1 FILLER_33_200 ();
 sg13g2_fill_1 FILLER_33_226 ();
 sg13g2_fill_2 FILLER_33_240 ();
 sg13g2_fill_1 FILLER_33_252 ();
 sg13g2_fill_2 FILLER_33_266 ();
 sg13g2_fill_2 FILLER_33_290 ();
 sg13g2_decap_8 FILLER_33_297 ();
 sg13g2_fill_2 FILLER_33_304 ();
 sg13g2_decap_8 FILLER_33_318 ();
 sg13g2_fill_2 FILLER_33_325 ();
 sg13g2_fill_1 FILLER_33_363 ();
 sg13g2_decap_4 FILLER_33_386 ();
 sg13g2_fill_1 FILLER_33_390 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_4 FILLER_34_21 ();
 sg13g2_fill_1 FILLER_34_25 ();
 sg13g2_fill_1 FILLER_34_78 ();
 sg13g2_fill_2 FILLER_34_141 ();
 sg13g2_fill_1 FILLER_34_143 ();
 sg13g2_fill_1 FILLER_34_177 ();
 sg13g2_fill_2 FILLER_34_227 ();
 sg13g2_fill_1 FILLER_34_229 ();
 sg13g2_decap_4 FILLER_34_288 ();
 sg13g2_fill_2 FILLER_34_292 ();
 sg13g2_decap_4 FILLER_34_319 ();
 sg13g2_decap_4 FILLER_34_327 ();
 sg13g2_fill_2 FILLER_34_337 ();
 sg13g2_decap_4 FILLER_34_347 ();
 sg13g2_fill_1 FILLER_34_351 ();
 sg13g2_decap_4 FILLER_34_379 ();
 sg13g2_fill_2 FILLER_34_383 ();
 sg13g2_fill_2 FILLER_34_389 ();
 sg13g2_fill_1 FILLER_34_391 ();
 sg13g2_decap_8 FILLER_34_401 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_fill_2 FILLER_35_35 ();
 sg13g2_fill_1 FILLER_35_37 ();
 sg13g2_fill_1 FILLER_35_65 ();
 sg13g2_fill_1 FILLER_35_80 ();
 sg13g2_fill_1 FILLER_35_144 ();
 sg13g2_fill_1 FILLER_35_173 ();
 sg13g2_fill_2 FILLER_35_182 ();
 sg13g2_fill_1 FILLER_35_187 ();
 sg13g2_fill_2 FILLER_35_191 ();
 sg13g2_fill_2 FILLER_35_197 ();
 sg13g2_fill_1 FILLER_35_199 ();
 sg13g2_decap_4 FILLER_35_282 ();
 sg13g2_fill_2 FILLER_35_286 ();
 sg13g2_fill_1 FILLER_35_310 ();
 sg13g2_fill_1 FILLER_35_329 ();
 sg13g2_decap_4 FILLER_35_355 ();
 sg13g2_fill_1 FILLER_35_379 ();
 sg13g2_fill_1 FILLER_35_386 ();
 sg13g2_fill_1 FILLER_35_394 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_fill_2 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_4 FILLER_36_63 ();
 sg13g2_fill_2 FILLER_36_153 ();
 sg13g2_fill_1 FILLER_36_184 ();
 sg13g2_decap_8 FILLER_36_194 ();
 sg13g2_fill_2 FILLER_36_201 ();
 sg13g2_fill_1 FILLER_36_203 ();
 sg13g2_fill_2 FILLER_36_212 ();
 sg13g2_fill_2 FILLER_36_264 ();
 sg13g2_fill_2 FILLER_36_351 ();
 sg13g2_decap_4 FILLER_36_363 ();
 sg13g2_fill_1 FILLER_36_367 ();
 sg13g2_fill_2 FILLER_36_378 ();
 sg13g2_fill_1 FILLER_36_380 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_fill_1 FILLER_37_56 ();
 sg13g2_fill_1 FILLER_37_111 ();
 sg13g2_fill_2 FILLER_37_122 ();
 sg13g2_fill_2 FILLER_37_142 ();
 sg13g2_fill_1 FILLER_37_149 ();
 sg13g2_fill_1 FILLER_37_169 ();
 sg13g2_decap_8 FILLER_37_204 ();
 sg13g2_fill_1 FILLER_37_288 ();
 sg13g2_decap_8 FILLER_37_341 ();
 sg13g2_fill_1 FILLER_37_348 ();
 sg13g2_fill_1 FILLER_37_353 ();
 sg13g2_decap_4 FILLER_37_366 ();
 sg13g2_fill_1 FILLER_37_377 ();
 sg13g2_fill_2 FILLER_37_384 ();
 sg13g2_fill_2 FILLER_37_391 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_4 FILLER_38_35 ();
 sg13g2_fill_1 FILLER_38_39 ();
 sg13g2_fill_2 FILLER_38_75 ();
 sg13g2_decap_8 FILLER_38_82 ();
 sg13g2_decap_4 FILLER_38_93 ();
 sg13g2_fill_2 FILLER_38_105 ();
 sg13g2_fill_1 FILLER_38_118 ();
 sg13g2_fill_1 FILLER_38_124 ();
 sg13g2_fill_2 FILLER_38_130 ();
 sg13g2_fill_1 FILLER_38_214 ();
 sg13g2_fill_2 FILLER_38_239 ();
 sg13g2_fill_1 FILLER_38_241 ();
 sg13g2_decap_4 FILLER_38_290 ();
 sg13g2_fill_2 FILLER_38_294 ();
 sg13g2_decap_8 FILLER_38_305 ();
 sg13g2_decap_8 FILLER_38_312 ();
 sg13g2_decap_4 FILLER_38_319 ();
 sg13g2_fill_2 FILLER_38_323 ();
 sg13g2_decap_8 FILLER_38_332 ();
 sg13g2_decap_8 FILLER_38_339 ();
 sg13g2_decap_4 FILLER_38_346 ();
 sg13g2_decap_8 FILLER_38_362 ();
 sg13g2_decap_8 FILLER_38_369 ();
 sg13g2_decap_4 FILLER_38_376 ();
 sg13g2_fill_1 FILLER_38_380 ();
 sg13g2_decap_8 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_4 FILLER_39_35 ();
 sg13g2_decap_4 FILLER_39_86 ();
 sg13g2_fill_2 FILLER_39_100 ();
 sg13g2_fill_1 FILLER_39_128 ();
 sg13g2_fill_2 FILLER_39_174 ();
 sg13g2_fill_2 FILLER_39_185 ();
 sg13g2_decap_4 FILLER_39_273 ();
 sg13g2_fill_2 FILLER_39_277 ();
 sg13g2_decap_4 FILLER_39_295 ();
 sg13g2_fill_1 FILLER_39_299 ();
 sg13g2_decap_8 FILLER_39_314 ();
 sg13g2_decap_8 FILLER_39_321 ();
 sg13g2_decap_8 FILLER_39_328 ();
 sg13g2_decap_4 FILLER_39_335 ();
 sg13g2_fill_1 FILLER_39_339 ();
 sg13g2_fill_1 FILLER_39_348 ();
 sg13g2_decap_8 FILLER_39_379 ();
 sg13g2_fill_1 FILLER_39_386 ();
 sg13g2_fill_1 FILLER_39_408 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_fill_1 FILLER_40_60 ();
 sg13g2_fill_1 FILLER_40_90 ();
 sg13g2_fill_2 FILLER_40_113 ();
 sg13g2_fill_2 FILLER_40_159 ();
 sg13g2_fill_1 FILLER_40_191 ();
 sg13g2_decap_8 FILLER_40_224 ();
 sg13g2_fill_2 FILLER_40_231 ();
 sg13g2_fill_2 FILLER_40_253 ();
 sg13g2_fill_1 FILLER_40_333 ();
 sg13g2_fill_2 FILLER_40_346 ();
 sg13g2_fill_2 FILLER_40_366 ();
 sg13g2_fill_1 FILLER_40_368 ();
 sg13g2_fill_1 FILLER_40_384 ();
 sg13g2_fill_2 FILLER_40_406 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_fill_2 FILLER_41_35 ();
 sg13g2_fill_2 FILLER_41_68 ();
 sg13g2_fill_1 FILLER_41_70 ();
 sg13g2_fill_1 FILLER_41_191 ();
 sg13g2_decap_8 FILLER_41_207 ();
 sg13g2_decap_4 FILLER_41_214 ();
 sg13g2_fill_1 FILLER_41_218 ();
 sg13g2_fill_1 FILLER_41_225 ();
 sg13g2_decap_8 FILLER_41_231 ();
 sg13g2_fill_1 FILLER_41_238 ();
 sg13g2_fill_2 FILLER_41_249 ();
 sg13g2_fill_1 FILLER_41_251 ();
 sg13g2_fill_1 FILLER_41_329 ();
 sg13g2_fill_1 FILLER_41_350 ();
 sg13g2_fill_2 FILLER_41_382 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_fill_2 FILLER_42_49 ();
 sg13g2_fill_1 FILLER_42_51 ();
 sg13g2_decap_4 FILLER_42_58 ();
 sg13g2_fill_2 FILLER_42_62 ();
 sg13g2_decap_4 FILLER_42_69 ();
 sg13g2_fill_2 FILLER_42_73 ();
 sg13g2_fill_2 FILLER_42_79 ();
 sg13g2_fill_2 FILLER_42_104 ();
 sg13g2_decap_4 FILLER_42_120 ();
 sg13g2_fill_1 FILLER_42_127 ();
 sg13g2_fill_2 FILLER_42_133 ();
 sg13g2_decap_8 FILLER_42_143 ();
 sg13g2_fill_1 FILLER_42_150 ();
 sg13g2_fill_2 FILLER_42_159 ();
 sg13g2_fill_2 FILLER_42_187 ();
 sg13g2_fill_2 FILLER_42_222 ();
 sg13g2_fill_1 FILLER_42_224 ();
 sg13g2_fill_1 FILLER_42_252 ();
 sg13g2_fill_2 FILLER_42_273 ();
 sg13g2_fill_2 FILLER_42_292 ();
 sg13g2_fill_1 FILLER_42_302 ();
 sg13g2_fill_2 FILLER_42_328 ();
 sg13g2_fill_1 FILLER_42_330 ();
 sg13g2_decap_8 FILLER_42_336 ();
 sg13g2_fill_1 FILLER_42_343 ();
 sg13g2_decap_8 FILLER_42_353 ();
 sg13g2_decap_4 FILLER_42_360 ();
 sg13g2_fill_2 FILLER_42_364 ();
 sg13g2_decap_8 FILLER_42_375 ();
 sg13g2_decap_8 FILLER_42_382 ();
 sg13g2_fill_2 FILLER_42_389 ();
 sg13g2_fill_1 FILLER_42_391 ();
 sg13g2_decap_8 FILLER_42_401 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_fill_1 FILLER_43_42 ();
 sg13g2_fill_2 FILLER_43_56 ();
 sg13g2_fill_1 FILLER_43_61 ();
 sg13g2_decap_8 FILLER_43_67 ();
 sg13g2_decap_8 FILLER_43_74 ();
 sg13g2_decap_4 FILLER_43_84 ();
 sg13g2_fill_1 FILLER_43_88 ();
 sg13g2_fill_2 FILLER_43_94 ();
 sg13g2_fill_1 FILLER_43_96 ();
 sg13g2_decap_4 FILLER_43_138 ();
 sg13g2_fill_2 FILLER_43_142 ();
 sg13g2_fill_2 FILLER_43_153 ();
 sg13g2_fill_1 FILLER_43_258 ();
 sg13g2_decap_8 FILLER_43_298 ();
 sg13g2_fill_2 FILLER_43_305 ();
 sg13g2_fill_1 FILLER_43_307 ();
 sg13g2_decap_4 FILLER_43_311 ();
 sg13g2_fill_1 FILLER_43_315 ();
 sg13g2_decap_8 FILLER_43_322 ();
 sg13g2_decap_8 FILLER_43_329 ();
 sg13g2_decap_8 FILLER_43_351 ();
 sg13g2_fill_2 FILLER_43_358 ();
 sg13g2_fill_1 FILLER_43_360 ();
 sg13g2_decap_4 FILLER_43_378 ();
 sg13g2_decap_8 FILLER_43_393 ();
 sg13g2_decap_8 FILLER_43_400 ();
 sg13g2_fill_2 FILLER_43_407 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_fill_2 FILLER_44_61 ();
 sg13g2_fill_2 FILLER_44_96 ();
 sg13g2_fill_1 FILLER_44_121 ();
 sg13g2_decap_8 FILLER_44_137 ();
 sg13g2_fill_2 FILLER_44_170 ();
 sg13g2_fill_1 FILLER_44_235 ();
 sg13g2_fill_1 FILLER_44_249 ();
 sg13g2_decap_8 FILLER_44_293 ();
 sg13g2_fill_2 FILLER_44_300 ();
 sg13g2_fill_2 FILLER_44_310 ();
 sg13g2_fill_1 FILLER_44_332 ();
 sg13g2_fill_1 FILLER_44_390 ();
 sg13g2_decap_8 FILLER_44_401 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_fill_1 FILLER_45_28 ();
 sg13g2_fill_1 FILLER_45_72 ();
 sg13g2_fill_1 FILLER_45_125 ();
 sg13g2_fill_2 FILLER_45_161 ();
 sg13g2_fill_1 FILLER_45_163 ();
 sg13g2_decap_4 FILLER_45_203 ();
 sg13g2_fill_2 FILLER_45_207 ();
 sg13g2_fill_1 FILLER_45_218 ();
 sg13g2_fill_2 FILLER_45_243 ();
 sg13g2_fill_1 FILLER_45_245 ();
 sg13g2_fill_2 FILLER_45_251 ();
 sg13g2_fill_2 FILLER_45_258 ();
 sg13g2_fill_1 FILLER_45_301 ();
 sg13g2_fill_1 FILLER_45_322 ();
 sg13g2_fill_2 FILLER_45_340 ();
 sg13g2_fill_1 FILLER_45_342 ();
 sg13g2_fill_1 FILLER_45_356 ();
 sg13g2_fill_2 FILLER_45_383 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_4 FILLER_46_28 ();
 sg13g2_fill_1 FILLER_46_32 ();
 sg13g2_fill_1 FILLER_46_59 ();
 sg13g2_fill_2 FILLER_46_73 ();
 sg13g2_fill_2 FILLER_46_128 ();
 sg13g2_fill_2 FILLER_46_161 ();
 sg13g2_decap_8 FILLER_46_194 ();
 sg13g2_decap_8 FILLER_46_201 ();
 sg13g2_decap_8 FILLER_46_208 ();
 sg13g2_fill_1 FILLER_46_215 ();
 sg13g2_fill_1 FILLER_46_241 ();
 sg13g2_decap_4 FILLER_46_256 ();
 sg13g2_fill_2 FILLER_46_260 ();
 sg13g2_fill_1 FILLER_46_299 ();
 sg13g2_fill_1 FILLER_46_363 ();
 sg13g2_fill_2 FILLER_46_372 ();
 sg13g2_fill_1 FILLER_46_374 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_4 FILLER_47_35 ();
 sg13g2_fill_1 FILLER_47_53 ();
 sg13g2_fill_2 FILLER_47_80 ();
 sg13g2_fill_1 FILLER_47_100 ();
 sg13g2_fill_1 FILLER_47_137 ();
 sg13g2_fill_1 FILLER_47_153 ();
 sg13g2_decap_8 FILLER_47_185 ();
 sg13g2_decap_4 FILLER_47_200 ();
 sg13g2_decap_4 FILLER_47_207 ();
 sg13g2_fill_1 FILLER_47_211 ();
 sg13g2_fill_1 FILLER_47_221 ();
 sg13g2_fill_2 FILLER_47_239 ();
 sg13g2_fill_1 FILLER_47_241 ();
 sg13g2_decap_8 FILLER_47_263 ();
 sg13g2_decap_4 FILLER_47_270 ();
 sg13g2_fill_1 FILLER_47_274 ();
 sg13g2_fill_1 FILLER_47_292 ();
 sg13g2_fill_2 FILLER_47_298 ();
 sg13g2_fill_1 FILLER_47_300 ();
 sg13g2_fill_1 FILLER_47_321 ();
 sg13g2_fill_1 FILLER_47_339 ();
 sg13g2_fill_2 FILLER_47_344 ();
 sg13g2_fill_1 FILLER_47_357 ();
 sg13g2_fill_1 FILLER_47_363 ();
 sg13g2_fill_2 FILLER_47_377 ();
 sg13g2_fill_1 FILLER_47_379 ();
 sg13g2_fill_1 FILLER_47_403 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_fill_2 FILLER_48_92 ();
 sg13g2_fill_2 FILLER_48_163 ();
 sg13g2_fill_1 FILLER_48_231 ();
 sg13g2_decap_8 FILLER_48_273 ();
 sg13g2_decap_4 FILLER_48_280 ();
 sg13g2_fill_1 FILLER_48_284 ();
 sg13g2_decap_8 FILLER_48_298 ();
 sg13g2_decap_4 FILLER_48_305 ();
 sg13g2_fill_2 FILLER_48_309 ();
 sg13g2_fill_2 FILLER_48_316 ();
 sg13g2_fill_2 FILLER_48_330 ();
 sg13g2_fill_1 FILLER_48_332 ();
 sg13g2_fill_1 FILLER_48_341 ();
 sg13g2_decap_8 FILLER_48_360 ();
 sg13g2_fill_2 FILLER_48_367 ();
 sg13g2_decap_4 FILLER_48_373 ();
 sg13g2_fill_2 FILLER_48_381 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_4 FILLER_49_42 ();
 sg13g2_fill_1 FILLER_49_46 ();
 sg13g2_fill_1 FILLER_49_77 ();
 sg13g2_fill_1 FILLER_49_102 ();
 sg13g2_fill_2 FILLER_49_130 ();
 sg13g2_decap_4 FILLER_49_191 ();
 sg13g2_fill_2 FILLER_49_195 ();
 sg13g2_fill_1 FILLER_49_226 ();
 sg13g2_fill_2 FILLER_49_267 ();
 sg13g2_decap_8 FILLER_49_300 ();
 sg13g2_decap_8 FILLER_49_307 ();
 sg13g2_fill_2 FILLER_49_314 ();
 sg13g2_decap_8 FILLER_49_334 ();
 sg13g2_decap_4 FILLER_49_341 ();
 sg13g2_fill_1 FILLER_49_345 ();
 sg13g2_decap_8 FILLER_49_350 ();
 sg13g2_decap_4 FILLER_49_357 ();
 sg13g2_fill_2 FILLER_49_361 ();
 sg13g2_decap_8 FILLER_49_367 ();
 sg13g2_fill_1 FILLER_49_374 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_4 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_43 ();
 sg13g2_decap_8 FILLER_50_50 ();
 sg13g2_fill_2 FILLER_50_161 ();
 sg13g2_decap_8 FILLER_50_184 ();
 sg13g2_decap_8 FILLER_50_191 ();
 sg13g2_fill_2 FILLER_50_216 ();
 sg13g2_fill_2 FILLER_50_249 ();
 sg13g2_fill_1 FILLER_50_251 ();
 sg13g2_fill_2 FILLER_50_261 ();
 sg13g2_fill_1 FILLER_50_263 ();
 sg13g2_fill_2 FILLER_50_295 ();
 sg13g2_fill_1 FILLER_50_325 ();
 sg13g2_decap_4 FILLER_50_341 ();
 sg13g2_fill_1 FILLER_50_363 ();
 sg13g2_decap_4 FILLER_50_380 ();
 sg13g2_fill_2 FILLER_50_406 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_fill_1 FILLER_51_54 ();
 sg13g2_fill_1 FILLER_51_95 ();
 sg13g2_fill_2 FILLER_51_106 ();
 sg13g2_fill_2 FILLER_51_174 ();
 sg13g2_fill_2 FILLER_51_218 ();
 sg13g2_fill_2 FILLER_51_241 ();
 sg13g2_fill_1 FILLER_51_295 ();
 sg13g2_fill_2 FILLER_51_361 ();
 sg13g2_decap_4 FILLER_51_392 ();
 sg13g2_decap_8 FILLER_51_400 ();
 sg13g2_fill_2 FILLER_51_407 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_4 FILLER_52_14 ();
 sg13g2_fill_2 FILLER_52_18 ();
 sg13g2_fill_2 FILLER_52_43 ();
 sg13g2_fill_2 FILLER_52_77 ();
 sg13g2_fill_2 FILLER_52_118 ();
 sg13g2_fill_1 FILLER_52_174 ();
 sg13g2_fill_2 FILLER_52_189 ();
 sg13g2_fill_1 FILLER_52_237 ();
 sg13g2_fill_1 FILLER_52_243 ();
 sg13g2_fill_1 FILLER_52_254 ();
 sg13g2_fill_2 FILLER_52_263 ();
 sg13g2_fill_1 FILLER_52_308 ();
 sg13g2_fill_1 FILLER_52_344 ();
 sg13g2_fill_1 FILLER_52_350 ();
 sg13g2_decap_8 FILLER_52_377 ();
 sg13g2_fill_2 FILLER_52_384 ();
 sg13g2_fill_1 FILLER_52_386 ();
 sg13g2_decap_8 FILLER_52_394 ();
 sg13g2_fill_2 FILLER_52_401 ();
 sg13g2_fill_2 FILLER_52_407 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_fill_1 FILLER_53_21 ();
 sg13g2_fill_2 FILLER_53_135 ();
 sg13g2_fill_1 FILLER_53_137 ();
 sg13g2_fill_1 FILLER_53_160 ();
 sg13g2_fill_1 FILLER_53_205 ();
 sg13g2_fill_2 FILLER_53_254 ();
 sg13g2_decap_4 FILLER_53_265 ();
 sg13g2_fill_2 FILLER_53_269 ();
 sg13g2_decap_4 FILLER_53_289 ();
 sg13g2_decap_8 FILLER_53_297 ();
 sg13g2_decap_8 FILLER_53_304 ();
 sg13g2_decap_4 FILLER_53_311 ();
 sg13g2_decap_4 FILLER_53_341 ();
 sg13g2_decap_8 FILLER_53_363 ();
 sg13g2_fill_1 FILLER_53_370 ();
 sg13g2_fill_2 FILLER_53_375 ();
 sg13g2_fill_1 FILLER_53_377 ();
 sg13g2_fill_1 FILLER_53_408 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_4 FILLER_54_7 ();
 sg13g2_fill_1 FILLER_54_65 ();
 sg13g2_fill_1 FILLER_54_92 ();
 sg13g2_fill_2 FILLER_54_110 ();
 sg13g2_fill_2 FILLER_54_156 ();
 sg13g2_fill_1 FILLER_54_185 ();
 sg13g2_fill_1 FILLER_54_230 ();
 sg13g2_decap_4 FILLER_54_266 ();
 sg13g2_fill_2 FILLER_54_275 ();
 sg13g2_fill_1 FILLER_54_277 ();
 sg13g2_decap_4 FILLER_54_283 ();
 sg13g2_fill_2 FILLER_54_291 ();
 sg13g2_fill_1 FILLER_54_293 ();
 sg13g2_decap_8 FILLER_54_299 ();
 sg13g2_decap_4 FILLER_54_306 ();
 sg13g2_fill_2 FILLER_54_321 ();
 sg13g2_fill_1 FILLER_54_328 ();
 sg13g2_decap_4 FILLER_54_333 ();
 sg13g2_fill_1 FILLER_54_337 ();
 sg13g2_fill_1 FILLER_54_351 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_fill_2 FILLER_55_14 ();
 sg13g2_decap_4 FILLER_55_88 ();
 sg13g2_fill_1 FILLER_55_92 ();
 sg13g2_decap_8 FILLER_55_114 ();
 sg13g2_fill_2 FILLER_55_121 ();
 sg13g2_fill_2 FILLER_55_132 ();
 sg13g2_fill_2 FILLER_55_178 ();
 sg13g2_fill_2 FILLER_55_308 ();
 sg13g2_fill_1 FILLER_55_310 ();
 sg13g2_fill_2 FILLER_55_336 ();
 sg13g2_fill_1 FILLER_55_362 ();
 sg13g2_fill_2 FILLER_55_377 ();
 sg13g2_fill_2 FILLER_55_407 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_fill_2 FILLER_56_21 ();
 sg13g2_fill_1 FILLER_56_23 ();
 sg13g2_fill_1 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_85 ();
 sg13g2_fill_2 FILLER_56_92 ();
 sg13g2_fill_1 FILLER_56_94 ();
 sg13g2_decap_4 FILLER_56_126 ();
 sg13g2_fill_1 FILLER_56_135 ();
 sg13g2_fill_2 FILLER_56_150 ();
 sg13g2_fill_1 FILLER_56_161 ();
 sg13g2_fill_1 FILLER_56_262 ();
 sg13g2_fill_1 FILLER_56_276 ();
 sg13g2_fill_2 FILLER_56_286 ();
 sg13g2_fill_1 FILLER_56_288 ();
 sg13g2_fill_1 FILLER_56_344 ();
 sg13g2_decap_8 FILLER_56_370 ();
 sg13g2_fill_2 FILLER_56_406 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_fill_1 FILLER_57_67 ();
 sg13g2_fill_1 FILLER_57_72 ();
 sg13g2_fill_1 FILLER_57_87 ();
 sg13g2_fill_2 FILLER_57_101 ();
 sg13g2_fill_1 FILLER_57_103 ();
 sg13g2_fill_1 FILLER_57_195 ();
 sg13g2_fill_1 FILLER_57_322 ();
 sg13g2_decap_4 FILLER_57_327 ();
 sg13g2_fill_2 FILLER_57_331 ();
 sg13g2_decap_8 FILLER_57_342 ();
 sg13g2_decap_4 FILLER_57_349 ();
 sg13g2_fill_2 FILLER_57_378 ();
 sg13g2_fill_2 FILLER_57_388 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_fill_1 FILLER_58_7 ();
 sg13g2_fill_2 FILLER_58_34 ();
 sg13g2_fill_1 FILLER_58_50 ();
 sg13g2_decap_4 FILLER_58_66 ();
 sg13g2_fill_1 FILLER_58_70 ();
 sg13g2_fill_1 FILLER_58_109 ();
 sg13g2_fill_1 FILLER_58_123 ();
 sg13g2_fill_2 FILLER_58_133 ();
 sg13g2_fill_1 FILLER_58_135 ();
 sg13g2_fill_1 FILLER_58_188 ();
 sg13g2_fill_2 FILLER_58_216 ();
 sg13g2_decap_8 FILLER_58_229 ();
 sg13g2_decap_4 FILLER_58_236 ();
 sg13g2_decap_4 FILLER_58_243 ();
 sg13g2_fill_2 FILLER_58_247 ();
 sg13g2_fill_1 FILLER_58_271 ();
 sg13g2_fill_1 FILLER_58_284 ();
 sg13g2_decap_8 FILLER_58_311 ();
 sg13g2_fill_1 FILLER_58_318 ();
 sg13g2_decap_8 FILLER_58_324 ();
 sg13g2_fill_2 FILLER_58_331 ();
 sg13g2_fill_1 FILLER_58_333 ();
 sg13g2_fill_2 FILLER_58_357 ();
 sg13g2_fill_1 FILLER_58_359 ();
 sg13g2_decap_4 FILLER_58_379 ();
 sg13g2_fill_1 FILLER_58_383 ();
 sg13g2_fill_2 FILLER_58_392 ();
 sg13g2_fill_1 FILLER_58_394 ();
 sg13g2_decap_4 FILLER_59_0 ();
 sg13g2_fill_1 FILLER_59_65 ();
 sg13g2_fill_1 FILLER_59_92 ();
 sg13g2_fill_2 FILLER_59_112 ();
 sg13g2_fill_1 FILLER_59_114 ();
 sg13g2_fill_2 FILLER_59_120 ();
 sg13g2_fill_1 FILLER_59_122 ();
 sg13g2_decap_4 FILLER_59_128 ();
 sg13g2_fill_2 FILLER_59_132 ();
 sg13g2_fill_2 FILLER_59_139 ();
 sg13g2_fill_1 FILLER_59_141 ();
 sg13g2_fill_1 FILLER_59_160 ();
 sg13g2_fill_2 FILLER_59_195 ();
 sg13g2_fill_2 FILLER_59_226 ();
 sg13g2_fill_1 FILLER_59_228 ();
 sg13g2_fill_1 FILLER_59_255 ();
 sg13g2_fill_2 FILLER_59_261 ();
 sg13g2_fill_1 FILLER_59_263 ();
 sg13g2_fill_2 FILLER_59_293 ();
 sg13g2_decap_4 FILLER_59_298 ();
 sg13g2_fill_2 FILLER_59_302 ();
 sg13g2_fill_1 FILLER_59_313 ();
 sg13g2_fill_1 FILLER_59_319 ();
 sg13g2_fill_2 FILLER_59_327 ();
 sg13g2_fill_1 FILLER_59_329 ();
 sg13g2_fill_2 FILLER_59_356 ();
 sg13g2_fill_1 FILLER_59_358 ();
 sg13g2_fill_2 FILLER_59_380 ();
 sg13g2_fill_2 FILLER_59_407 ();
 sg13g2_fill_1 FILLER_60_73 ();
 sg13g2_fill_2 FILLER_60_83 ();
 sg13g2_fill_1 FILLER_60_103 ();
 sg13g2_fill_2 FILLER_60_120 ();
 sg13g2_fill_1 FILLER_60_122 ();
 sg13g2_fill_2 FILLER_60_128 ();
 sg13g2_fill_2 FILLER_60_135 ();
 sg13g2_fill_2 FILLER_60_142 ();
 sg13g2_fill_2 FILLER_60_153 ();
 sg13g2_fill_2 FILLER_60_195 ();
 sg13g2_fill_2 FILLER_60_228 ();
 sg13g2_decap_8 FILLER_60_253 ();
 sg13g2_fill_2 FILLER_60_260 ();
 sg13g2_fill_2 FILLER_60_268 ();
 sg13g2_fill_1 FILLER_60_270 ();
 sg13g2_fill_2 FILLER_60_293 ();
 sg13g2_fill_1 FILLER_60_295 ();
 sg13g2_decap_4 FILLER_60_300 ();
 sg13g2_fill_1 FILLER_60_304 ();
 sg13g2_fill_1 FILLER_60_333 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_7 ();
 sg13g2_fill_2 FILLER_61_55 ();
 sg13g2_fill_1 FILLER_61_71 ();
 sg13g2_fill_2 FILLER_61_120 ();
 sg13g2_fill_1 FILLER_61_148 ();
 sg13g2_fill_1 FILLER_61_184 ();
 sg13g2_fill_2 FILLER_61_221 ();
 sg13g2_fill_2 FILLER_61_280 ();
 sg13g2_fill_1 FILLER_61_282 ();
 sg13g2_fill_2 FILLER_61_309 ();
 sg13g2_decap_8 FILLER_61_332 ();
 sg13g2_decap_4 FILLER_61_339 ();
 sg13g2_fill_1 FILLER_61_343 ();
 sg13g2_decap_4 FILLER_61_372 ();
 sg13g2_fill_1 FILLER_61_376 ();
 sg13g2_decap_4 FILLER_62_0 ();
 sg13g2_fill_2 FILLER_62_4 ();
 sg13g2_fill_1 FILLER_62_63 ();
 sg13g2_fill_1 FILLER_62_89 ();
 sg13g2_fill_2 FILLER_62_124 ();
 sg13g2_fill_2 FILLER_62_131 ();
 sg13g2_fill_2 FILLER_62_141 ();
 sg13g2_fill_1 FILLER_62_143 ();
 sg13g2_fill_1 FILLER_62_149 ();
 sg13g2_fill_1 FILLER_62_167 ();
 sg13g2_fill_1 FILLER_62_199 ();
 sg13g2_fill_1 FILLER_62_214 ();
 sg13g2_fill_1 FILLER_62_243 ();
 sg13g2_fill_2 FILLER_62_330 ();
 sg13g2_decap_8 FILLER_62_350 ();
 sg13g2_decap_4 FILLER_62_357 ();
 sg13g2_decap_8 FILLER_62_366 ();
 sg13g2_decap_8 FILLER_62_373 ();
 sg13g2_fill_2 FILLER_62_380 ();
 sg13g2_fill_1 FILLER_62_382 ();
 sg13g2_fill_1 FILLER_62_387 ();
 sg13g2_decap_4 FILLER_62_392 ();
 sg13g2_fill_1 FILLER_62_396 ();
 sg13g2_fill_2 FILLER_62_406 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_4 FILLER_63_7 ();
 sg13g2_fill_1 FILLER_63_11 ();
 sg13g2_fill_1 FILLER_63_131 ();
 sg13g2_fill_2 FILLER_63_163 ();
 sg13g2_fill_2 FILLER_63_182 ();
 sg13g2_fill_2 FILLER_63_193 ();
 sg13g2_fill_2 FILLER_63_200 ();
 sg13g2_fill_2 FILLER_63_331 ();
 sg13g2_fill_1 FILLER_63_333 ();
 sg13g2_fill_1 FILLER_63_347 ();
 sg13g2_decap_4 FILLER_63_362 ();
 sg13g2_fill_2 FILLER_63_366 ();
 sg13g2_fill_1 FILLER_63_382 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_fill_1 FILLER_64_7 ();
 sg13g2_fill_1 FILLER_64_34 ();
 sg13g2_fill_2 FILLER_64_88 ();
 sg13g2_fill_1 FILLER_64_129 ();
 sg13g2_fill_2 FILLER_64_135 ();
 sg13g2_fill_1 FILLER_64_219 ();
 sg13g2_fill_2 FILLER_64_243 ();
 sg13g2_fill_2 FILLER_64_312 ();
 sg13g2_fill_1 FILLER_64_314 ();
 sg13g2_fill_2 FILLER_64_372 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_fill_2 FILLER_65_52 ();
 sg13g2_fill_1 FILLER_65_54 ();
 sg13g2_fill_1 FILLER_65_81 ();
 sg13g2_fill_2 FILLER_65_90 ();
 sg13g2_fill_1 FILLER_65_170 ();
 sg13g2_fill_2 FILLER_65_209 ();
 sg13g2_fill_1 FILLER_65_229 ();
 sg13g2_fill_2 FILLER_65_235 ();
 sg13g2_fill_2 FILLER_65_241 ();
 sg13g2_decap_8 FILLER_65_337 ();
 sg13g2_decap_8 FILLER_65_344 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_fill_2 FILLER_66_7 ();
 sg13g2_fill_1 FILLER_66_75 ();
 sg13g2_fill_1 FILLER_66_98 ();
 sg13g2_fill_2 FILLER_66_108 ();
 sg13g2_fill_1 FILLER_66_110 ();
 sg13g2_fill_1 FILLER_66_115 ();
 sg13g2_fill_2 FILLER_66_124 ();
 sg13g2_fill_1 FILLER_66_150 ();
 sg13g2_fill_1 FILLER_66_212 ();
 sg13g2_fill_2 FILLER_66_362 ();
 sg13g2_fill_2 FILLER_66_398 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_4 FILLER_67_14 ();
 sg13g2_fill_2 FILLER_67_18 ();
 sg13g2_fill_2 FILLER_67_60 ();
 sg13g2_fill_1 FILLER_67_62 ();
 sg13g2_fill_1 FILLER_67_81 ();
 sg13g2_decap_4 FILLER_67_102 ();
 sg13g2_fill_1 FILLER_67_106 ();
 sg13g2_fill_2 FILLER_67_137 ();
 sg13g2_fill_1 FILLER_67_139 ();
 sg13g2_fill_2 FILLER_67_149 ();
 sg13g2_fill_2 FILLER_67_184 ();
 sg13g2_fill_2 FILLER_67_195 ();
 sg13g2_fill_1 FILLER_67_281 ();
 sg13g2_fill_2 FILLER_67_331 ();
 sg13g2_fill_1 FILLER_67_333 ();
 sg13g2_decap_8 FILLER_67_338 ();
 sg13g2_decap_8 FILLER_67_345 ();
 sg13g2_fill_1 FILLER_67_352 ();
 sg13g2_fill_2 FILLER_67_366 ();
 sg13g2_fill_1 FILLER_67_368 ();
 sg13g2_fill_1 FILLER_67_388 ();
 sg13g2_fill_2 FILLER_67_406 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_fill_2 FILLER_68_21 ();
 sg13g2_fill_2 FILLER_68_102 ();
 sg13g2_fill_1 FILLER_68_104 ();
 sg13g2_fill_1 FILLER_68_113 ();
 sg13g2_fill_1 FILLER_68_237 ();
 sg13g2_fill_2 FILLER_68_299 ();
 sg13g2_decap_4 FILLER_68_321 ();
 sg13g2_fill_1 FILLER_68_381 ();
 sg13g2_decap_4 FILLER_68_390 ();
 sg13g2_fill_2 FILLER_68_406 ();
 sg13g2_fill_1 FILLER_68_408 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_fill_2 FILLER_69_14 ();
 sg13g2_fill_1 FILLER_69_74 ();
 sg13g2_fill_1 FILLER_69_103 ();
 sg13g2_fill_2 FILLER_69_146 ();
 sg13g2_fill_1 FILLER_69_304 ();
 sg13g2_fill_2 FILLER_69_335 ();
 sg13g2_fill_1 FILLER_69_347 ();
 sg13g2_fill_1 FILLER_69_367 ();
 sg13g2_fill_2 FILLER_69_380 ();
 sg13g2_fill_1 FILLER_69_382 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_4 FILLER_70_14 ();
 sg13g2_fill_2 FILLER_70_88 ();
 sg13g2_fill_2 FILLER_70_95 ();
 sg13g2_fill_1 FILLER_70_97 ();
 sg13g2_decap_8 FILLER_70_129 ();
 sg13g2_fill_2 FILLER_70_136 ();
 sg13g2_fill_1 FILLER_70_142 ();
 sg13g2_decap_8 FILLER_70_148 ();
 sg13g2_fill_1 FILLER_70_155 ();
 sg13g2_fill_2 FILLER_70_186 ();
 sg13g2_fill_1 FILLER_70_188 ();
 sg13g2_fill_2 FILLER_70_211 ();
 sg13g2_decap_4 FILLER_70_239 ();
 sg13g2_decap_8 FILLER_70_249 ();
 sg13g2_fill_1 FILLER_70_256 ();
 sg13g2_fill_1 FILLER_70_269 ();
 sg13g2_fill_2 FILLER_70_340 ();
 sg13g2_fill_1 FILLER_70_384 ();
 sg13g2_fill_2 FILLER_70_402 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_fill_2 FILLER_71_7 ();
 sg13g2_fill_1 FILLER_71_9 ();
 sg13g2_fill_1 FILLER_71_42 ();
 sg13g2_fill_1 FILLER_71_52 ();
 sg13g2_fill_1 FILLER_71_100 ();
 sg13g2_fill_2 FILLER_71_113 ();
 sg13g2_fill_1 FILLER_71_115 ();
 sg13g2_fill_2 FILLER_71_135 ();
 sg13g2_fill_1 FILLER_71_137 ();
 sg13g2_decap_8 FILLER_71_143 ();
 sg13g2_decap_8 FILLER_71_150 ();
 sg13g2_decap_8 FILLER_71_157 ();
 sg13g2_decap_4 FILLER_71_164 ();
 sg13g2_fill_2 FILLER_71_168 ();
 sg13g2_decap_4 FILLER_71_174 ();
 sg13g2_fill_2 FILLER_71_178 ();
 sg13g2_fill_2 FILLER_71_184 ();
 sg13g2_decap_4 FILLER_71_190 ();
 sg13g2_fill_1 FILLER_71_194 ();
 sg13g2_decap_8 FILLER_71_207 ();
 sg13g2_fill_1 FILLER_71_214 ();
 sg13g2_decap_4 FILLER_71_266 ();
 sg13g2_fill_2 FILLER_71_353 ();
 sg13g2_fill_2 FILLER_71_376 ();
 sg13g2_fill_1 FILLER_71_383 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_fill_2 FILLER_72_14 ();
 sg13g2_fill_2 FILLER_72_48 ();
 sg13g2_fill_1 FILLER_72_76 ();
 sg13g2_fill_2 FILLER_72_92 ();
 sg13g2_fill_1 FILLER_72_94 ();
 sg13g2_fill_2 FILLER_72_105 ();
 sg13g2_fill_1 FILLER_72_112 ();
 sg13g2_fill_2 FILLER_72_123 ();
 sg13g2_fill_1 FILLER_72_189 ();
 sg13g2_decap_8 FILLER_72_199 ();
 sg13g2_decap_8 FILLER_72_206 ();
 sg13g2_fill_2 FILLER_72_213 ();
 sg13g2_fill_1 FILLER_72_215 ();
 sg13g2_fill_1 FILLER_72_237 ();
 sg13g2_fill_1 FILLER_72_264 ();
 sg13g2_fill_2 FILLER_72_291 ();
 sg13g2_decap_4 FILLER_72_297 ();
 sg13g2_fill_2 FILLER_72_301 ();
 sg13g2_fill_2 FILLER_72_321 ();
 sg13g2_fill_2 FILLER_72_328 ();
 sg13g2_fill_1 FILLER_72_330 ();
 sg13g2_decap_8 FILLER_72_336 ();
 sg13g2_fill_2 FILLER_72_343 ();
 sg13g2_fill_1 FILLER_72_357 ();
 sg13g2_fill_1 FILLER_72_370 ();
 sg13g2_fill_2 FILLER_72_393 ();
 sg13g2_fill_1 FILLER_72_395 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_fill_2 FILLER_73_21 ();
 sg13g2_fill_2 FILLER_73_64 ();
 sg13g2_fill_1 FILLER_73_105 ();
 sg13g2_fill_2 FILLER_73_141 ();
 sg13g2_fill_2 FILLER_73_174 ();
 sg13g2_fill_2 FILLER_73_211 ();
 sg13g2_fill_2 FILLER_73_220 ();
 sg13g2_fill_2 FILLER_73_244 ();
 sg13g2_fill_1 FILLER_73_259 ();
 sg13g2_decap_4 FILLER_73_283 ();
 sg13g2_fill_2 FILLER_73_326 ();
 sg13g2_fill_1 FILLER_73_328 ();
 sg13g2_decap_4 FILLER_73_338 ();
 sg13g2_decap_8 FILLER_73_347 ();
 sg13g2_fill_2 FILLER_73_354 ();
 sg13g2_decap_8 FILLER_73_374 ();
 sg13g2_fill_2 FILLER_73_381 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_4 FILLER_74_21 ();
 sg13g2_fill_1 FILLER_74_51 ();
 sg13g2_fill_1 FILLER_74_61 ();
 sg13g2_fill_2 FILLER_74_87 ();
 sg13g2_fill_1 FILLER_74_89 ();
 sg13g2_fill_2 FILLER_74_100 ();
 sg13g2_fill_1 FILLER_74_102 ();
 sg13g2_fill_1 FILLER_74_129 ();
 sg13g2_fill_2 FILLER_74_144 ();
 sg13g2_fill_1 FILLER_74_146 ();
 sg13g2_fill_2 FILLER_74_225 ();
 sg13g2_decap_4 FILLER_74_299 ();
 sg13g2_fill_1 FILLER_74_303 ();
 sg13g2_decap_8 FILLER_74_356 ();
 sg13g2_decap_8 FILLER_74_363 ();
 sg13g2_fill_2 FILLER_74_370 ();
 sg13g2_fill_2 FILLER_74_407 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_4 FILLER_75_28 ();
 sg13g2_fill_1 FILLER_75_48 ();
 sg13g2_fill_1 FILLER_75_84 ();
 sg13g2_fill_2 FILLER_75_135 ();
 sg13g2_fill_1 FILLER_75_147 ();
 sg13g2_decap_4 FILLER_75_153 ();
 sg13g2_fill_2 FILLER_75_157 ();
 sg13g2_fill_1 FILLER_75_167 ();
 sg13g2_fill_1 FILLER_75_203 ();
 sg13g2_fill_2 FILLER_75_296 ();
 sg13g2_fill_1 FILLER_75_328 ();
 sg13g2_fill_2 FILLER_75_338 ();
 sg13g2_fill_1 FILLER_75_340 ();
 sg13g2_fill_1 FILLER_75_349 ();
 sg13g2_fill_2 FILLER_75_363 ();
 sg13g2_decap_4 FILLER_75_378 ();
 sg13g2_fill_1 FILLER_75_382 ();
 sg13g2_decap_8 FILLER_75_396 ();
 sg13g2_decap_4 FILLER_75_403 ();
 sg13g2_fill_2 FILLER_75_407 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_4 FILLER_76_21 ();
 sg13g2_fill_2 FILLER_76_47 ();
 sg13g2_fill_2 FILLER_76_58 ();
 sg13g2_fill_1 FILLER_76_60 ();
 sg13g2_fill_2 FILLER_76_69 ();
 sg13g2_fill_2 FILLER_76_105 ();
 sg13g2_fill_2 FILLER_76_111 ();
 sg13g2_fill_1 FILLER_76_113 ();
 sg13g2_decap_4 FILLER_76_133 ();
 sg13g2_decap_4 FILLER_76_147 ();
 sg13g2_fill_2 FILLER_76_188 ();
 sg13g2_fill_1 FILLER_76_212 ();
 sg13g2_fill_1 FILLER_76_218 ();
 sg13g2_fill_1 FILLER_76_228 ();
 sg13g2_fill_1 FILLER_76_287 ();
 sg13g2_decap_4 FILLER_76_304 ();
 sg13g2_fill_1 FILLER_76_308 ();
 sg13g2_fill_2 FILLER_76_317 ();
 sg13g2_fill_1 FILLER_76_327 ();
 sg13g2_fill_1 FILLER_76_333 ();
 sg13g2_fill_2 FILLER_76_337 ();
 sg13g2_fill_1 FILLER_76_344 ();
 sg13g2_decap_8 FILLER_76_349 ();
 sg13g2_fill_1 FILLER_76_356 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_fill_2 FILLER_77_21 ();
 sg13g2_fill_1 FILLER_77_53 ();
 sg13g2_fill_2 FILLER_77_122 ();
 sg13g2_fill_1 FILLER_77_227 ();
 sg13g2_fill_2 FILLER_77_238 ();
 sg13g2_fill_1 FILLER_77_266 ();
 sg13g2_decap_8 FILLER_77_399 ();
 sg13g2_fill_2 FILLER_77_406 ();
 sg13g2_fill_1 FILLER_77_408 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_fill_2 FILLER_78_124 ();
 sg13g2_fill_1 FILLER_78_126 ();
 sg13g2_fill_2 FILLER_78_185 ();
 sg13g2_fill_2 FILLER_78_240 ();
 sg13g2_fill_1 FILLER_78_251 ();
 sg13g2_fill_2 FILLER_78_261 ();
 sg13g2_fill_1 FILLER_78_315 ();
 sg13g2_fill_2 FILLER_78_342 ();
 sg13g2_fill_1 FILLER_78_376 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_fill_2 FILLER_79_35 ();
 sg13g2_fill_2 FILLER_79_45 ();
 sg13g2_fill_1 FILLER_79_47 ();
 sg13g2_decap_4 FILLER_79_57 ();
 sg13g2_fill_2 FILLER_79_61 ();
 sg13g2_decap_4 FILLER_79_100 ();
 sg13g2_fill_2 FILLER_79_104 ();
 sg13g2_fill_1 FILLER_79_137 ();
 sg13g2_fill_1 FILLER_79_190 ();
 sg13g2_fill_2 FILLER_79_221 ();
 sg13g2_fill_1 FILLER_79_275 ();
 sg13g2_fill_2 FILLER_79_295 ();
 sg13g2_fill_2 FILLER_79_349 ();
 sg13g2_fill_2 FILLER_79_363 ();
 sg13g2_decap_4 FILLER_79_405 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_fill_1 FILLER_80_76 ();
 sg13g2_fill_2 FILLER_80_94 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_fill_1 FILLER_80_216 ();
 sg13g2_fill_2 FILLER_80_272 ();
 sg13g2_fill_2 FILLER_80_350 ();
 sg13g2_fill_2 FILLER_80_373 ();
 sg13g2_fill_1 FILLER_80_375 ();
 sg13g2_decap_8 FILLER_80_402 ();
 assign uio_oe[0] = net9;
 assign uio_oe[1] = net10;
 assign uio_oe[2] = net11;
 assign uio_oe[3] = net12;
 assign uio_oe[4] = net13;
 assign uio_oe[5] = net14;
 assign uio_oe[6] = net15;
 assign uio_oe[7] = net16;
 assign uio_out[0] = net17;
 assign uio_out[1] = net18;
 assign uio_out[2] = net19;
 assign uio_out[3] = net20;
 assign uio_out[4] = net21;
 assign uio_out[5] = net22;
 assign uio_out[6] = net23;
 assign uio_out[7] = net24;
 assign uo_out[7] = net25;
endmodule
