module tt_um_kianV_rv32ima_uLinux_SoC (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire _14944_;
 wire _14945_;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14983_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire _14990_;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire _14994_;
 wire _14995_;
 wire _14996_;
 wire _14997_;
 wire _14998_;
 wire _14999_;
 wire _15000_;
 wire _15001_;
 wire _15002_;
 wire _15003_;
 wire _15004_;
 wire _15005_;
 wire _15006_;
 wire _15007_;
 wire _15008_;
 wire _15009_;
 wire _15010_;
 wire _15011_;
 wire _15012_;
 wire _15013_;
 wire _15014_;
 wire _15015_;
 wire _15016_;
 wire _15017_;
 wire _15018_;
 wire _15019_;
 wire _15020_;
 wire _15021_;
 wire _15022_;
 wire _15023_;
 wire _15024_;
 wire _15025_;
 wire _15026_;
 wire _15027_;
 wire _15028_;
 wire _15029_;
 wire _15030_;
 wire _15031_;
 wire _15032_;
 wire _15033_;
 wire _15034_;
 wire _15035_;
 wire _15036_;
 wire _15037_;
 wire _15038_;
 wire _15039_;
 wire _15040_;
 wire _15041_;
 wire _15042_;
 wire _15043_;
 wire _15044_;
 wire _15045_;
 wire _15046_;
 wire _15047_;
 wire _15048_;
 wire _15049_;
 wire _15050_;
 wire _15051_;
 wire _15052_;
 wire _15053_;
 wire _15054_;
 wire _15055_;
 wire _15056_;
 wire _15057_;
 wire _15058_;
 wire _15059_;
 wire _15060_;
 wire _15061_;
 wire _15062_;
 wire _15063_;
 wire _15064_;
 wire _15065_;
 wire _15066_;
 wire _15067_;
 wire _15068_;
 wire _15069_;
 wire _15070_;
 wire _15071_;
 wire _15072_;
 wire _15073_;
 wire _15074_;
 wire _15075_;
 wire _15076_;
 wire _15077_;
 wire _15078_;
 wire _15079_;
 wire _15080_;
 wire _15081_;
 wire _15082_;
 wire _15083_;
 wire _15084_;
 wire _15085_;
 wire _15086_;
 wire _15087_;
 wire _15088_;
 wire _15089_;
 wire _15090_;
 wire _15091_;
 wire _15092_;
 wire _15093_;
 wire _15094_;
 wire _15095_;
 wire _15096_;
 wire _15097_;
 wire _15098_;
 wire _15099_;
 wire _15100_;
 wire _15101_;
 wire _15102_;
 wire _15103_;
 wire _15104_;
 wire _15105_;
 wire _15106_;
 wire _15107_;
 wire _15108_;
 wire _15109_;
 wire _15110_;
 wire _15111_;
 wire _15112_;
 wire _15113_;
 wire _15114_;
 wire _15115_;
 wire _15116_;
 wire _15117_;
 wire _15118_;
 wire _15119_;
 wire _15120_;
 wire _15121_;
 wire _15122_;
 wire _15123_;
 wire _15124_;
 wire _15125_;
 wire _15126_;
 wire _15127_;
 wire _15128_;
 wire _15129_;
 wire _15130_;
 wire _15131_;
 wire _15132_;
 wire _15133_;
 wire _15134_;
 wire _15135_;
 wire _15136_;
 wire _15137_;
 wire _15138_;
 wire _15139_;
 wire _15140_;
 wire _15141_;
 wire _15142_;
 wire _15143_;
 wire _15144_;
 wire _15145_;
 wire _15146_;
 wire _15147_;
 wire _15148_;
 wire _15149_;
 wire _15150_;
 wire _15151_;
 wire _15152_;
 wire _15153_;
 wire _15154_;
 wire _15155_;
 wire _15156_;
 wire _15157_;
 wire _15158_;
 wire _15159_;
 wire _15160_;
 wire _15161_;
 wire _15162_;
 wire _15163_;
 wire _15164_;
 wire _15165_;
 wire _15166_;
 wire _15167_;
 wire _15168_;
 wire _15169_;
 wire _15170_;
 wire _15171_;
 wire _15172_;
 wire _15173_;
 wire _15174_;
 wire _15175_;
 wire _15176_;
 wire _15177_;
 wire _15178_;
 wire _15179_;
 wire _15180_;
 wire _15181_;
 wire _15182_;
 wire _15183_;
 wire _15184_;
 wire _15185_;
 wire _15186_;
 wire _15187_;
 wire _15188_;
 wire _15189_;
 wire _15190_;
 wire _15191_;
 wire _15192_;
 wire _15193_;
 wire _15194_;
 wire _15195_;
 wire _15196_;
 wire _15197_;
 wire _15198_;
 wire _15199_;
 wire _15200_;
 wire _15201_;
 wire _15202_;
 wire _15203_;
 wire _15204_;
 wire _15205_;
 wire _15206_;
 wire _15207_;
 wire _15208_;
 wire _15209_;
 wire _15210_;
 wire _15211_;
 wire _15212_;
 wire _15213_;
 wire _15214_;
 wire _15215_;
 wire _15216_;
 wire _15217_;
 wire _15218_;
 wire _15219_;
 wire _15220_;
 wire _15221_;
 wire _15222_;
 wire _15223_;
 wire _15224_;
 wire _15225_;
 wire _15226_;
 wire _15227_;
 wire _15228_;
 wire _15229_;
 wire _15230_;
 wire _15231_;
 wire _15232_;
 wire _15233_;
 wire _15234_;
 wire _15235_;
 wire _15236_;
 wire _15237_;
 wire _15238_;
 wire _15239_;
 wire _15240_;
 wire _15241_;
 wire _15242_;
 wire _15243_;
 wire _15244_;
 wire _15245_;
 wire _15246_;
 wire _15247_;
 wire _15248_;
 wire _15249_;
 wire _15250_;
 wire _15251_;
 wire _15252_;
 wire _15253_;
 wire _15254_;
 wire _15255_;
 wire _15256_;
 wire _15257_;
 wire _15258_;
 wire _15259_;
 wire _15260_;
 wire _15261_;
 wire _15262_;
 wire _15263_;
 wire _15264_;
 wire _15265_;
 wire _15266_;
 wire _15267_;
 wire _15268_;
 wire _15269_;
 wire _15270_;
 wire _15271_;
 wire _15272_;
 wire _15273_;
 wire _15274_;
 wire _15275_;
 wire _15276_;
 wire _15277_;
 wire _15278_;
 wire _15279_;
 wire _15280_;
 wire _15281_;
 wire _15282_;
 wire _15283_;
 wire _15284_;
 wire _15285_;
 wire _15286_;
 wire _15287_;
 wire _15288_;
 wire _15289_;
 wire _15290_;
 wire _15291_;
 wire _15292_;
 wire _15293_;
 wire _15294_;
 wire _15295_;
 wire _15296_;
 wire _15297_;
 wire _15298_;
 wire _15299_;
 wire _15300_;
 wire _15301_;
 wire _15302_;
 wire _15303_;
 wire _15304_;
 wire _15305_;
 wire _15306_;
 wire _15307_;
 wire _15308_;
 wire _15309_;
 wire _15310_;
 wire _15311_;
 wire _15312_;
 wire _15313_;
 wire _15314_;
 wire _15315_;
 wire _15316_;
 wire _15317_;
 wire _15318_;
 wire _15319_;
 wire _15320_;
 wire _15321_;
 wire _15322_;
 wire _15323_;
 wire _15324_;
 wire _15325_;
 wire _15326_;
 wire _15327_;
 wire _15328_;
 wire _15329_;
 wire _15330_;
 wire _15331_;
 wire _15332_;
 wire _15333_;
 wire _15334_;
 wire _15335_;
 wire _15336_;
 wire _15337_;
 wire _15338_;
 wire _15339_;
 wire _15340_;
 wire _15341_;
 wire _15342_;
 wire _15343_;
 wire _15344_;
 wire _15345_;
 wire _15346_;
 wire _15347_;
 wire _15348_;
 wire _15349_;
 wire _15350_;
 wire _15351_;
 wire _15352_;
 wire _15353_;
 wire _15354_;
 wire _15355_;
 wire _15356_;
 wire _15357_;
 wire _15358_;
 wire _15359_;
 wire _15360_;
 wire _15361_;
 wire _15362_;
 wire _15363_;
 wire _15364_;
 wire _15365_;
 wire _15366_;
 wire _15367_;
 wire _15368_;
 wire _15369_;
 wire _15370_;
 wire _15371_;
 wire _15372_;
 wire _15373_;
 wire _15374_;
 wire _15375_;
 wire _15376_;
 wire _15377_;
 wire _15378_;
 wire _15379_;
 wire _15380_;
 wire _15381_;
 wire _15382_;
 wire _15383_;
 wire _15384_;
 wire _15385_;
 wire _15386_;
 wire _15387_;
 wire _15388_;
 wire _15389_;
 wire _15390_;
 wire _15391_;
 wire _15392_;
 wire _15393_;
 wire _15394_;
 wire _15395_;
 wire _15396_;
 wire _15397_;
 wire _15398_;
 wire _15399_;
 wire _15400_;
 wire _15401_;
 wire _15402_;
 wire _15403_;
 wire _15404_;
 wire _15405_;
 wire _15406_;
 wire _15407_;
 wire _15408_;
 wire _15409_;
 wire _15410_;
 wire _15411_;
 wire _15412_;
 wire _15413_;
 wire _15414_;
 wire _15415_;
 wire _15416_;
 wire _15417_;
 wire _15418_;
 wire _15419_;
 wire _15420_;
 wire _15421_;
 wire _15422_;
 wire _15423_;
 wire _15424_;
 wire _15425_;
 wire _15426_;
 wire _15427_;
 wire _15428_;
 wire _15429_;
 wire _15430_;
 wire _15431_;
 wire _15432_;
 wire _15433_;
 wire _15434_;
 wire _15435_;
 wire _15436_;
 wire _15437_;
 wire _15438_;
 wire _15439_;
 wire _15440_;
 wire _15441_;
 wire _15442_;
 wire _15443_;
 wire _15444_;
 wire _15445_;
 wire _15446_;
 wire _15447_;
 wire _15448_;
 wire _15449_;
 wire _15450_;
 wire _15451_;
 wire _15452_;
 wire _15453_;
 wire _15454_;
 wire _15455_;
 wire _15456_;
 wire _15457_;
 wire _15458_;
 wire _15459_;
 wire _15460_;
 wire _15461_;
 wire _15462_;
 wire _15463_;
 wire _15464_;
 wire _15465_;
 wire _15466_;
 wire _15467_;
 wire _15468_;
 wire _15469_;
 wire _15470_;
 wire _15471_;
 wire _15472_;
 wire _15473_;
 wire _15474_;
 wire _15475_;
 wire _15476_;
 wire _15477_;
 wire _15478_;
 wire _15479_;
 wire _15480_;
 wire _15481_;
 wire _15482_;
 wire _15483_;
 wire _15484_;
 wire _15485_;
 wire _15486_;
 wire _15487_;
 wire _15488_;
 wire _15489_;
 wire _15490_;
 wire _15491_;
 wire _15492_;
 wire _15493_;
 wire _15494_;
 wire _15495_;
 wire _15496_;
 wire _15497_;
 wire _15498_;
 wire _15499_;
 wire _15500_;
 wire _15501_;
 wire _15502_;
 wire _15503_;
 wire _15504_;
 wire _15505_;
 wire _15506_;
 wire _15507_;
 wire _15508_;
 wire _15509_;
 wire _15510_;
 wire _15511_;
 wire _15512_;
 wire _15513_;
 wire _15514_;
 wire _15515_;
 wire _15516_;
 wire _15517_;
 wire _15518_;
 wire _15519_;
 wire _15520_;
 wire _15521_;
 wire _15522_;
 wire _15523_;
 wire _15524_;
 wire _15525_;
 wire _15526_;
 wire _15527_;
 wire _15528_;
 wire _15529_;
 wire _15530_;
 wire _15531_;
 wire _15532_;
 wire _15533_;
 wire _15534_;
 wire _15535_;
 wire _15536_;
 wire _15537_;
 wire _15538_;
 wire _15539_;
 wire _15540_;
 wire _15541_;
 wire _15542_;
 wire _15543_;
 wire _15544_;
 wire _15545_;
 wire _15546_;
 wire _15547_;
 wire _15548_;
 wire _15549_;
 wire _15550_;
 wire _15551_;
 wire _15552_;
 wire _15553_;
 wire _15554_;
 wire _15555_;
 wire _15556_;
 wire _15557_;
 wire _15558_;
 wire _15559_;
 wire _15560_;
 wire _15561_;
 wire _15562_;
 wire _15563_;
 wire _15564_;
 wire _15565_;
 wire _15566_;
 wire _15567_;
 wire _15568_;
 wire _15569_;
 wire _15570_;
 wire _15571_;
 wire _15572_;
 wire _15573_;
 wire _15574_;
 wire _15575_;
 wire _15576_;
 wire _15577_;
 wire _15578_;
 wire _15579_;
 wire _15580_;
 wire _15581_;
 wire _15582_;
 wire _15583_;
 wire _15584_;
 wire _15585_;
 wire _15586_;
 wire _15587_;
 wire _15588_;
 wire _15589_;
 wire _15590_;
 wire _15591_;
 wire _15592_;
 wire _15593_;
 wire _15594_;
 wire _15595_;
 wire _15596_;
 wire _15597_;
 wire _15598_;
 wire _15599_;
 wire _15600_;
 wire _15601_;
 wire _15602_;
 wire _15603_;
 wire _15604_;
 wire _15605_;
 wire _15606_;
 wire _15607_;
 wire _15608_;
 wire _15609_;
 wire _15610_;
 wire _15611_;
 wire _15612_;
 wire _15613_;
 wire _15614_;
 wire _15615_;
 wire _15616_;
 wire _15617_;
 wire _15618_;
 wire _15619_;
 wire _15620_;
 wire _15621_;
 wire _15622_;
 wire _15623_;
 wire _15624_;
 wire _15625_;
 wire _15626_;
 wire _15627_;
 wire _15628_;
 wire _15629_;
 wire _15630_;
 wire _15631_;
 wire _15632_;
 wire _15633_;
 wire _15634_;
 wire _15635_;
 wire _15636_;
 wire _15637_;
 wire _15638_;
 wire _15639_;
 wire _15640_;
 wire _15641_;
 wire _15642_;
 wire _15643_;
 wire _15644_;
 wire _15645_;
 wire _15646_;
 wire _15647_;
 wire _15648_;
 wire _15649_;
 wire _15650_;
 wire _15651_;
 wire _15652_;
 wire _15653_;
 wire _15654_;
 wire _15655_;
 wire _15656_;
 wire _15657_;
 wire _15658_;
 wire _15659_;
 wire _15660_;
 wire _15661_;
 wire _15662_;
 wire _15663_;
 wire _15664_;
 wire _15665_;
 wire _15666_;
 wire _15667_;
 wire _15668_;
 wire _15669_;
 wire _15670_;
 wire _15671_;
 wire _15672_;
 wire _15673_;
 wire _15674_;
 wire _15675_;
 wire _15676_;
 wire _15677_;
 wire _15678_;
 wire _15679_;
 wire _15680_;
 wire _15681_;
 wire _15682_;
 wire _15683_;
 wire _15684_;
 wire _15685_;
 wire _15686_;
 wire _15687_;
 wire _15688_;
 wire _15689_;
 wire _15690_;
 wire _15691_;
 wire _15692_;
 wire _15693_;
 wire _15694_;
 wire _15695_;
 wire _15696_;
 wire _15697_;
 wire _15698_;
 wire _15699_;
 wire _15700_;
 wire _15701_;
 wire _15702_;
 wire _15703_;
 wire _15704_;
 wire _15705_;
 wire _15706_;
 wire _15707_;
 wire _15708_;
 wire _15709_;
 wire _15710_;
 wire _15711_;
 wire _15712_;
 wire _15713_;
 wire _15714_;
 wire _15715_;
 wire _15716_;
 wire _15717_;
 wire _15718_;
 wire _15719_;
 wire _15720_;
 wire _15721_;
 wire _15722_;
 wire _15723_;
 wire _15724_;
 wire _15725_;
 wire _15726_;
 wire _15727_;
 wire _15728_;
 wire _15729_;
 wire _15730_;
 wire _15731_;
 wire _15732_;
 wire _15733_;
 wire _15734_;
 wire _15735_;
 wire _15736_;
 wire _15737_;
 wire _15738_;
 wire _15739_;
 wire _15740_;
 wire _15741_;
 wire _15742_;
 wire _15743_;
 wire _15744_;
 wire _15745_;
 wire _15746_;
 wire _15747_;
 wire _15748_;
 wire _15749_;
 wire _15750_;
 wire _15751_;
 wire _15752_;
 wire _15753_;
 wire _15754_;
 wire _15755_;
 wire _15756_;
 wire _15757_;
 wire _15758_;
 wire _15759_;
 wire _15760_;
 wire _15761_;
 wire _15762_;
 wire _15763_;
 wire _15764_;
 wire _15765_;
 wire _15766_;
 wire _15767_;
 wire _15768_;
 wire _15769_;
 wire _15770_;
 wire _15771_;
 wire _15772_;
 wire _15773_;
 wire _15774_;
 wire _15775_;
 wire _15776_;
 wire _15777_;
 wire _15778_;
 wire _15779_;
 wire _15780_;
 wire _15781_;
 wire _15782_;
 wire _15783_;
 wire _15784_;
 wire _15785_;
 wire _15786_;
 wire _15787_;
 wire _15788_;
 wire _15789_;
 wire _15790_;
 wire _15791_;
 wire _15792_;
 wire _15793_;
 wire _15794_;
 wire _15795_;
 wire _15796_;
 wire _15797_;
 wire _15798_;
 wire _15799_;
 wire _15800_;
 wire _15801_;
 wire _15802_;
 wire _15803_;
 wire _15804_;
 wire _15805_;
 wire _15806_;
 wire _15807_;
 wire _15808_;
 wire _15809_;
 wire _15810_;
 wire _15811_;
 wire _15812_;
 wire _15813_;
 wire _15814_;
 wire _15815_;
 wire _15816_;
 wire _15817_;
 wire _15818_;
 wire _15819_;
 wire _15820_;
 wire _15821_;
 wire _15822_;
 wire _15823_;
 wire _15824_;
 wire _15825_;
 wire _15826_;
 wire _15827_;
 wire _15828_;
 wire _15829_;
 wire _15830_;
 wire _15831_;
 wire _15832_;
 wire _15833_;
 wire _15834_;
 wire _15835_;
 wire _15836_;
 wire _15837_;
 wire _15838_;
 wire _15839_;
 wire _15840_;
 wire _15841_;
 wire _15842_;
 wire _15843_;
 wire _15844_;
 wire _15845_;
 wire _15846_;
 wire _15847_;
 wire _15848_;
 wire _15849_;
 wire _15850_;
 wire _15851_;
 wire _15852_;
 wire _15853_;
 wire _15854_;
 wire _15855_;
 wire _15856_;
 wire _15857_;
 wire _15858_;
 wire _15859_;
 wire _15860_;
 wire _15861_;
 wire _15862_;
 wire _15863_;
 wire _15864_;
 wire _15865_;
 wire _15866_;
 wire _15867_;
 wire _15868_;
 wire _15869_;
 wire _15870_;
 wire _15871_;
 wire _15872_;
 wire _15873_;
 wire _15874_;
 wire _15875_;
 wire _15876_;
 wire _15877_;
 wire _15878_;
 wire _15879_;
 wire _15880_;
 wire _15881_;
 wire _15882_;
 wire _15883_;
 wire _15884_;
 wire _15885_;
 wire _15886_;
 wire _15887_;
 wire _15888_;
 wire _15889_;
 wire _15890_;
 wire _15891_;
 wire _15892_;
 wire _15893_;
 wire _15894_;
 wire _15895_;
 wire _15896_;
 wire _15897_;
 wire _15898_;
 wire _15899_;
 wire _15900_;
 wire _15901_;
 wire _15902_;
 wire _15903_;
 wire _15904_;
 wire _15905_;
 wire _15906_;
 wire _15907_;
 wire _15908_;
 wire _15909_;
 wire _15910_;
 wire _15911_;
 wire _15912_;
 wire _15913_;
 wire _15914_;
 wire _15915_;
 wire _15916_;
 wire _15917_;
 wire _15918_;
 wire _15919_;
 wire _15920_;
 wire _15921_;
 wire _15922_;
 wire _15923_;
 wire _15924_;
 wire _15925_;
 wire _15926_;
 wire _15927_;
 wire _15928_;
 wire _15929_;
 wire _15930_;
 wire _15931_;
 wire _15932_;
 wire _15933_;
 wire _15934_;
 wire _15935_;
 wire _15936_;
 wire _15937_;
 wire _15938_;
 wire _15939_;
 wire _15940_;
 wire _15941_;
 wire _15942_;
 wire _15943_;
 wire _15944_;
 wire _15945_;
 wire _15946_;
 wire _15947_;
 wire _15948_;
 wire _15949_;
 wire _15950_;
 wire _15951_;
 wire _15952_;
 wire _15953_;
 wire _15954_;
 wire _15955_;
 wire _15956_;
 wire _15957_;
 wire _15958_;
 wire _15959_;
 wire _15960_;
 wire _15961_;
 wire _15962_;
 wire _15963_;
 wire _15964_;
 wire _15965_;
 wire _15966_;
 wire _15967_;
 wire _15968_;
 wire _15969_;
 wire _15970_;
 wire _15971_;
 wire _15972_;
 wire _15973_;
 wire _15974_;
 wire _15975_;
 wire _15976_;
 wire _15977_;
 wire _15978_;
 wire _15979_;
 wire _15980_;
 wire _15981_;
 wire _15982_;
 wire _15983_;
 wire _15984_;
 wire _15985_;
 wire _15986_;
 wire _15987_;
 wire _15988_;
 wire _15989_;
 wire _15990_;
 wire _15991_;
 wire _15992_;
 wire _15993_;
 wire _15994_;
 wire _15995_;
 wire _15996_;
 wire _15997_;
 wire _15998_;
 wire _15999_;
 wire _16000_;
 wire _16001_;
 wire _16002_;
 wire _16003_;
 wire _16004_;
 wire _16005_;
 wire _16006_;
 wire _16007_;
 wire _16008_;
 wire _16009_;
 wire _16010_;
 wire _16011_;
 wire _16012_;
 wire _16013_;
 wire _16014_;
 wire _16015_;
 wire _16016_;
 wire _16017_;
 wire _16018_;
 wire _16019_;
 wire _16020_;
 wire _16021_;
 wire _16022_;
 wire _16023_;
 wire _16024_;
 wire _16025_;
 wire _16026_;
 wire _16027_;
 wire _16028_;
 wire _16029_;
 wire _16030_;
 wire _16031_;
 wire _16032_;
 wire _16033_;
 wire _16034_;
 wire _16035_;
 wire _16036_;
 wire _16037_;
 wire _16038_;
 wire _16039_;
 wire _16040_;
 wire _16041_;
 wire _16042_;
 wire _16043_;
 wire _16044_;
 wire _16045_;
 wire _16046_;
 wire _16047_;
 wire _16048_;
 wire _16049_;
 wire _16050_;
 wire _16051_;
 wire _16052_;
 wire _16053_;
 wire _16054_;
 wire _16055_;
 wire _16056_;
 wire _16057_;
 wire _16058_;
 wire _16059_;
 wire _16060_;
 wire _16061_;
 wire _16062_;
 wire _16063_;
 wire _16064_;
 wire _16065_;
 wire _16066_;
 wire _16067_;
 wire _16068_;
 wire _16069_;
 wire _16070_;
 wire _16071_;
 wire _16072_;
 wire _16073_;
 wire _16074_;
 wire _16075_;
 wire _16076_;
 wire _16077_;
 wire _16078_;
 wire _16079_;
 wire _16080_;
 wire _16081_;
 wire _16082_;
 wire _16083_;
 wire _16084_;
 wire _16085_;
 wire _16086_;
 wire _16087_;
 wire _16088_;
 wire _16089_;
 wire _16090_;
 wire _16091_;
 wire _16092_;
 wire _16093_;
 wire _16094_;
 wire _16095_;
 wire _16096_;
 wire _16097_;
 wire _16098_;
 wire _16099_;
 wire _16100_;
 wire _16101_;
 wire _16102_;
 wire _16103_;
 wire _16104_;
 wire _16105_;
 wire _16106_;
 wire _16107_;
 wire _16108_;
 wire _16109_;
 wire _16110_;
 wire _16111_;
 wire _16112_;
 wire _16113_;
 wire _16114_;
 wire _16115_;
 wire _16116_;
 wire _16117_;
 wire _16118_;
 wire _16119_;
 wire _16120_;
 wire _16121_;
 wire _16122_;
 wire _16123_;
 wire _16124_;
 wire _16125_;
 wire _16126_;
 wire _16127_;
 wire _16128_;
 wire _16129_;
 wire _16130_;
 wire _16131_;
 wire _16132_;
 wire _16133_;
 wire _16134_;
 wire _16135_;
 wire _16136_;
 wire _16137_;
 wire _16138_;
 wire _16139_;
 wire _16140_;
 wire _16141_;
 wire _16142_;
 wire _16143_;
 wire _16144_;
 wire _16145_;
 wire _16146_;
 wire _16147_;
 wire _16148_;
 wire _16149_;
 wire _16150_;
 wire _16151_;
 wire _16152_;
 wire _16153_;
 wire _16154_;
 wire _16155_;
 wire _16156_;
 wire _16157_;
 wire _16158_;
 wire _16159_;
 wire _16160_;
 wire _16161_;
 wire _16162_;
 wire _16163_;
 wire _16164_;
 wire _16165_;
 wire _16166_;
 wire _16167_;
 wire _16168_;
 wire _16169_;
 wire _16170_;
 wire _16171_;
 wire _16172_;
 wire _16173_;
 wire _16174_;
 wire _16175_;
 wire _16176_;
 wire _16177_;
 wire _16178_;
 wire _16179_;
 wire _16180_;
 wire _16181_;
 wire _16182_;
 wire _16183_;
 wire _16184_;
 wire _16185_;
 wire _16186_;
 wire _16187_;
 wire _16188_;
 wire _16189_;
 wire _16190_;
 wire _16191_;
 wire _16192_;
 wire _16193_;
 wire _16194_;
 wire _16195_;
 wire _16196_;
 wire _16197_;
 wire _16198_;
 wire _16199_;
 wire _16200_;
 wire _16201_;
 wire _16202_;
 wire _16203_;
 wire _16204_;
 wire _16205_;
 wire _16206_;
 wire _16207_;
 wire _16208_;
 wire _16209_;
 wire _16210_;
 wire _16211_;
 wire _16212_;
 wire _16213_;
 wire _16214_;
 wire _16215_;
 wire _16216_;
 wire _16217_;
 wire _16218_;
 wire _16219_;
 wire _16220_;
 wire _16221_;
 wire _16222_;
 wire _16223_;
 wire _16224_;
 wire _16225_;
 wire _16226_;
 wire _16227_;
 wire _16228_;
 wire _16229_;
 wire _16230_;
 wire _16231_;
 wire _16232_;
 wire _16233_;
 wire _16234_;
 wire _16235_;
 wire _16236_;
 wire _16237_;
 wire _16238_;
 wire _16239_;
 wire _16240_;
 wire _16241_;
 wire _16242_;
 wire _16243_;
 wire _16244_;
 wire _16245_;
 wire _16246_;
 wire _16247_;
 wire _16248_;
 wire _16249_;
 wire _16250_;
 wire _16251_;
 wire _16252_;
 wire _16253_;
 wire _16254_;
 wire _16255_;
 wire _16256_;
 wire _16257_;
 wire _16258_;
 wire _16259_;
 wire _16260_;
 wire _16261_;
 wire _16262_;
 wire _16263_;
 wire _16264_;
 wire _16265_;
 wire _16266_;
 wire _16267_;
 wire _16268_;
 wire _16269_;
 wire _16270_;
 wire _16271_;
 wire _16272_;
 wire _16273_;
 wire _16274_;
 wire _16275_;
 wire _16276_;
 wire _16277_;
 wire _16278_;
 wire _16279_;
 wire _16280_;
 wire _16281_;
 wire _16282_;
 wire _16283_;
 wire _16284_;
 wire _16285_;
 wire _16286_;
 wire _16287_;
 wire _16288_;
 wire _16289_;
 wire _16290_;
 wire _16291_;
 wire _16292_;
 wire _16293_;
 wire _16294_;
 wire _16295_;
 wire _16296_;
 wire _16297_;
 wire _16298_;
 wire _16299_;
 wire _16300_;
 wire _16301_;
 wire _16302_;
 wire _16303_;
 wire _16304_;
 wire _16305_;
 wire _16306_;
 wire _16307_;
 wire _16308_;
 wire _16309_;
 wire _16310_;
 wire _16311_;
 wire _16312_;
 wire _16313_;
 wire _16314_;
 wire _16315_;
 wire _16316_;
 wire _16317_;
 wire _16318_;
 wire _16319_;
 wire _16320_;
 wire _16321_;
 wire _16322_;
 wire _16323_;
 wire _16324_;
 wire _16325_;
 wire _16326_;
 wire _16327_;
 wire _16328_;
 wire _16329_;
 wire _16330_;
 wire _16331_;
 wire _16332_;
 wire _16333_;
 wire _16334_;
 wire _16335_;
 wire _16336_;
 wire _16337_;
 wire _16338_;
 wire _16339_;
 wire _16340_;
 wire _16341_;
 wire _16342_;
 wire _16343_;
 wire _16344_;
 wire _16345_;
 wire _16346_;
 wire _16347_;
 wire _16348_;
 wire _16349_;
 wire _16350_;
 wire _16351_;
 wire _16352_;
 wire _16353_;
 wire _16354_;
 wire _16355_;
 wire _16356_;
 wire _16357_;
 wire _16358_;
 wire _16359_;
 wire _16360_;
 wire _16361_;
 wire _16362_;
 wire _16363_;
 wire _16364_;
 wire _16365_;
 wire _16366_;
 wire _16367_;
 wire _16368_;
 wire _16369_;
 wire _16370_;
 wire _16371_;
 wire _16372_;
 wire _16373_;
 wire _16374_;
 wire _16375_;
 wire _16376_;
 wire _16377_;
 wire _16378_;
 wire _16379_;
 wire _16380_;
 wire _16381_;
 wire _16382_;
 wire _16383_;
 wire _16384_;
 wire _16385_;
 wire _16386_;
 wire _16387_;
 wire _16388_;
 wire _16389_;
 wire _16390_;
 wire _16391_;
 wire _16392_;
 wire _16393_;
 wire _16394_;
 wire _16395_;
 wire _16396_;
 wire _16397_;
 wire _16398_;
 wire _16399_;
 wire _16400_;
 wire _16401_;
 wire _16402_;
 wire _16403_;
 wire _16404_;
 wire _16405_;
 wire _16406_;
 wire _16407_;
 wire _16408_;
 wire _16409_;
 wire _16410_;
 wire _16411_;
 wire _16412_;
 wire _16413_;
 wire _16414_;
 wire _16415_;
 wire _16416_;
 wire _16417_;
 wire _16418_;
 wire _16419_;
 wire _16420_;
 wire _16421_;
 wire _16422_;
 wire _16423_;
 wire _16424_;
 wire _16425_;
 wire _16426_;
 wire _16427_;
 wire _16428_;
 wire _16429_;
 wire _16430_;
 wire _16431_;
 wire _16432_;
 wire _16433_;
 wire _16434_;
 wire _16435_;
 wire _16436_;
 wire _16437_;
 wire _16438_;
 wire _16439_;
 wire _16440_;
 wire _16441_;
 wire _16442_;
 wire _16443_;
 wire _16444_;
 wire _16445_;
 wire _16446_;
 wire _16447_;
 wire _16448_;
 wire _16449_;
 wire _16450_;
 wire _16451_;
 wire _16452_;
 wire _16453_;
 wire _16454_;
 wire _16455_;
 wire _16456_;
 wire _16457_;
 wire _16458_;
 wire _16459_;
 wire _16460_;
 wire _16461_;
 wire _16462_;
 wire _16463_;
 wire _16464_;
 wire _16465_;
 wire _16466_;
 wire _16467_;
 wire _16468_;
 wire _16469_;
 wire _16470_;
 wire _16471_;
 wire _16472_;
 wire _16473_;
 wire _16474_;
 wire _16475_;
 wire _16476_;
 wire _16477_;
 wire _16478_;
 wire _16479_;
 wire _16480_;
 wire _16481_;
 wire _16482_;
 wire _16483_;
 wire _16484_;
 wire _16485_;
 wire _16486_;
 wire _16487_;
 wire _16488_;
 wire _16489_;
 wire _16490_;
 wire _16491_;
 wire _16492_;
 wire _16493_;
 wire _16494_;
 wire _16495_;
 wire _16496_;
 wire _16497_;
 wire _16498_;
 wire _16499_;
 wire _16500_;
 wire _16501_;
 wire _16502_;
 wire _16503_;
 wire _16504_;
 wire _16505_;
 wire _16506_;
 wire _16507_;
 wire _16508_;
 wire _16509_;
 wire _16510_;
 wire _16511_;
 wire _16512_;
 wire _16513_;
 wire _16514_;
 wire _16515_;
 wire _16516_;
 wire _16517_;
 wire _16518_;
 wire _16519_;
 wire _16520_;
 wire _16521_;
 wire _16522_;
 wire _16523_;
 wire _16524_;
 wire _16525_;
 wire _16526_;
 wire _16527_;
 wire _16528_;
 wire _16529_;
 wire _16530_;
 wire _16531_;
 wire _16532_;
 wire _16533_;
 wire _16534_;
 wire _16535_;
 wire _16536_;
 wire _16537_;
 wire _16538_;
 wire _16539_;
 wire _16540_;
 wire _16541_;
 wire _16542_;
 wire _16543_;
 wire _16544_;
 wire _16545_;
 wire _16546_;
 wire _16547_;
 wire _16548_;
 wire _16549_;
 wire _16550_;
 wire _16551_;
 wire _16552_;
 wire _16553_;
 wire _16554_;
 wire _16555_;
 wire _16556_;
 wire _16557_;
 wire _16558_;
 wire _16559_;
 wire _16560_;
 wire _16561_;
 wire _16562_;
 wire _16563_;
 wire _16564_;
 wire _16565_;
 wire _16566_;
 wire _16567_;
 wire _16568_;
 wire _16569_;
 wire _16570_;
 wire _16571_;
 wire _16572_;
 wire _16573_;
 wire _16574_;
 wire _16575_;
 wire _16576_;
 wire _16577_;
 wire _16578_;
 wire _16579_;
 wire _16580_;
 wire _16581_;
 wire _16582_;
 wire _16583_;
 wire _16584_;
 wire _16585_;
 wire _16586_;
 wire _16587_;
 wire _16588_;
 wire _16589_;
 wire _16590_;
 wire _16591_;
 wire _16592_;
 wire _16593_;
 wire _16594_;
 wire _16595_;
 wire _16596_;
 wire _16597_;
 wire _16598_;
 wire _16599_;
 wire _16600_;
 wire _16601_;
 wire _16602_;
 wire _16603_;
 wire _16604_;
 wire _16605_;
 wire _16606_;
 wire _16607_;
 wire _16608_;
 wire _16609_;
 wire _16610_;
 wire _16611_;
 wire _16612_;
 wire _16613_;
 wire _16614_;
 wire _16615_;
 wire _16616_;
 wire _16617_;
 wire _16618_;
 wire _16619_;
 wire _16620_;
 wire _16621_;
 wire _16622_;
 wire _16623_;
 wire _16624_;
 wire _16625_;
 wire _16626_;
 wire _16627_;
 wire _16628_;
 wire _16629_;
 wire _16630_;
 wire _16631_;
 wire _16632_;
 wire _16633_;
 wire _16634_;
 wire _16635_;
 wire _16636_;
 wire _16637_;
 wire _16638_;
 wire _16639_;
 wire _16640_;
 wire _16641_;
 wire _16642_;
 wire _16643_;
 wire _16644_;
 wire _16645_;
 wire _16646_;
 wire _16647_;
 wire _16648_;
 wire _16649_;
 wire _16650_;
 wire _16651_;
 wire _16652_;
 wire _16653_;
 wire _16654_;
 wire _16655_;
 wire _16656_;
 wire _16657_;
 wire _16658_;
 wire _16659_;
 wire _16660_;
 wire _16661_;
 wire _16662_;
 wire _16663_;
 wire _16664_;
 wire _16665_;
 wire _16666_;
 wire _16667_;
 wire _16668_;
 wire _16669_;
 wire _16670_;
 wire _16671_;
 wire _16672_;
 wire _16673_;
 wire _16674_;
 wire _16675_;
 wire _16676_;
 wire _16677_;
 wire _16678_;
 wire _16679_;
 wire _16680_;
 wire _16681_;
 wire _16682_;
 wire _16683_;
 wire _16684_;
 wire _16685_;
 wire _16686_;
 wire _16687_;
 wire _16688_;
 wire _16689_;
 wire _16690_;
 wire _16691_;
 wire _16692_;
 wire _16693_;
 wire _16694_;
 wire _16695_;
 wire _16696_;
 wire _16697_;
 wire _16698_;
 wire _16699_;
 wire _16700_;
 wire _16701_;
 wire _16702_;
 wire _16703_;
 wire _16704_;
 wire _16705_;
 wire _16706_;
 wire _16707_;
 wire _16708_;
 wire _16709_;
 wire _16710_;
 wire _16711_;
 wire _16712_;
 wire _16713_;
 wire _16714_;
 wire _16715_;
 wire _16716_;
 wire _16717_;
 wire _16718_;
 wire _16719_;
 wire _16720_;
 wire _16721_;
 wire _16722_;
 wire _16723_;
 wire _16724_;
 wire _16725_;
 wire _16726_;
 wire _16727_;
 wire _16728_;
 wire _16729_;
 wire _16730_;
 wire _16731_;
 wire _16732_;
 wire _16733_;
 wire _16734_;
 wire _16735_;
 wire _16736_;
 wire _16737_;
 wire _16738_;
 wire _16739_;
 wire _16740_;
 wire _16741_;
 wire _16742_;
 wire _16743_;
 wire _16744_;
 wire _16745_;
 wire _16746_;
 wire _16747_;
 wire _16748_;
 wire _16749_;
 wire _16750_;
 wire _16751_;
 wire _16752_;
 wire _16753_;
 wire _16754_;
 wire _16755_;
 wire _16756_;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire \gpio_uo_en[0] ;
 wire \gpio_uo_en[1] ;
 wire \gpio_uo_en[2] ;
 wire \gpio_uo_en[3] ;
 wire \gpio_uo_en[4] ;
 wire \gpio_uo_en[5] ;
 wire \gpio_uo_en[6] ;
 wire \gpio_uo_en[7] ;
 wire \gpio_uo_out[0] ;
 wire \gpio_uo_out[1] ;
 wire \gpio_uo_out[2] ;
 wire \gpio_uo_out[3] ;
 wire \gpio_uo_out[4] ;
 wire \gpio_uo_out[5] ;
 wire \gpio_uo_out[6] ;
 wire \gpio_uo_out[7] ;
 wire \led[0] ;
 wire \led[1] ;
 wire \led[2] ;
 wire \led[3] ;
 wire sclk;
 wire sio0_si_mosi_o;
 wire sio1_so_miso_o;
 wire sio2_o;
 wire sio3_o;
 wire \soc_I.IRQ3 ;
 wire \soc_I.PC[0] ;
 wire \soc_I.PC[10] ;
 wire \soc_I.PC[11] ;
 wire \soc_I.PC[12] ;
 wire \soc_I.PC[13] ;
 wire \soc_I.PC[14] ;
 wire \soc_I.PC[15] ;
 wire \soc_I.PC[1] ;
 wire \soc_I.PC[20] ;
 wire \soc_I.PC[21] ;
 wire \soc_I.PC[22] ;
 wire \soc_I.PC[23] ;
 wire \soc_I.PC[24] ;
 wire \soc_I.PC[25] ;
 wire \soc_I.PC[26] ;
 wire \soc_I.PC[27] ;
 wire \soc_I.PC[28] ;
 wire \soc_I.PC[29] ;
 wire \soc_I.PC[2] ;
 wire \soc_I.PC[30] ;
 wire \soc_I.PC[31] ;
 wire \soc_I.PC[3] ;
 wire \soc_I.PC[4] ;
 wire \soc_I.PC[5] ;
 wire \soc_I.PC[6] ;
 wire \soc_I.PC[7] ;
 wire \soc_I.PC[8] ;
 wire \soc_I.PC[9] ;
 wire \soc_I.clint_I.addr[0] ;
 wire \soc_I.clint_I.addr[1] ;
 wire \soc_I.clint_I.div[0] ;
 wire \soc_I.clint_I.div[10] ;
 wire \soc_I.clint_I.div[11] ;
 wire \soc_I.clint_I.div[12] ;
 wire \soc_I.clint_I.div[13] ;
 wire \soc_I.clint_I.div[14] ;
 wire \soc_I.clint_I.div[15] ;
 wire \soc_I.clint_I.div[1] ;
 wire \soc_I.clint_I.div[2] ;
 wire \soc_I.clint_I.div[3] ;
 wire \soc_I.clint_I.div[4] ;
 wire \soc_I.clint_I.div[5] ;
 wire \soc_I.clint_I.div[6] ;
 wire \soc_I.clint_I.div[7] ;
 wire \soc_I.clint_I.div[8] ;
 wire \soc_I.clint_I.div[9] ;
 wire \soc_I.clint_I.mtime[0] ;
 wire \soc_I.clint_I.mtime[10] ;
 wire \soc_I.clint_I.mtime[11] ;
 wire \soc_I.clint_I.mtime[12] ;
 wire \soc_I.clint_I.mtime[13] ;
 wire \soc_I.clint_I.mtime[14] ;
 wire \soc_I.clint_I.mtime[15] ;
 wire \soc_I.clint_I.mtime[16] ;
 wire \soc_I.clint_I.mtime[17] ;
 wire \soc_I.clint_I.mtime[18] ;
 wire \soc_I.clint_I.mtime[19] ;
 wire \soc_I.clint_I.mtime[1] ;
 wire \soc_I.clint_I.mtime[20] ;
 wire \soc_I.clint_I.mtime[21] ;
 wire \soc_I.clint_I.mtime[22] ;
 wire \soc_I.clint_I.mtime[23] ;
 wire \soc_I.clint_I.mtime[24] ;
 wire \soc_I.clint_I.mtime[25] ;
 wire \soc_I.clint_I.mtime[26] ;
 wire \soc_I.clint_I.mtime[27] ;
 wire \soc_I.clint_I.mtime[28] ;
 wire \soc_I.clint_I.mtime[29] ;
 wire \soc_I.clint_I.mtime[2] ;
 wire \soc_I.clint_I.mtime[30] ;
 wire \soc_I.clint_I.mtime[31] ;
 wire \soc_I.clint_I.mtime[32] ;
 wire \soc_I.clint_I.mtime[33] ;
 wire \soc_I.clint_I.mtime[34] ;
 wire \soc_I.clint_I.mtime[35] ;
 wire \soc_I.clint_I.mtime[36] ;
 wire \soc_I.clint_I.mtime[37] ;
 wire \soc_I.clint_I.mtime[38] ;
 wire \soc_I.clint_I.mtime[39] ;
 wire \soc_I.clint_I.mtime[3] ;
 wire \soc_I.clint_I.mtime[40] ;
 wire \soc_I.clint_I.mtime[41] ;
 wire \soc_I.clint_I.mtime[42] ;
 wire \soc_I.clint_I.mtime[43] ;
 wire \soc_I.clint_I.mtime[44] ;
 wire \soc_I.clint_I.mtime[45] ;
 wire \soc_I.clint_I.mtime[46] ;
 wire \soc_I.clint_I.mtime[47] ;
 wire \soc_I.clint_I.mtime[48] ;
 wire \soc_I.clint_I.mtime[49] ;
 wire \soc_I.clint_I.mtime[4] ;
 wire \soc_I.clint_I.mtime[50] ;
 wire \soc_I.clint_I.mtime[51] ;
 wire \soc_I.clint_I.mtime[52] ;
 wire \soc_I.clint_I.mtime[53] ;
 wire \soc_I.clint_I.mtime[54] ;
 wire \soc_I.clint_I.mtime[55] ;
 wire \soc_I.clint_I.mtime[56] ;
 wire \soc_I.clint_I.mtime[57] ;
 wire \soc_I.clint_I.mtime[58] ;
 wire \soc_I.clint_I.mtime[59] ;
 wire \soc_I.clint_I.mtime[5] ;
 wire \soc_I.clint_I.mtime[60] ;
 wire \soc_I.clint_I.mtime[61] ;
 wire \soc_I.clint_I.mtime[62] ;
 wire \soc_I.clint_I.mtime[63] ;
 wire \soc_I.clint_I.mtime[6] ;
 wire \soc_I.clint_I.mtime[7] ;
 wire \soc_I.clint_I.mtime[8] ;
 wire \soc_I.clint_I.mtime[9] ;
 wire \soc_I.clint_I.mtimecmp[0] ;
 wire \soc_I.clint_I.mtimecmp[10] ;
 wire \soc_I.clint_I.mtimecmp[11] ;
 wire \soc_I.clint_I.mtimecmp[12] ;
 wire \soc_I.clint_I.mtimecmp[13] ;
 wire \soc_I.clint_I.mtimecmp[14] ;
 wire \soc_I.clint_I.mtimecmp[15] ;
 wire \soc_I.clint_I.mtimecmp[16] ;
 wire \soc_I.clint_I.mtimecmp[17] ;
 wire \soc_I.clint_I.mtimecmp[18] ;
 wire \soc_I.clint_I.mtimecmp[19] ;
 wire \soc_I.clint_I.mtimecmp[1] ;
 wire \soc_I.clint_I.mtimecmp[20] ;
 wire \soc_I.clint_I.mtimecmp[21] ;
 wire \soc_I.clint_I.mtimecmp[22] ;
 wire \soc_I.clint_I.mtimecmp[23] ;
 wire \soc_I.clint_I.mtimecmp[24] ;
 wire \soc_I.clint_I.mtimecmp[25] ;
 wire \soc_I.clint_I.mtimecmp[26] ;
 wire \soc_I.clint_I.mtimecmp[27] ;
 wire \soc_I.clint_I.mtimecmp[28] ;
 wire \soc_I.clint_I.mtimecmp[29] ;
 wire \soc_I.clint_I.mtimecmp[2] ;
 wire \soc_I.clint_I.mtimecmp[30] ;
 wire \soc_I.clint_I.mtimecmp[31] ;
 wire \soc_I.clint_I.mtimecmp[32] ;
 wire \soc_I.clint_I.mtimecmp[33] ;
 wire \soc_I.clint_I.mtimecmp[34] ;
 wire \soc_I.clint_I.mtimecmp[35] ;
 wire \soc_I.clint_I.mtimecmp[36] ;
 wire \soc_I.clint_I.mtimecmp[37] ;
 wire \soc_I.clint_I.mtimecmp[38] ;
 wire \soc_I.clint_I.mtimecmp[39] ;
 wire \soc_I.clint_I.mtimecmp[3] ;
 wire \soc_I.clint_I.mtimecmp[40] ;
 wire \soc_I.clint_I.mtimecmp[41] ;
 wire \soc_I.clint_I.mtimecmp[42] ;
 wire \soc_I.clint_I.mtimecmp[43] ;
 wire \soc_I.clint_I.mtimecmp[44] ;
 wire \soc_I.clint_I.mtimecmp[45] ;
 wire \soc_I.clint_I.mtimecmp[46] ;
 wire \soc_I.clint_I.mtimecmp[47] ;
 wire \soc_I.clint_I.mtimecmp[48] ;
 wire \soc_I.clint_I.mtimecmp[49] ;
 wire \soc_I.clint_I.mtimecmp[4] ;
 wire \soc_I.clint_I.mtimecmp[50] ;
 wire \soc_I.clint_I.mtimecmp[51] ;
 wire \soc_I.clint_I.mtimecmp[52] ;
 wire \soc_I.clint_I.mtimecmp[53] ;
 wire \soc_I.clint_I.mtimecmp[54] ;
 wire \soc_I.clint_I.mtimecmp[55] ;
 wire \soc_I.clint_I.mtimecmp[56] ;
 wire \soc_I.clint_I.mtimecmp[57] ;
 wire \soc_I.clint_I.mtimecmp[58] ;
 wire \soc_I.clint_I.mtimecmp[59] ;
 wire \soc_I.clint_I.mtimecmp[5] ;
 wire \soc_I.clint_I.mtimecmp[60] ;
 wire \soc_I.clint_I.mtimecmp[61] ;
 wire \soc_I.clint_I.mtimecmp[62] ;
 wire \soc_I.clint_I.mtimecmp[63] ;
 wire \soc_I.clint_I.mtimecmp[6] ;
 wire \soc_I.clint_I.mtimecmp[7] ;
 wire \soc_I.clint_I.mtimecmp[8] ;
 wire \soc_I.clint_I.mtimecmp[9] ;
 wire \soc_I.clint_I.ready ;
 wire \soc_I.clint_I.resetn ;
 wire \soc_I.clint_I.tick_cnt[0] ;
 wire \soc_I.clint_I.tick_cnt[10] ;
 wire \soc_I.clint_I.tick_cnt[11] ;
 wire \soc_I.clint_I.tick_cnt[12] ;
 wire \soc_I.clint_I.tick_cnt[13] ;
 wire \soc_I.clint_I.tick_cnt[14] ;
 wire \soc_I.clint_I.tick_cnt[15] ;
 wire \soc_I.clint_I.tick_cnt[16] ;
 wire \soc_I.clint_I.tick_cnt[17] ;
 wire \soc_I.clint_I.tick_cnt[1] ;
 wire \soc_I.clint_I.tick_cnt[2] ;
 wire \soc_I.clint_I.tick_cnt[3] ;
 wire \soc_I.clint_I.tick_cnt[4] ;
 wire \soc_I.clint_I.tick_cnt[5] ;
 wire \soc_I.clint_I.tick_cnt[6] ;
 wire \soc_I.clint_I.tick_cnt[7] ;
 wire \soc_I.clint_I.tick_cnt[8] ;
 wire \soc_I.clint_I.tick_cnt[9] ;
 wire \soc_I.div_ready ;
 wire \soc_I.div_reg[0] ;
 wire \soc_I.div_reg[10] ;
 wire \soc_I.div_reg[11] ;
 wire \soc_I.div_reg[12] ;
 wire \soc_I.div_reg[13] ;
 wire \soc_I.div_reg[14] ;
 wire \soc_I.div_reg[15] ;
 wire \soc_I.div_reg[1] ;
 wire \soc_I.div_reg[2] ;
 wire \soc_I.div_reg[3] ;
 wire \soc_I.div_reg[4] ;
 wire \soc_I.div_reg[5] ;
 wire \soc_I.div_reg[6] ;
 wire \soc_I.div_reg[7] ;
 wire \soc_I.div_reg[8] ;
 wire \soc_I.div_reg[9] ;
 wire \soc_I.gpio0_I.rdata[0] ;
 wire \soc_I.gpio0_I.rdata[1] ;
 wire \soc_I.gpio0_I.rdata[2] ;
 wire \soc_I.gpio0_I.rdata[3] ;
 wire \soc_I.gpio0_I.rdata[4] ;
 wire \soc_I.gpio0_I.rdata[5] ;
 wire \soc_I.gpio0_I.rdata[6] ;
 wire \soc_I.gpio0_I.rdata[7] ;
 wire \soc_I.gpio0_I.ready ;
 wire \soc_I.kianv_I.Instr[0] ;
 wire \soc_I.kianv_I.Instr[10] ;
 wire \soc_I.kianv_I.Instr[11] ;
 wire \soc_I.kianv_I.Instr[12] ;
 wire \soc_I.kianv_I.Instr[13] ;
 wire \soc_I.kianv_I.Instr[14] ;
 wire \soc_I.kianv_I.Instr[15] ;
 wire \soc_I.kianv_I.Instr[16] ;
 wire \soc_I.kianv_I.Instr[17] ;
 wire \soc_I.kianv_I.Instr[18] ;
 wire \soc_I.kianv_I.Instr[19] ;
 wire \soc_I.kianv_I.Instr[1] ;
 wire \soc_I.kianv_I.Instr[20] ;
 wire \soc_I.kianv_I.Instr[21] ;
 wire \soc_I.kianv_I.Instr[22] ;
 wire \soc_I.kianv_I.Instr[23] ;
 wire \soc_I.kianv_I.Instr[24] ;
 wire \soc_I.kianv_I.Instr[25] ;
 wire \soc_I.kianv_I.Instr[26] ;
 wire \soc_I.kianv_I.Instr[27] ;
 wire \soc_I.kianv_I.Instr[28] ;
 wire \soc_I.kianv_I.Instr[29] ;
 wire \soc_I.kianv_I.Instr[2] ;
 wire \soc_I.kianv_I.Instr[30] ;
 wire \soc_I.kianv_I.Instr[31] ;
 wire \soc_I.kianv_I.Instr[3] ;
 wire \soc_I.kianv_I.Instr[4] ;
 wire \soc_I.kianv_I.Instr[5] ;
 wire \soc_I.kianv_I.Instr[6] ;
 wire \soc_I.kianv_I.Instr[7] ;
 wire \soc_I.kianv_I.Instr[8] ;
 wire \soc_I.kianv_I.Instr[9] ;
 wire \soc_I.kianv_I.amo_reserved_state_load ;
 wire \soc_I.kianv_I.control_unit_I.div_ready ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[0] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[10] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[11] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[12] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[13] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[14] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[15] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[16] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[17] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[18] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[19] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[1] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[20] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[21] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[22] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[23] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[24] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[25] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[26] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[27] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[28] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[29] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[2] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[30] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[31] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[3] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[4] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[5] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[6] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[7] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[8] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mie[9] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mip[3] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mip[7] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[0] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[10] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[11] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[12] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[13] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[14] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[15] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[16] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[17] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[18] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[19] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[1] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[20] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[21] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[22] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[23] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[24] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[25] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[26] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[27] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[28] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[29] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[2] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[30] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[31] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[3] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[4] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[5] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[6] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[7] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[8] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[9] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.privilege_mode[0] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.privilege_mode[1] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.state[0] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.state[1] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.state[2] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.state[3] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.state[4] ;
 wire \soc_I.kianv_I.control_unit_I.main_fsm_I.state[5] ;
 wire \soc_I.kianv_I.control_unit_I.mul_ready ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[5] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[6] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[7] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.A1[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[5] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[6] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[7] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.A2[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.ADDR_I.q[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.ADDR_I.q[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[5] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[6] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[7] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.ALUOut[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[5] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[6] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[7] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[5] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[6] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[7] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRDataOut[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[5] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[6] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[7] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.CSRData[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[5] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[6] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[7] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.DataLatched[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[5] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[6] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[7] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.Data[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[5] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[6] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[7] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResultOut[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[5] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[6] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[7] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.MULExtResult[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[5] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[6] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[7] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.OldPC[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[5] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[6] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[7] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.Result_I.d5[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[32] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[33] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[34] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[35] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[36] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[37] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[38] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[39] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[40] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[41] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[42] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[43] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[44] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[45] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[46] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[47] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[48] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[49] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[50] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[51] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[52] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[53] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[54] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[55] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[56] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[57] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[58] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[59] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[5] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[60] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[61] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[62] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[63] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[6] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[7] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[5] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[6] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[7] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_select ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[32] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[33] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[34] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[35] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[36] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[37] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[38] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[39] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[40] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[41] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[42] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[43] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[44] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[45] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[46] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[47] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[48] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[49] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[50] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[51] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[52] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[53] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[54] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[55] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[56] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[57] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[58] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[59] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[5] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[60] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[61] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[62] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[63] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[6] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[7] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[5] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[6] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[7] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[5] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[6] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[7] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[5] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[6] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[7] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[5] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[6] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[7] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[5] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[6] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[7] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.bit_idx[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.bit_idx[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.bit_idx[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.bit_idx[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.bit_idx[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[5] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[6] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[7] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_state[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_state[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.div_state[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[5] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[6] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[7] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.bit_idx[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.bit_idx[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.bit_idx[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.bit_idx[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.bit_idx[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[5] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[6] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[7] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[5] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[6] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[7] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[10] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[11] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[12] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[13] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[14] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[15] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[16] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[17] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[18] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[19] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[20] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[21] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[22] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[23] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[24] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[25] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[26] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[27] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[28] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[29] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[30] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[31] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[32] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[33] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[34] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[35] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[36] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[37] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[38] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[39] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[3] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[40] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[41] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[42] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[43] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[44] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[45] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[46] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[47] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[48] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[49] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[4] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[50] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[51] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[52] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[53] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[54] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[55] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[56] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[57] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[58] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[59] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[5] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[60] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[61] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[62] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[63] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[6] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[7] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[8] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.rslt[9] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.state[0] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.state[1] ;
 wire \soc_I.kianv_I.datapath_unit_I.mul_I.state[2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][9] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][0] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][10] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][11] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][12] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][13] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][14] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][15] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][16] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][17] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][18] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][19] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][1] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][20] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][21] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][22] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][23] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][24] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][25] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][26] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][27] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][28] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][29] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][2] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][30] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][31] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][3] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][4] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][5] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][6] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][7] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][8] ;
 wire \soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][9] ;
 wire \soc_I.qqspi_I.is_quad ;
 wire \soc_I.qqspi_I.rdata[0] ;
 wire \soc_I.qqspi_I.rdata[10] ;
 wire \soc_I.qqspi_I.rdata[11] ;
 wire \soc_I.qqspi_I.rdata[12] ;
 wire \soc_I.qqspi_I.rdata[13] ;
 wire \soc_I.qqspi_I.rdata[14] ;
 wire \soc_I.qqspi_I.rdata[15] ;
 wire \soc_I.qqspi_I.rdata[16] ;
 wire \soc_I.qqspi_I.rdata[17] ;
 wire \soc_I.qqspi_I.rdata[18] ;
 wire \soc_I.qqspi_I.rdata[19] ;
 wire \soc_I.qqspi_I.rdata[1] ;
 wire \soc_I.qqspi_I.rdata[20] ;
 wire \soc_I.qqspi_I.rdata[21] ;
 wire \soc_I.qqspi_I.rdata[22] ;
 wire \soc_I.qqspi_I.rdata[23] ;
 wire \soc_I.qqspi_I.rdata[24] ;
 wire \soc_I.qqspi_I.rdata[25] ;
 wire \soc_I.qqspi_I.rdata[26] ;
 wire \soc_I.qqspi_I.rdata[27] ;
 wire \soc_I.qqspi_I.rdata[28] ;
 wire \soc_I.qqspi_I.rdata[29] ;
 wire \soc_I.qqspi_I.rdata[2] ;
 wire \soc_I.qqspi_I.rdata[30] ;
 wire \soc_I.qqspi_I.rdata[31] ;
 wire \soc_I.qqspi_I.rdata[3] ;
 wire \soc_I.qqspi_I.rdata[4] ;
 wire \soc_I.qqspi_I.rdata[5] ;
 wire \soc_I.qqspi_I.rdata[6] ;
 wire \soc_I.qqspi_I.rdata[7] ;
 wire \soc_I.qqspi_I.rdata[8] ;
 wire \soc_I.qqspi_I.rdata[9] ;
 wire \soc_I.qqspi_I.ready ;
 wire \soc_I.qqspi_I.spi_buf[0] ;
 wire \soc_I.qqspi_I.spi_buf[10] ;
 wire \soc_I.qqspi_I.spi_buf[11] ;
 wire \soc_I.qqspi_I.spi_buf[12] ;
 wire \soc_I.qqspi_I.spi_buf[13] ;
 wire \soc_I.qqspi_I.spi_buf[14] ;
 wire \soc_I.qqspi_I.spi_buf[15] ;
 wire \soc_I.qqspi_I.spi_buf[16] ;
 wire \soc_I.qqspi_I.spi_buf[17] ;
 wire \soc_I.qqspi_I.spi_buf[18] ;
 wire \soc_I.qqspi_I.spi_buf[19] ;
 wire \soc_I.qqspi_I.spi_buf[1] ;
 wire \soc_I.qqspi_I.spi_buf[20] ;
 wire \soc_I.qqspi_I.spi_buf[21] ;
 wire \soc_I.qqspi_I.spi_buf[22] ;
 wire \soc_I.qqspi_I.spi_buf[23] ;
 wire \soc_I.qqspi_I.spi_buf[24] ;
 wire \soc_I.qqspi_I.spi_buf[25] ;
 wire \soc_I.qqspi_I.spi_buf[26] ;
 wire \soc_I.qqspi_I.spi_buf[27] ;
 wire \soc_I.qqspi_I.spi_buf[28] ;
 wire \soc_I.qqspi_I.spi_buf[29] ;
 wire \soc_I.qqspi_I.spi_buf[2] ;
 wire \soc_I.qqspi_I.spi_buf[30] ;
 wire \soc_I.qqspi_I.spi_buf[31] ;
 wire \soc_I.qqspi_I.spi_buf[3] ;
 wire \soc_I.qqspi_I.spi_buf[4] ;
 wire \soc_I.qqspi_I.spi_buf[5] ;
 wire \soc_I.qqspi_I.spi_buf[6] ;
 wire \soc_I.qqspi_I.spi_buf[7] ;
 wire \soc_I.qqspi_I.spi_buf[8] ;
 wire \soc_I.qqspi_I.spi_buf[9] ;
 wire \soc_I.qqspi_I.state[0] ;
 wire \soc_I.qqspi_I.state[1] ;
 wire \soc_I.qqspi_I.state[2] ;
 wire \soc_I.qqspi_I.state[3] ;
 wire \soc_I.qqspi_I.state[4] ;
 wire \soc_I.qqspi_I.state[5] ;
 wire \soc_I.qqspi_I.state[6] ;
 wire \soc_I.qqspi_I.xfer_cycles[0] ;
 wire \soc_I.qqspi_I.xfer_cycles[1] ;
 wire \soc_I.qqspi_I.xfer_cycles[2] ;
 wire \soc_I.qqspi_I.xfer_cycles[3] ;
 wire \soc_I.qqspi_I.xfer_cycles[4] ;
 wire \soc_I.qqspi_I.xfer_cycles[5] ;
 wire \soc_I.rst_cnt[0] ;
 wire \soc_I.rst_cnt[1] ;
 wire \soc_I.rst_cnt[2] ;
 wire \soc_I.rx_uart_i.bit_idx[0] ;
 wire \soc_I.rx_uart_i.bit_idx[1] ;
 wire \soc_I.rx_uart_i.bit_idx[2] ;
 wire \soc_I.rx_uart_i.data_rd ;
 wire \soc_I.rx_uart_i.fifo_i.cnt[0] ;
 wire \soc_I.rx_uart_i.fifo_i.cnt[1] ;
 wire \soc_I.rx_uart_i.fifo_i.cnt[2] ;
 wire \soc_I.rx_uart_i.fifo_i.cnt[3] ;
 wire \soc_I.rx_uart_i.fifo_i.cnt[4] ;
 wire \soc_I.rx_uart_i.fifo_i.din[0] ;
 wire \soc_I.rx_uart_i.fifo_i.din[1] ;
 wire \soc_I.rx_uart_i.fifo_i.din[2] ;
 wire \soc_I.rx_uart_i.fifo_i.din[3] ;
 wire \soc_I.rx_uart_i.fifo_i.din[4] ;
 wire \soc_I.rx_uart_i.fifo_i.din[5] ;
 wire \soc_I.rx_uart_i.fifo_i.din[6] ;
 wire \soc_I.rx_uart_i.fifo_i.din[7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[0][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[0][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[0][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[0][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[0][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[0][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[0][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[0][7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[10][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[10][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[10][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[10][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[10][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[10][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[10][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[10][7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[11][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[11][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[11][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[11][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[11][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[11][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[11][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[11][7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[12][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[12][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[12][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[12][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[12][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[12][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[12][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[12][7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[13][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[13][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[13][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[13][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[13][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[13][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[13][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[13][7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[14][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[14][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[14][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[14][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[14][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[14][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[14][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[14][7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[15][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[15][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[15][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[15][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[15][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[15][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[15][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[15][7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[1][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[1][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[1][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[1][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[1][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[1][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[1][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[1][7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[2][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[2][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[2][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[2][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[2][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[2][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[2][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[2][7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[3][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[3][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[3][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[3][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[3][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[3][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[3][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[3][7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[4][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[4][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[4][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[4][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[4][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[4][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[4][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[4][7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[5][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[5][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[5][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[5][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[5][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[5][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[5][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[5][7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[6][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[6][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[6][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[6][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[6][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[6][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[6][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[6][7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[7][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[7][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[7][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[7][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[7][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[7][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[7][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[7][7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[8][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[8][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[8][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[8][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[8][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[8][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[8][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[8][7] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[9][0] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[9][1] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[9][2] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[9][3] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[9][4] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[9][5] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[9][6] ;
 wire \soc_I.rx_uart_i.fifo_i.ram[9][7] ;
 wire \soc_I.rx_uart_i.fifo_i.rd_ptr[0] ;
 wire \soc_I.rx_uart_i.fifo_i.rd_ptr[1] ;
 wire \soc_I.rx_uart_i.fifo_i.rd_ptr[2] ;
 wire \soc_I.rx_uart_i.fifo_i.rd_ptr[3] ;
 wire \soc_I.rx_uart_i.fifo_i.wr_ptr[0] ;
 wire \soc_I.rx_uart_i.fifo_i.wr_ptr[1] ;
 wire \soc_I.rx_uart_i.fifo_i.wr_ptr[2] ;
 wire \soc_I.rx_uart_i.fifo_i.wr_ptr[3] ;
 wire \soc_I.rx_uart_i.ready ;
 wire \soc_I.rx_uart_i.return_state[0] ;
 wire \soc_I.rx_uart_i.return_state[1] ;
 wire \soc_I.rx_uart_i.rx_in_sync[0] ;
 wire \soc_I.rx_uart_i.rx_in_sync[1] ;
 wire \soc_I.rx_uart_i.rx_in_sync[2] ;
 wire \soc_I.rx_uart_i.state[0] ;
 wire \soc_I.rx_uart_i.state[1] ;
 wire \soc_I.rx_uart_i.state[2] ;
 wire \soc_I.rx_uart_i.wait_states[0] ;
 wire \soc_I.rx_uart_i.wait_states[10] ;
 wire \soc_I.rx_uart_i.wait_states[11] ;
 wire \soc_I.rx_uart_i.wait_states[12] ;
 wire \soc_I.rx_uart_i.wait_states[13] ;
 wire \soc_I.rx_uart_i.wait_states[14] ;
 wire \soc_I.rx_uart_i.wait_states[15] ;
 wire \soc_I.rx_uart_i.wait_states[16] ;
 wire \soc_I.rx_uart_i.wait_states[1] ;
 wire \soc_I.rx_uart_i.wait_states[2] ;
 wire \soc_I.rx_uart_i.wait_states[3] ;
 wire \soc_I.rx_uart_i.wait_states[4] ;
 wire \soc_I.rx_uart_i.wait_states[5] ;
 wire \soc_I.rx_uart_i.wait_states[6] ;
 wire \soc_I.rx_uart_i.wait_states[7] ;
 wire \soc_I.rx_uart_i.wait_states[8] ;
 wire \soc_I.rx_uart_i.wait_states[9] ;
 wire \soc_I.spi0_I.cen ;
 wire \soc_I.spi0_I.div[0] ;
 wire \soc_I.spi0_I.div[10] ;
 wire \soc_I.spi0_I.div[11] ;
 wire \soc_I.spi0_I.div[12] ;
 wire \soc_I.spi0_I.div[13] ;
 wire \soc_I.spi0_I.div[14] ;
 wire \soc_I.spi0_I.div[15] ;
 wire \soc_I.spi0_I.div[1] ;
 wire \soc_I.spi0_I.div[2] ;
 wire \soc_I.spi0_I.div[3] ;
 wire \soc_I.spi0_I.div[4] ;
 wire \soc_I.spi0_I.div[5] ;
 wire \soc_I.spi0_I.div[6] ;
 wire \soc_I.spi0_I.div[7] ;
 wire \soc_I.spi0_I.div[8] ;
 wire \soc_I.spi0_I.div[9] ;
 wire \soc_I.spi0_I.ready_ctrl ;
 wire \soc_I.spi0_I.ready_xfer ;
 wire \soc_I.spi0_I.rx_data[0] ;
 wire \soc_I.spi0_I.rx_data[1] ;
 wire \soc_I.spi0_I.rx_data[2] ;
 wire \soc_I.spi0_I.rx_data[3] ;
 wire \soc_I.spi0_I.rx_data[4] ;
 wire \soc_I.spi0_I.rx_data[5] ;
 wire \soc_I.spi0_I.rx_data[6] ;
 wire \soc_I.spi0_I.rx_data[7] ;
 wire \soc_I.spi0_I.sclk ;
 wire \soc_I.spi0_I.sio0_si_mosi ;
 wire \soc_I.spi0_I.spi_buf[0] ;
 wire \soc_I.spi0_I.spi_buf[1] ;
 wire \soc_I.spi0_I.spi_buf[2] ;
 wire \soc_I.spi0_I.spi_buf[3] ;
 wire \soc_I.spi0_I.spi_buf[4] ;
 wire \soc_I.spi0_I.spi_buf[5] ;
 wire \soc_I.spi0_I.spi_buf[6] ;
 wire \soc_I.spi0_I.spi_buf[7] ;
 wire \soc_I.spi0_I.state ;
 wire \soc_I.spi0_I.tick_cnt[0] ;
 wire \soc_I.spi0_I.tick_cnt[10] ;
 wire \soc_I.spi0_I.tick_cnt[11] ;
 wire \soc_I.spi0_I.tick_cnt[12] ;
 wire \soc_I.spi0_I.tick_cnt[13] ;
 wire \soc_I.spi0_I.tick_cnt[14] ;
 wire \soc_I.spi0_I.tick_cnt[15] ;
 wire \soc_I.spi0_I.tick_cnt[16] ;
 wire \soc_I.spi0_I.tick_cnt[17] ;
 wire \soc_I.spi0_I.tick_cnt[1] ;
 wire \soc_I.spi0_I.tick_cnt[2] ;
 wire \soc_I.spi0_I.tick_cnt[3] ;
 wire \soc_I.spi0_I.tick_cnt[4] ;
 wire \soc_I.spi0_I.tick_cnt[5] ;
 wire \soc_I.spi0_I.tick_cnt[6] ;
 wire \soc_I.spi0_I.tick_cnt[7] ;
 wire \soc_I.spi0_I.tick_cnt[8] ;
 wire \soc_I.spi0_I.tick_cnt[9] ;
 wire \soc_I.spi0_I.xfer_cycles[0] ;
 wire \soc_I.spi0_I.xfer_cycles[1] ;
 wire \soc_I.spi0_I.xfer_cycles[2] ;
 wire \soc_I.spi0_I.xfer_cycles[3] ;
 wire \soc_I.spi0_I.xfer_cycles[4] ;
 wire \soc_I.spi0_I.xfer_cycles[5] ;
 wire \soc_I.spi_div_ready ;
 wire \soc_I.spi_div_reg[16] ;
 wire \soc_I.spi_div_reg[17] ;
 wire \soc_I.spi_div_reg[18] ;
 wire \soc_I.spi_div_reg[19] ;
 wire \soc_I.spi_div_reg[20] ;
 wire \soc_I.spi_div_reg[21] ;
 wire \soc_I.spi_div_reg[22] ;
 wire \soc_I.spi_div_reg[23] ;
 wire \soc_I.spi_div_reg[24] ;
 wire \soc_I.spi_div_reg[25] ;
 wire \soc_I.spi_div_reg[26] ;
 wire \soc_I.spi_div_reg[27] ;
 wire \soc_I.spi_div_reg[28] ;
 wire \soc_I.spi_div_reg[29] ;
 wire \soc_I.spi_div_reg[30] ;
 wire \soc_I.spi_div_reg[31] ;
 wire \soc_I.tx_uart_i.bit_idx[0] ;
 wire \soc_I.tx_uart_i.bit_idx[1] ;
 wire \soc_I.tx_uart_i.bit_idx[2] ;
 wire \soc_I.tx_uart_i.ready ;
 wire \soc_I.tx_uart_i.return_state[0] ;
 wire \soc_I.tx_uart_i.return_state[1] ;
 wire \soc_I.tx_uart_i.state[0] ;
 wire \soc_I.tx_uart_i.state[1] ;
 wire \soc_I.tx_uart_i.tx_data_reg[0] ;
 wire \soc_I.tx_uart_i.tx_data_reg[1] ;
 wire \soc_I.tx_uart_i.tx_data_reg[2] ;
 wire \soc_I.tx_uart_i.tx_data_reg[3] ;
 wire \soc_I.tx_uart_i.tx_data_reg[4] ;
 wire \soc_I.tx_uart_i.tx_data_reg[5] ;
 wire \soc_I.tx_uart_i.tx_data_reg[6] ;
 wire \soc_I.tx_uart_i.tx_data_reg[7] ;
 wire \soc_I.tx_uart_i.tx_out ;
 wire \soc_I.tx_uart_i.wait_states[0] ;
 wire \soc_I.tx_uart_i.wait_states[10] ;
 wire \soc_I.tx_uart_i.wait_states[11] ;
 wire \soc_I.tx_uart_i.wait_states[12] ;
 wire \soc_I.tx_uart_i.wait_states[13] ;
 wire \soc_I.tx_uart_i.wait_states[14] ;
 wire \soc_I.tx_uart_i.wait_states[15] ;
 wire \soc_I.tx_uart_i.wait_states[1] ;
 wire \soc_I.tx_uart_i.wait_states[2] ;
 wire \soc_I.tx_uart_i.wait_states[3] ;
 wire \soc_I.tx_uart_i.wait_states[4] ;
 wire \soc_I.tx_uart_i.wait_states[5] ;
 wire \soc_I.tx_uart_i.wait_states[6] ;
 wire \soc_I.tx_uart_i.wait_states[7] ;
 wire \soc_I.tx_uart_i.wait_states[8] ;
 wire \soc_I.tx_uart_i.wait_states[9] ;
 wire \soc_I.uart_lsr_rdy ;
 wire \soc_I.uart_tx_ready ;
 wire net2595;
 wire net2596;
 wire net2597;
 wire clknet_leaf_0_clk;
 wire net7326;
 wire net7327;
 wire net7328;
 wire net7329;
 wire net7330;
 wire net7331;
 wire net7332;
 wire net7333;
 wire net7334;
 wire net7335;
 wire net7336;
 wire net7337;
 wire net7338;
 wire net7339;
 wire net7340;
 wire net7341;
 wire net7342;
 wire net7343;
 wire net7344;
 wire net7345;
 wire net7346;
 wire net7347;
 wire net7348;
 wire net7349;
 wire net7350;
 wire net7351;
 wire net7352;
 wire net7353;
 wire net7354;
 wire net7355;
 wire net7356;
 wire net7357;
 wire net7358;
 wire net7359;
 wire net7360;
 wire net7361;
 wire net7362;
 wire net7363;
 wire net7364;
 wire net7365;
 wire net7366;
 wire net7367;
 wire net7368;
 wire net7369;
 wire net7370;
 wire net7371;
 wire net7372;
 wire net7373;
 wire net7374;
 wire net7375;
 wire net7376;
 wire net7377;
 wire net7378;
 wire net7379;
 wire net7380;
 wire net7381;
 wire net7382;
 wire net7383;
 wire net7384;
 wire net7385;
 wire net7386;
 wire net7387;
 wire net7388;
 wire net7389;
 wire net7390;
 wire net7391;
 wire net7392;
 wire net7393;
 wire net7394;
 wire net7395;
 wire net7396;
 wire net7397;
 wire net7398;
 wire net7399;
 wire net7400;
 wire net7401;
 wire net7402;
 wire net7403;
 wire net7404;
 wire net7405;
 wire net7406;
 wire net7407;
 wire net7408;
 wire net7409;
 wire net7410;
 wire net7411;
 wire net7412;
 wire net7413;
 wire net7414;
 wire net7415;
 wire net7416;
 wire net7417;
 wire net7418;
 wire net7419;
 wire net7420;
 wire net7421;
 wire net7422;
 wire net7423;
 wire net7424;
 wire net7425;
 wire net7426;
 wire net7427;
 wire net7428;
 wire net7429;
 wire net7430;
 wire net7431;
 wire net7432;
 wire net7433;
 wire net7434;
 wire net7435;
 wire net7436;
 wire net7437;
 wire net7438;
 wire net7439;
 wire net7440;
 wire net7441;
 wire net7442;
 wire net7443;
 wire net7444;
 wire net7445;
 wire net7446;
 wire net7447;
 wire net7448;
 wire net7449;
 wire net7450;
 wire net7451;
 wire net7452;
 wire net7453;
 wire net7454;
 wire net7455;
 wire net7456;
 wire net7457;
 wire net7458;
 wire net7459;
 wire net7460;
 wire net7461;
 wire net7462;
 wire net7463;
 wire net7464;
 wire net7465;
 wire net7466;
 wire net7467;
 wire net7468;
 wire net7469;
 wire net7470;
 wire net7471;
 wire net7472;
 wire net7473;
 wire net7474;
 wire net7475;
 wire net7476;
 wire net7477;
 wire net7478;
 wire net7479;
 wire net7480;
 wire net7481;
 wire net7482;
 wire net7483;
 wire net7484;
 wire net7485;
 wire net7486;
 wire net7487;
 wire net7488;
 wire net7489;
 wire net7490;
 wire net7491;
 wire net7492;
 wire net7493;
 wire net7494;
 wire net7495;
 wire net7496;
 wire net7497;
 wire net7498;
 wire net7499;
 wire net7500;
 wire net7501;
 wire net7502;
 wire net7503;
 wire net7504;
 wire net7505;
 wire net7506;
 wire net7507;
 wire net7508;
 wire net7509;
 wire net7510;
 wire net7511;
 wire net7512;
 wire net7513;
 wire net7514;
 wire net7515;
 wire net7516;
 wire net7517;
 wire net7518;
 wire net7519;
 wire net7520;
 wire net7521;
 wire net7522;
 wire net7523;
 wire net7524;
 wire net7525;
 wire net7526;
 wire net7527;
 wire net7528;
 wire net7529;
 wire net7530;
 wire net7531;
 wire net7532;
 wire net7533;
 wire net7534;
 wire net7535;
 wire net7536;
 wire net7537;
 wire net7538;
 wire net7539;
 wire net7540;
 wire net7541;
 wire net7542;
 wire net7543;
 wire net7544;
 wire net7545;
 wire net7546;
 wire net7547;
 wire net7548;
 wire net7549;
 wire net7550;
 wire net7551;
 wire net7552;
 wire net7553;
 wire net7554;
 wire net7555;
 wire net7556;
 wire net7557;
 wire net7558;
 wire net7559;
 wire net7560;
 wire net7561;
 wire net7562;
 wire net7563;
 wire net7564;
 wire net7565;
 wire net7566;
 wire net7567;
 wire net7568;
 wire net7569;
 wire net7570;
 wire net7571;
 wire net7572;
 wire net7573;
 wire net7574;
 wire net7575;
 wire net7576;
 wire net7577;
 wire net7578;
 wire net7579;
 wire net7580;
 wire net7581;
 wire net7582;
 wire net7583;
 wire net7584;
 wire net7585;
 wire net7586;
 wire net7587;
 wire net7588;
 wire net7589;
 wire net7590;
 wire net7591;
 wire net7592;
 wire net7593;
 wire net7594;
 wire net7595;
 wire net7596;
 wire net7597;
 wire net7598;
 wire net7599;
 wire net7600;
 wire net7601;
 wire net7602;
 wire net7603;
 wire net7604;
 wire net7605;
 wire net7606;
 wire net7607;
 wire net7608;
 wire net7609;
 wire net7610;
 wire net7611;
 wire net7612;
 wire net7613;
 wire net7614;
 wire net7615;
 wire net7616;
 wire net7617;
 wire net7618;
 wire net7619;
 wire net7620;
 wire net7621;
 wire net7622;
 wire net7623;
 wire net7624;
 wire net7625;
 wire net7626;
 wire net7627;
 wire net7628;
 wire net7629;
 wire net7630;
 wire net7631;
 wire net7632;
 wire net7633;
 wire net7634;
 wire net7635;
 wire net7636;
 wire net7637;
 wire net7638;
 wire net7639;
 wire net7640;
 wire net7641;
 wire net7642;
 wire net7643;
 wire net7644;
 wire net7645;
 wire net7646;
 wire net7647;
 wire net7648;
 wire net7649;
 wire net7650;
 wire net7651;
 wire net7652;
 wire net7653;
 wire net7654;
 wire net7655;
 wire net7656;
 wire net7657;
 wire net7658;
 wire net7659;
 wire net7660;
 wire net7661;
 wire net7662;
 wire net7663;
 wire net7664;
 wire net7665;
 wire net7666;
 wire net7667;
 wire net7668;
 wire net7669;
 wire net7670;
 wire net7671;
 wire net7672;
 wire net7673;
 wire net7674;
 wire net7675;
 wire net7676;
 wire net7677;
 wire net7678;
 wire net7679;
 wire net7680;
 wire net7681;
 wire net7682;
 wire net7683;
 wire net7684;
 wire net7685;
 wire net7686;
 wire net7687;
 wire net7688;
 wire net7689;
 wire net7690;
 wire net7691;
 wire net7692;
 wire net7693;
 wire net7694;
 wire net7695;
 wire net7696;
 wire net7697;
 wire net7698;
 wire net7699;
 wire net7700;
 wire net7701;
 wire net7702;
 wire net7703;
 wire net7704;
 wire net7705;
 wire net7706;
 wire net7707;
 wire net7708;
 wire net7709;
 wire net7710;
 wire net7711;
 wire net7712;
 wire net7713;
 wire net7714;
 wire net7715;
 wire net7716;
 wire net7717;
 wire net7718;
 wire net7719;
 wire net7720;
 wire net7721;
 wire net7722;
 wire net7723;
 wire net7724;
 wire net7725;
 wire net7726;
 wire net7727;
 wire net7728;
 wire net7729;
 wire net7730;
 wire net7731;
 wire net7732;
 wire net7733;
 wire net7734;
 wire net7735;
 wire net7736;
 wire net7737;
 wire net7738;
 wire net7739;
 wire net7740;
 wire net7741;
 wire net7742;
 wire net7743;
 wire net7744;
 wire net7745;
 wire net7746;
 wire net7747;
 wire net7748;
 wire net7749;
 wire net7750;
 wire net7751;
 wire net7752;
 wire net7753;
 wire net7754;
 wire net7755;
 wire net7756;
 wire net7757;
 wire net7758;
 wire net7759;
 wire net7760;
 wire net7761;
 wire net7762;
 wire net7763;
 wire net7764;
 wire net7765;
 wire net7766;
 wire net7767;
 wire net7768;
 wire net7769;
 wire net7770;
 wire net7771;
 wire net7772;
 wire net7773;
 wire net7774;
 wire net7775;
 wire net7776;
 wire net7777;
 wire net7778;
 wire net7779;
 wire net7780;
 wire net7781;
 wire net7782;
 wire net7783;
 wire net7784;
 wire net7785;
 wire net7786;
 wire net7787;
 wire net7788;
 wire net7789;
 wire net7790;
 wire net7791;
 wire net7792;
 wire net7793;
 wire net7794;
 wire net7795;
 wire net7796;
 wire net7797;
 wire net7798;
 wire net7799;
 wire net7800;
 wire net7801;
 wire net7802;
 wire net7803;
 wire net7804;
 wire net7805;
 wire net7806;
 wire net7807;
 wire net7808;
 wire net7809;
 wire net7810;
 wire net7811;
 wire net7812;
 wire net7813;
 wire net7814;
 wire net7815;
 wire net7816;
 wire net7817;
 wire net7818;
 wire net7819;
 wire net7820;
 wire net7821;
 wire net7822;
 wire net7823;
 wire net7824;
 wire net7825;
 wire net7826;
 wire net7827;
 wire net7828;
 wire net7829;
 wire net7830;
 wire net7831;
 wire net7832;
 wire net7833;
 wire net7834;
 wire net7835;
 wire net7836;
 wire net7837;
 wire net7838;
 wire net7839;
 wire net7840;
 wire net7841;
 wire net7842;
 wire net7843;
 wire net7844;
 wire net7845;
 wire net7846;
 wire net7847;
 wire net7848;
 wire net7849;
 wire net7850;
 wire net7851;
 wire net7852;
 wire net7853;
 wire net7854;
 wire net7855;
 wire net7856;
 wire net7857;
 wire net7858;
 wire net7859;
 wire net7860;
 wire net7861;
 wire net7862;
 wire net7863;
 wire net7864;
 wire net7865;
 wire net7866;
 wire net7867;
 wire net7868;
 wire net7869;
 wire net7870;
 wire net7871;
 wire net7872;
 wire net7873;
 wire net7874;
 wire net7875;
 wire net7876;
 wire net7877;
 wire net7878;
 wire net7879;
 wire net7880;
 wire net7881;
 wire net7882;
 wire net7883;
 wire net7884;
 wire net7885;
 wire net7886;
 wire net7887;
 wire net7888;
 wire net7889;
 wire net7890;
 wire net7891;
 wire net7892;
 wire net7893;
 wire net7894;
 wire net7895;
 wire net7896;
 wire net7897;
 wire net7898;
 wire net7899;
 wire net7900;
 wire net7901;
 wire net7902;
 wire net7903;
 wire net7904;
 wire net7905;
 wire net7906;
 wire net7907;
 wire net7908;
 wire net7909;
 wire net7910;
 wire net7911;
 wire net7912;
 wire net7913;
 wire net7914;
 wire net7915;
 wire net7916;
 wire net7917;
 wire net7918;
 wire net7919;
 wire net7920;
 wire net7921;
 wire net7922;
 wire net7923;
 wire net7924;
 wire net7925;
 wire net7926;
 wire net7927;
 wire net7928;
 wire net7929;
 wire net7930;
 wire net7931;
 wire net7932;
 wire net7933;
 wire net7934;
 wire net7935;
 wire net7936;
 wire net7937;
 wire net7938;
 wire net7939;
 wire net7940;
 wire net7941;
 wire net7942;
 wire net7943;
 wire net7944;
 wire net7945;
 wire net7946;
 wire net7947;
 wire net7948;
 wire net7949;
 wire net7950;
 wire net7951;
 wire net7952;
 wire net7953;
 wire net7954;
 wire net7955;
 wire net7956;
 wire net7957;
 wire net7958;
 wire net7959;
 wire net7960;
 wire net7961;
 wire net7962;
 wire net7963;
 wire net7964;
 wire net7965;
 wire net7966;
 wire net7967;
 wire net7968;
 wire net7969;
 wire net7970;
 wire net7971;
 wire net7972;
 wire net7973;
 wire net7974;
 wire net7975;
 wire net7976;
 wire net7977;
 wire net7978;
 wire net7979;
 wire net7980;
 wire net7981;
 wire net7982;
 wire net7983;
 wire net7984;
 wire net7985;
 wire net7986;
 wire net7987;
 wire net7988;
 wire net7989;
 wire net7990;
 wire net7991;
 wire net7992;
 wire net7993;
 wire net7994;
 wire net7995;
 wire net7996;
 wire net7997;
 wire net7998;
 wire net7999;
 wire net8000;
 wire net8001;
 wire net8002;
 wire net8003;
 wire net8004;
 wire net8005;
 wire net8006;
 wire net8007;
 wire net8008;
 wire net8009;
 wire net8010;
 wire net8011;
 wire net8012;
 wire net8013;
 wire net8014;
 wire net8015;
 wire net8016;
 wire net8017;
 wire net8018;
 wire net8019;
 wire net8020;
 wire net8021;
 wire net8022;
 wire net8023;
 wire net8024;
 wire net8025;
 wire net8026;
 wire net8027;
 wire net8028;
 wire net8029;
 wire net8030;
 wire net8031;
 wire net8032;
 wire net8033;
 wire net8034;
 wire net8035;
 wire net8036;
 wire net8037;
 wire net8038;
 wire net8039;
 wire net8040;
 wire net8041;
 wire net8042;
 wire net8043;
 wire net8044;
 wire net8045;
 wire net8046;
 wire net8047;
 wire net8048;
 wire net8049;
 wire net8050;
 wire net8051;
 wire net8052;
 wire net8053;
 wire net8054;
 wire net8055;
 wire net8056;
 wire net8057;
 wire net8058;
 wire net8059;
 wire net8060;
 wire net8061;
 wire net8062;
 wire net8063;
 wire net8064;
 wire net8065;
 wire net8066;
 wire net8067;
 wire net8068;
 wire net8069;
 wire net8070;
 wire net8071;
 wire net8072;
 wire net8073;
 wire net8074;
 wire net8075;
 wire net8076;
 wire net8077;
 wire net8078;
 wire net8079;
 wire net8080;
 wire net8081;
 wire net8082;
 wire net8083;
 wire net8084;
 wire net8085;
 wire net8086;
 wire net8087;
 wire net8088;
 wire net8089;
 wire net8090;
 wire net8091;
 wire net8092;
 wire net8093;
 wire net8094;
 wire net8095;
 wire net8096;
 wire net8097;
 wire net8098;
 wire net8099;
 wire net8100;
 wire net8101;
 wire net8102;
 wire net8103;
 wire net8104;
 wire net8105;
 wire net8106;
 wire net8107;
 wire net8108;
 wire net8109;
 wire net8110;
 wire net8111;
 wire net8112;
 wire net8113;
 wire net8114;
 wire net8115;
 wire net8116;
 wire net8117;
 wire net8118;
 wire net8119;
 wire net8120;
 wire net8121;
 wire net8122;
 wire net8123;
 wire net8124;
 wire net8125;
 wire net8126;
 wire net8127;
 wire net8128;
 wire net8129;
 wire net8130;
 wire net8131;
 wire net8132;
 wire net8133;
 wire net8134;
 wire net8135;
 wire net8136;
 wire net8137;
 wire net8138;
 wire net8139;
 wire net8140;
 wire net8141;
 wire net8142;
 wire net8143;
 wire net8144;
 wire net8145;
 wire net8146;
 wire net8147;
 wire net8148;
 wire net8149;
 wire net8150;
 wire net8151;
 wire net8152;
 wire net8153;
 wire net8154;
 wire net8155;
 wire net8156;
 wire net8157;
 wire net8158;
 wire net8159;
 wire net8160;
 wire net8161;
 wire net8162;
 wire net8163;
 wire net8164;
 wire net8165;
 wire net8166;
 wire net8167;
 wire net8168;
 wire net8169;
 wire net8170;
 wire net8171;
 wire net8172;
 wire net8173;
 wire net8174;
 wire net8175;
 wire net8176;
 wire net8177;
 wire net8178;
 wire net8179;
 wire net8180;
 wire net8181;
 wire net8182;
 wire net8183;
 wire net8184;
 wire net8185;
 wire net8186;
 wire net8187;
 wire net8188;
 wire net8189;
 wire net8190;
 wire net8191;
 wire net8192;
 wire net8193;
 wire net8194;
 wire net8195;
 wire net8196;
 wire net8197;
 wire net8198;
 wire net8199;
 wire net8200;
 wire net8201;
 wire net8202;
 wire net8203;
 wire net8204;
 wire net8205;
 wire net8206;
 wire net8207;
 wire net8208;
 wire net8209;
 wire net8210;
 wire net8211;
 wire net8212;
 wire net8213;
 wire net8214;
 wire net8215;
 wire net8216;
 wire net8217;
 wire net8218;
 wire net8219;
 wire net8220;
 wire net8221;
 wire net8222;
 wire net8223;
 wire net8224;
 wire net8225;
 wire net8226;
 wire net8227;
 wire net8228;
 wire net8229;
 wire net8230;
 wire net8231;
 wire net8232;
 wire net8233;
 wire net8234;
 wire net8235;
 wire net8236;
 wire net8237;
 wire net8238;
 wire net8239;
 wire net8240;
 wire net8241;
 wire net8242;
 wire net8243;
 wire net8244;
 wire net8245;
 wire net8246;
 wire net8247;
 wire net8248;
 wire net8249;
 wire net8250;
 wire net8251;
 wire net8252;
 wire net8253;
 wire net8254;
 wire net8255;
 wire net8256;
 wire net8257;
 wire net8258;
 wire net8259;
 wire net8260;
 wire net8261;
 wire net8262;
 wire net8263;
 wire net8264;
 wire net8265;
 wire net8266;
 wire net8267;
 wire net8268;
 wire net8269;
 wire net8270;
 wire net8271;
 wire net8272;
 wire net8273;
 wire net8274;
 wire net8275;
 wire net8276;
 wire net8277;
 wire net8278;
 wire net8279;
 wire net8280;
 wire net8281;
 wire net8282;
 wire net8283;
 wire net8284;
 wire net8285;
 wire net8286;
 wire net8287;
 wire net8288;
 wire net8289;
 wire net8290;
 wire net8291;
 wire net8292;
 wire net8293;
 wire net8294;
 wire net8295;
 wire net8296;
 wire net8297;
 wire net8298;
 wire net8299;
 wire net8300;
 wire net8301;
 wire net8302;
 wire net8303;
 wire net8304;
 wire net8305;
 wire net8306;
 wire net8307;
 wire net8308;
 wire net8309;
 wire net8310;
 wire net8311;
 wire net8312;
 wire net8313;
 wire net8314;
 wire net8315;
 wire net8316;
 wire net8317;
 wire net8318;
 wire net8319;
 wire net8320;
 wire net8321;
 wire net8322;
 wire net8323;
 wire net8324;
 wire net8325;
 wire net8326;
 wire net8327;
 wire net8328;
 wire net8329;
 wire net8330;
 wire net8331;
 wire net8332;
 wire net8333;
 wire net8334;
 wire net8335;
 wire net8336;
 wire net8337;
 wire net8338;
 wire net8339;
 wire net8340;
 wire net8341;
 wire net8342;
 wire net8343;
 wire net8344;
 wire net8345;
 wire net8346;
 wire net8347;
 wire net8348;
 wire net8349;
 wire net8350;
 wire net8351;
 wire net8352;
 wire net8353;
 wire net8354;
 wire net8355;
 wire net8356;
 wire net8357;
 wire net8358;
 wire net8359;
 wire net8360;
 wire net8361;
 wire net8362;
 wire net8363;
 wire net8364;
 wire net8365;
 wire net8366;
 wire net8367;
 wire net8368;
 wire net8369;
 wire net8370;
 wire net8371;
 wire net8372;
 wire net8373;
 wire net8374;
 wire net8375;
 wire net8376;
 wire net8377;
 wire net8378;
 wire net8379;
 wire net8380;
 wire net8381;
 wire net8382;
 wire net8383;
 wire net8384;
 wire net8385;
 wire net8386;
 wire net8387;
 wire net8388;
 wire net8389;
 wire net8390;
 wire net8391;
 wire net8392;
 wire net8393;
 wire net8394;
 wire net8395;
 wire net8396;
 wire net8397;
 wire net8398;
 wire net8399;
 wire net8400;
 wire net8401;
 wire net8402;
 wire net8403;
 wire net8404;
 wire net8405;
 wire net8406;
 wire net8407;
 wire net8408;
 wire net8409;
 wire net8410;
 wire net8411;
 wire net8412;
 wire net8413;
 wire net8414;
 wire net8415;
 wire net8416;
 wire net8417;
 wire net8418;
 wire net8419;
 wire net8420;
 wire net8421;
 wire net8422;
 wire net8423;
 wire net8424;
 wire net8425;
 wire net8426;
 wire net8427;
 wire net8428;
 wire net8429;
 wire net8430;
 wire net8431;
 wire net8432;
 wire net8433;
 wire net8434;
 wire net8435;
 wire net8436;
 wire net8437;
 wire net8438;
 wire net8439;
 wire net8440;
 wire net8441;
 wire net8442;
 wire net8443;
 wire net8444;
 wire net8445;
 wire net8446;
 wire net8447;
 wire net8448;
 wire net8449;
 wire net8450;
 wire net8451;
 wire net8452;
 wire net8453;
 wire net8454;
 wire net8455;
 wire net8456;
 wire net8457;
 wire net8458;
 wire net8459;
 wire net8460;
 wire net8461;
 wire net8462;
 wire net8463;
 wire net8464;
 wire net8465;
 wire net8466;
 wire net8467;
 wire net8468;
 wire net8469;
 wire net8470;
 wire net8471;
 wire net8472;
 wire net8473;
 wire net8474;
 wire net8475;
 wire net8476;
 wire net8477;
 wire net8478;
 wire net8479;
 wire net8480;
 wire net8481;
 wire net8482;
 wire net8483;
 wire net8484;
 wire net8485;
 wire net8486;
 wire net8487;
 wire net8488;
 wire net8489;
 wire net8490;
 wire net8491;
 wire net8492;
 wire net8493;
 wire net8494;
 wire net8495;
 wire net8496;
 wire net8497;
 wire net8498;
 wire net8499;
 wire net8500;
 wire net8501;
 wire net8502;
 wire net8503;
 wire net8504;
 wire net8505;
 wire net8506;
 wire net8507;
 wire net8508;
 wire net8509;
 wire net8510;
 wire net8511;
 wire net8512;
 wire net8513;
 wire net8514;
 wire net8515;
 wire net8516;
 wire net8517;
 wire net8518;
 wire net8519;
 wire net8520;
 wire net8521;
 wire net8522;
 wire net8523;
 wire net8524;
 wire net8525;
 wire net8526;
 wire net8527;
 wire net8528;
 wire net8529;
 wire net8530;
 wire net8531;
 wire net8532;
 wire net8533;
 wire net8534;
 wire net8535;
 wire net8536;
 wire net8537;
 wire net8538;
 wire net8539;
 wire net8540;
 wire net8541;
 wire net8542;
 wire net8543;
 wire net8544;
 wire net8545;
 wire net8546;
 wire net8547;
 wire net8548;
 wire net8549;
 wire net8550;
 wire net8551;
 wire net8552;
 wire net8553;
 wire net8554;
 wire net8555;
 wire net8556;
 wire net8557;
 wire net8558;
 wire net8559;
 wire net8560;
 wire net8561;
 wire net8562;
 wire net8563;
 wire net8564;
 wire net8565;
 wire net8566;
 wire net8567;
 wire net8568;
 wire net8569;
 wire net8570;
 wire net8571;
 wire net8572;
 wire net8573;
 wire net8574;
 wire net8575;
 wire net8576;
 wire net8577;
 wire net8578;
 wire net8579;
 wire net8580;
 wire net8581;
 wire net8582;
 wire net8583;
 wire net8584;
 wire net8585;
 wire net8586;
 wire net8587;
 wire net8588;
 wire net8589;
 wire net8590;
 wire net8591;
 wire net8592;
 wire net8593;
 wire net8594;
 wire net8595;
 wire net8596;
 wire net8597;
 wire net8598;
 wire net8599;
 wire net8600;
 wire net8601;
 wire net8602;
 wire net8603;
 wire net8604;
 wire net8605;
 wire net8606;
 wire net8607;
 wire net8608;
 wire net8609;
 wire net8610;
 wire net8611;
 wire net8612;
 wire net8613;
 wire net8614;
 wire net8615;
 wire net8616;
 wire net8617;
 wire net8618;
 wire net8619;
 wire net8620;
 wire net8621;
 wire net8622;
 wire net8623;
 wire net8624;
 wire net8625;
 wire net8626;
 wire net8627;
 wire net8628;
 wire net8629;
 wire net8630;
 wire net8631;
 wire net8632;
 wire net8633;
 wire net8634;
 wire net8635;
 wire net8636;
 wire net8637;
 wire net8638;
 wire net8639;
 wire net8640;
 wire net8641;
 wire net8642;
 wire net8643;
 wire net8644;
 wire net8645;
 wire net8646;
 wire net8647;
 wire net8648;
 wire net8649;
 wire net8650;
 wire net8651;
 wire net8652;
 wire net8653;
 wire net8654;
 wire net8655;
 wire net8656;
 wire net8657;
 wire net8658;
 wire net8659;
 wire net8660;
 wire net8661;
 wire net8662;
 wire net8663;
 wire net8664;
 wire net8665;
 wire net8666;
 wire net8667;
 wire net8668;
 wire net8669;
 wire net8670;
 wire net8671;
 wire net8672;
 wire net8673;
 wire net8674;
 wire net8675;
 wire net8676;
 wire net8677;
 wire net8678;
 wire net8679;
 wire net8680;
 wire net8681;
 wire net8682;
 wire net8683;
 wire net8684;
 wire net8685;
 wire net8686;
 wire net8687;
 wire net8688;
 wire net8689;
 wire net8690;
 wire net8691;
 wire net8692;
 wire net8693;
 wire net8694;
 wire net8695;
 wire net8696;
 wire net8697;
 wire net8698;
 wire net8699;
 wire net8700;
 wire net8701;
 wire net8702;
 wire net8703;
 wire net8704;
 wire net8705;
 wire net8706;
 wire net8707;
 wire net8708;
 wire net8709;
 wire net8710;
 wire net8711;
 wire net8712;
 wire net8713;
 wire net8714;
 wire net8715;
 wire net8716;
 wire net8717;
 wire net8718;
 wire net8719;
 wire net8720;
 wire net8721;
 wire net8722;
 wire net8723;
 wire net8724;
 wire net8725;
 wire net8726;
 wire net8727;
 wire net8728;
 wire net8729;
 wire net8730;
 wire net8731;
 wire net8732;
 wire net8733;
 wire net8734;
 wire net8735;
 wire net8736;
 wire net8737;
 wire net8738;
 wire net8739;
 wire net8740;
 wire net8741;
 wire net8742;
 wire net8743;
 wire net8744;
 wire net8745;
 wire net8746;
 wire net8747;
 wire net8748;
 wire net8749;
 wire net8750;
 wire net8751;
 wire net8752;
 wire net8753;
 wire net8754;
 wire net8755;
 wire net8756;
 wire net8757;
 wire net8758;
 wire net8759;
 wire net8760;
 wire net8761;
 wire net8762;
 wire net8763;
 wire net8764;
 wire net8765;
 wire net8766;
 wire net8767;
 wire net8768;
 wire net8769;
 wire net8770;
 wire net8771;
 wire net8772;
 wire net8773;
 wire net8774;
 wire net8775;
 wire net8776;
 wire net8777;
 wire net8778;
 wire net8779;
 wire net8780;
 wire net8781;
 wire net8782;
 wire net8783;
 wire net8784;
 wire net8785;
 wire net8786;
 wire net8787;
 wire net8788;
 wire net8789;
 wire net8790;
 wire net8791;
 wire net8792;
 wire net8793;
 wire net8794;
 wire net8795;
 wire net8796;
 wire net8797;
 wire net8798;
 wire net8799;
 wire net8800;
 wire net8801;
 wire net8802;
 wire net8803;
 wire net8804;
 wire net8805;
 wire net8806;
 wire net8807;
 wire net8808;
 wire net8809;
 wire net8810;
 wire net8811;
 wire net8812;
 wire net8813;
 wire net8814;
 wire net8815;
 wire net8816;
 wire net8817;
 wire net8818;
 wire net8819;
 wire net8820;
 wire net8821;
 wire net8822;
 wire net8823;
 wire net8824;
 wire net8825;
 wire net8826;
 wire net8827;
 wire net8828;
 wire net8829;
 wire net8830;
 wire net8831;
 wire net8832;
 wire net8833;
 wire net8834;
 wire net8835;
 wire net8836;
 wire net8837;
 wire net8838;
 wire net8839;
 wire net8840;
 wire net8841;
 wire net8842;
 wire net8843;
 wire net8844;
 wire net8845;
 wire net8846;
 wire net8847;
 wire net8848;
 wire net8849;
 wire net8850;
 wire net8851;
 wire net8852;
 wire net8853;
 wire net8854;
 wire net8855;
 wire net8856;
 wire net8857;
 wire net8858;
 wire net8859;
 wire net8860;
 wire net8861;
 wire net8862;
 wire net8863;
 wire net8864;
 wire net8865;
 wire net8866;
 wire net8867;
 wire net8868;
 wire net8869;
 wire net8870;
 wire net8871;
 wire net8872;
 wire net8873;
 wire net8874;
 wire net8875;
 wire net8876;
 wire net8877;
 wire net8878;
 wire net8879;
 wire net8880;
 wire net8881;
 wire net8882;
 wire net8883;
 wire net8884;
 wire net8885;
 wire net8886;
 wire net8887;
 wire net8888;
 wire net8889;
 wire net8890;
 wire net8891;
 wire net8892;
 wire net8893;
 wire net8894;
 wire net8895;
 wire net8896;
 wire net8897;
 wire net8898;
 wire net8899;
 wire net8900;
 wire net8901;
 wire net8902;
 wire net8903;
 wire net8904;
 wire net8905;
 wire net8906;
 wire net8907;
 wire net8908;
 wire net8909;
 wire net8910;
 wire net8911;
 wire net8912;
 wire net8913;
 wire net8914;
 wire net8915;
 wire net8916;
 wire net8917;
 wire net8918;
 wire net8919;
 wire net8920;
 wire net8921;
 wire net8922;
 wire net8923;
 wire net8924;
 wire net8925;
 wire net8926;
 wire net8927;
 wire net8928;
 wire net8929;
 wire net8930;
 wire net8931;
 wire net8932;
 wire net8933;
 wire net8934;
 wire net8935;
 wire net8936;
 wire net8937;
 wire net8938;
 wire net8939;
 wire net8940;
 wire net8941;
 wire net8942;
 wire net8943;
 wire net8944;
 wire net8945;
 wire net8946;
 wire net8947;
 wire net8948;
 wire net8949;
 wire net8950;
 wire net8951;
 wire net8952;
 wire net8953;
 wire net8954;
 wire net8955;
 wire net8956;
 wire net8957;
 wire net8958;
 wire net8959;
 wire net8960;
 wire net8961;
 wire net8962;
 wire net8963;
 wire net8964;
 wire net8965;
 wire net8966;
 wire net8967;
 wire net8968;
 wire net8969;
 wire net8970;
 wire net8971;
 wire net8972;
 wire net8973;
 wire net8974;
 wire net8975;
 wire net8976;
 wire net8977;
 wire net8978;
 wire net8979;
 wire net8980;
 wire net8981;
 wire net8982;
 wire net8983;
 wire net8984;
 wire net8985;
 wire net8986;
 wire net8987;
 wire net8988;
 wire net8989;
 wire net8990;
 wire net8991;
 wire net8992;
 wire net8993;
 wire net8994;
 wire net8995;
 wire net8996;
 wire net8997;
 wire net8998;
 wire net8999;
 wire net9000;
 wire net9001;
 wire net9002;
 wire net9003;
 wire net9004;
 wire net9005;
 wire net9006;
 wire net9007;
 wire net9008;
 wire net9009;
 wire net9010;
 wire net9011;
 wire net9012;
 wire net9013;
 wire net9014;
 wire net9015;
 wire net9016;
 wire net9017;
 wire net9018;
 wire net9019;
 wire net9020;
 wire net9021;
 wire net9022;
 wire net9023;
 wire net9024;
 wire net9025;
 wire net9026;
 wire net9027;
 wire net9028;
 wire net9029;
 wire net9030;
 wire net9031;
 wire net9032;
 wire net9033;
 wire net9034;
 wire net9035;
 wire net9036;
 wire net9037;
 wire net9038;
 wire net9039;
 wire net9040;
 wire net9041;
 wire net9042;
 wire net9043;
 wire net9044;
 wire net9045;
 wire net9046;
 wire net9047;
 wire net9048;
 wire net9049;
 wire net9050;
 wire net9051;
 wire net9052;
 wire net9053;
 wire net9054;
 wire net9055;
 wire net9056;
 wire net9057;
 wire net9058;
 wire net9059;
 wire net9060;
 wire net9061;
 wire net9062;
 wire net9063;
 wire net9064;
 wire net9065;
 wire net9066;
 wire net9067;
 wire net9068;
 wire net9069;
 wire net9070;
 wire net9071;
 wire net9072;
 wire net9073;
 wire net9074;
 wire net9075;
 wire net9076;
 wire net9077;
 wire net9078;
 wire net9079;
 wire net9080;
 wire net9081;
 wire net9082;
 wire net9083;
 wire net9084;
 wire net9085;
 wire net9086;
 wire net9087;
 wire net9088;
 wire net9089;
 wire net9090;
 wire net9091;
 wire net9092;
 wire net9093;
 wire net9094;
 wire net9095;
 wire net9096;
 wire net9097;
 wire net9098;
 wire net9099;
 wire net9100;
 wire net9101;
 wire net9102;
 wire net9103;
 wire net9104;
 wire net9105;
 wire net9106;
 wire net9107;
 wire net9108;
 wire net9109;
 wire net9110;
 wire net9111;
 wire net9112;
 wire net9113;
 wire net9114;
 wire net9115;
 wire net9116;
 wire net9117;
 wire net9118;
 wire net9119;
 wire net9120;
 wire net9121;
 wire net9122;
 wire net9123;
 wire net9124;
 wire net9125;
 wire net9126;
 wire net9127;
 wire net9128;
 wire net9129;
 wire net9130;
 wire net9131;
 wire net9132;
 wire net9133;
 wire net9134;
 wire net9135;
 wire net9136;
 wire net9137;
 wire net9138;
 wire net9139;
 wire net9140;
 wire net9141;
 wire net9142;
 wire net9143;
 wire net9144;
 wire net9145;
 wire net9146;
 wire net9147;
 wire net9148;
 wire net9149;
 wire net9150;
 wire net9151;
 wire net9152;
 wire net9153;
 wire net9154;
 wire net9155;
 wire net9156;
 wire net9157;
 wire net9158;
 wire net9159;
 wire net9160;
 wire net9161;
 wire net9162;
 wire net9163;
 wire net9164;
 wire net9165;
 wire net9166;
 wire net9167;
 wire net9168;
 wire net9169;
 wire net9170;
 wire net9171;
 wire net9172;
 wire net9173;
 wire net9174;
 wire net9175;
 wire net9176;
 wire net9177;
 wire net9178;
 wire net9179;
 wire net9180;
 wire net9181;
 wire net9182;
 wire net9183;
 wire net9184;
 wire net9185;
 wire net9186;
 wire net9187;
 wire net9188;
 wire net9189;
 wire net9190;
 wire net9191;
 wire net9192;
 wire net9193;
 wire net9194;
 wire net9195;
 wire net9196;
 wire net9197;
 wire net9198;
 wire net9199;
 wire net9200;
 wire net9201;
 wire net9202;
 wire net9203;
 wire net9204;
 wire net9205;
 wire net9206;
 wire net9207;
 wire net9208;
 wire net9209;
 wire net9210;
 wire net9211;
 wire net9212;
 wire net9213;
 wire net9214;
 wire net9215;
 wire net9216;
 wire net9217;
 wire net9218;
 wire net9219;
 wire net9220;
 wire net9221;
 wire net9222;
 wire net9223;
 wire net9224;
 wire net9225;
 wire net9226;
 wire net9227;
 wire net9228;
 wire net9229;
 wire net9230;
 wire net9231;
 wire net9232;
 wire net9233;
 wire net9234;
 wire net9235;
 wire net9236;
 wire net9237;
 wire net9238;
 wire net9239;
 wire net9240;
 wire net9241;
 wire net9242;
 wire net9243;
 wire net9244;
 wire net9245;
 wire net9246;
 wire net9247;
 wire net9248;
 wire net9249;
 wire net9250;
 wire net9251;
 wire net9252;
 wire net9253;
 wire net9254;
 wire net9255;
 wire net9256;
 wire net9257;
 wire net9258;
 wire net9259;
 wire net9260;
 wire net9261;
 wire net9262;
 wire net9263;
 wire net9264;
 wire net9265;
 wire net9266;
 wire net9267;
 wire net9268;
 wire net9269;
 wire net9270;
 wire net9271;
 wire net9272;
 wire net9273;
 wire net9274;
 wire net9275;
 wire net9276;
 wire net9277;
 wire net9278;
 wire net9279;
 wire net9280;
 wire net9281;
 wire net9282;
 wire net9283;
 wire net9284;
 wire net9285;
 wire net9286;
 wire net9287;
 wire net9288;
 wire net9289;
 wire net9290;
 wire net9291;
 wire net9292;
 wire net9293;
 wire net9294;
 wire net9295;
 wire net9296;
 wire net9297;
 wire net9298;
 wire net9299;
 wire net9300;
 wire net9301;
 wire net9302;
 wire net9303;
 wire net9304;
 wire net9305;
 wire net9306;
 wire net9307;
 wire net9308;
 wire net9309;
 wire net9310;
 wire net9311;
 wire net9312;
 wire net9313;
 wire net9314;
 wire net9315;
 wire net9316;
 wire net9317;
 wire net9318;
 wire net9319;
 wire net9320;
 wire net9321;
 wire net9322;
 wire net9323;
 wire net9324;
 wire net9325;
 wire net9326;
 wire net9327;
 wire net9328;
 wire net9329;
 wire net9330;
 wire net9331;
 wire net9332;
 wire net9333;
 wire net9334;
 wire net9335;
 wire net9336;
 wire net9337;
 wire net9338;
 wire net9339;
 wire net9340;
 wire net9341;
 wire net9342;
 wire net9343;
 wire net9344;
 wire net9345;
 wire net9346;
 wire net9347;
 wire net9348;
 wire net9349;
 wire net9350;
 wire net9351;
 wire net9352;
 wire net9353;
 wire net9354;
 wire net9355;
 wire net9356;
 wire net9357;
 wire net9358;
 wire net9359;
 wire net9360;
 wire net9361;
 wire net9362;
 wire net9363;
 wire net9364;
 wire net9365;
 wire net9366;
 wire net9367;
 wire net9368;
 wire net9369;
 wire net9370;
 wire net9371;
 wire net9372;
 wire net9373;
 wire net9374;
 wire net9375;
 wire net9376;
 wire net9377;
 wire net9378;
 wire net9379;
 wire net9380;
 wire net9381;
 wire net9382;
 wire net9383;
 wire net9384;
 wire net9385;
 wire net9386;
 wire net9387;
 wire net9388;
 wire net9389;
 wire net9390;
 wire net9391;
 wire net9392;
 wire net9393;
 wire net9394;
 wire net9395;
 wire net9396;
 wire net9397;
 wire net9398;
 wire net9399;
 wire net9400;
 wire net9401;
 wire net9402;
 wire net9403;
 wire net9404;
 wire net9405;
 wire net9406;
 wire net9407;
 wire net9408;
 wire net9409;
 wire net9410;
 wire net9411;
 wire net9412;
 wire net9413;
 wire net9414;
 wire net9415;
 wire net9416;
 wire net9417;
 wire net9418;
 wire net9419;
 wire net9420;
 wire net9421;
 wire net9422;
 wire net9423;
 wire net9424;
 wire net9425;
 wire net9426;
 wire net9427;
 wire net9428;
 wire net9429;
 wire net9430;
 wire net9431;
 wire net9432;
 wire net9433;
 wire net9434;
 wire net9435;
 wire net9436;
 wire net9437;
 wire net9438;
 wire net9439;
 wire net9440;
 wire net9441;
 wire net9442;
 wire net9443;
 wire net9444;
 wire net9445;
 wire net9446;
 wire net9447;
 wire net9448;
 wire net9449;
 wire net9450;
 wire net9451;
 wire net9452;
 wire net9453;
 wire net9454;
 wire net9455;
 wire net9456;
 wire net9457;
 wire net9458;
 wire net9459;
 wire net9460;
 wire net9461;
 wire net9462;
 wire net9463;
 wire net9464;
 wire net9465;
 wire net9466;
 wire net9467;
 wire net9468;
 wire net9469;
 wire net9470;
 wire net9471;
 wire net9472;
 wire net9473;
 wire net9474;
 wire net9475;
 wire net9476;
 wire net9477;
 wire net9478;
 wire net9479;
 wire net9480;
 wire net9481;
 wire net9482;
 wire net9483;
 wire net9484;
 wire net9485;
 wire net9486;
 wire net9487;
 wire net9488;
 wire net9489;
 wire net9490;
 wire net9491;
 wire net9492;
 wire net9493;
 wire net9494;
 wire net9495;
 wire net9496;
 wire net9497;
 wire net9498;
 wire net9499;
 wire net9500;
 wire net9501;
 wire net9502;
 wire net9503;
 wire net9504;
 wire net9505;
 wire net9506;
 wire net9507;
 wire net9508;
 wire net9509;
 wire net9510;
 wire net9511;
 wire net9512;
 wire net9513;
 wire net9514;
 wire net9515;
 wire net9516;
 wire net9517;
 wire net9518;
 wire net9519;
 wire net9520;
 wire net9521;
 wire net9522;
 wire net9523;
 wire net9524;
 wire net9525;
 wire net9526;
 wire net9527;
 wire net9528;
 wire net9529;
 wire net9530;
 wire net9531;
 wire net9532;
 wire net9533;
 wire net9534;
 wire net9535;
 wire net9536;
 wire net9537;
 wire net9538;
 wire net9539;
 wire net9540;
 wire net9541;
 wire net9542;
 wire net9543;
 wire net9544;
 wire net9545;
 wire net9546;
 wire net9547;
 wire net9548;
 wire net9549;
 wire net9550;
 wire net9551;
 wire net9552;
 wire net9553;
 wire net9554;
 wire net9555;
 wire net9556;
 wire net9557;
 wire net9558;
 wire net9559;
 wire net9560;
 wire net9561;
 wire net9562;
 wire net9563;
 wire net9564;
 wire net9565;
 wire net9566;
 wire net9567;
 wire net9568;
 wire net9569;
 wire net9570;
 wire net9571;
 wire net9572;
 wire net9573;
 wire net9574;
 wire net9575;
 wire net9576;
 wire net9577;
 wire net9578;
 wire net9579;
 wire net9580;
 wire net9581;
 wire net9582;
 wire net9583;
 wire net9584;
 wire net9585;
 wire net9586;
 wire net9587;
 wire net9588;
 wire net9589;
 wire net9590;
 wire net9591;
 wire net9592;
 wire net9593;
 wire net9594;
 wire net9595;
 wire net9596;
 wire net9597;
 wire net9598;
 wire net9599;
 wire net9600;
 wire net9601;
 wire net9602;
 wire net9603;
 wire net9604;
 wire net9605;
 wire net9606;
 wire net9607;
 wire net9608;
 wire net9609;
 wire net9610;
 wire net9611;
 wire net9612;
 wire net9613;
 wire net9614;
 wire net9615;
 wire net9616;
 wire net9617;
 wire net9618;
 wire net9619;
 wire net9620;
 wire net9621;
 wire net9622;
 wire net9623;
 wire net9624;
 wire net9625;
 wire net9626;
 wire net9627;
 wire net9628;
 wire net9629;
 wire net9630;
 wire net9631;
 wire net9632;
 wire net9633;
 wire net9634;
 wire net9635;
 wire net9636;
 wire net9637;
 wire net9638;
 wire net9639;
 wire net9640;
 wire net9641;
 wire net9642;
 wire net9643;
 wire net9644;
 wire net9645;
 wire net9646;
 wire net9647;
 wire net9648;
 wire net9649;
 wire net9650;
 wire net9651;
 wire net9652;
 wire net9653;
 wire net9654;
 wire net9655;
 wire net9656;
 wire net9657;
 wire net9658;
 wire net9659;
 wire net9660;
 wire net9661;
 wire net9662;
 wire net9663;
 wire net9664;
 wire net9665;
 wire net9666;
 wire net9667;
 wire net9668;
 wire net9669;
 wire net9670;
 wire net9671;
 wire net9672;
 wire net9673;
 wire net9674;
 wire net9675;
 wire net9676;
 wire net9677;
 wire net9678;
 wire net9679;
 wire net9680;
 wire net9681;
 wire net9682;
 wire net9683;
 wire net9684;
 wire net9685;
 wire net9686;
 wire net9687;
 wire net9688;
 wire net9689;
 wire net9690;
 wire net9691;
 wire net9692;
 wire net9693;
 wire net9694;
 wire net9695;
 wire net9696;
 wire net9697;
 wire net9698;
 wire net9699;
 wire net9700;
 wire net9701;
 wire net9702;
 wire net9703;
 wire net9704;
 wire net9705;
 wire net9706;
 wire net9707;
 wire net9708;
 wire net9709;
 wire net9710;
 wire net9711;
 wire net9712;
 wire net9713;
 wire net9714;
 wire net9715;
 wire net9716;
 wire net9717;
 wire net9718;
 wire net9719;
 wire net9720;
 wire net9721;
 wire net9722;
 wire net9723;
 wire net9724;
 wire net9725;
 wire net9726;
 wire net9727;
 wire net9728;
 wire net9729;
 wire net9730;
 wire net9731;
 wire net9732;
 wire net9733;
 wire net9734;
 wire net9735;
 wire net9736;
 wire net9737;
 wire net9738;
 wire net9739;
 wire net9740;
 wire net9741;
 wire net9742;
 wire net9743;
 wire net9744;
 wire net9745;
 wire net9746;
 wire net9747;
 wire net9748;
 wire net9749;
 wire net9750;
 wire net9751;
 wire net9752;
 wire net9753;
 wire net9754;
 wire net9755;
 wire net9756;
 wire net9757;
 wire net9758;
 wire net9759;
 wire net9760;
 wire net9761;
 wire net9762;
 wire net9763;
 wire net9764;
 wire net9765;
 wire net9766;
 wire net9767;
 wire net9768;
 wire net9769;
 wire net9770;
 wire net9771;
 wire net9772;
 wire net9773;
 wire net9774;
 wire net9775;
 wire net9776;
 wire net9777;
 wire net9778;
 wire net9779;
 wire net9780;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_237_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_245_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_247_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_251_clk;
 wire clknet_leaf_252_clk;
 wire clknet_leaf_253_clk;
 wire clknet_leaf_254_clk;
 wire clknet_leaf_255_clk;
 wire clknet_leaf_256_clk;
 wire clknet_leaf_257_clk;
 wire clknet_leaf_258_clk;
 wire clknet_leaf_259_clk;
 wire clknet_leaf_260_clk;
 wire clknet_leaf_261_clk;
 wire clknet_leaf_262_clk;
 wire clknet_leaf_263_clk;
 wire clknet_leaf_264_clk;
 wire clknet_leaf_265_clk;
 wire clknet_leaf_266_clk;
 wire clknet_leaf_267_clk;
 wire clknet_leaf_268_clk;
 wire clknet_leaf_269_clk;
 wire clknet_leaf_270_clk;
 wire clknet_leaf_271_clk;
 wire clknet_leaf_272_clk;
 wire clknet_leaf_273_clk;
 wire clknet_leaf_274_clk;
 wire clknet_leaf_275_clk;
 wire clknet_leaf_276_clk;
 wire clknet_leaf_277_clk;
 wire clknet_leaf_278_clk;
 wire clknet_leaf_279_clk;
 wire clknet_leaf_280_clk;
 wire clknet_leaf_281_clk;
 wire clknet_leaf_282_clk;
 wire clknet_leaf_283_clk;
 wire clknet_leaf_284_clk;
 wire clknet_leaf_285_clk;
 wire clknet_leaf_286_clk;
 wire clknet_leaf_287_clk;
 wire clknet_leaf_288_clk;
 wire clknet_leaf_289_clk;
 wire clknet_leaf_290_clk;
 wire clknet_leaf_291_clk;
 wire clknet_leaf_292_clk;
 wire clknet_leaf_293_clk;
 wire clknet_leaf_294_clk;
 wire clknet_leaf_295_clk;
 wire clknet_leaf_296_clk;
 wire clknet_leaf_297_clk;
 wire clknet_leaf_298_clk;
 wire clknet_leaf_299_clk;
 wire clknet_leaf_300_clk;
 wire clknet_leaf_301_clk;
 wire clknet_leaf_302_clk;
 wire clknet_leaf_303_clk;
 wire clknet_leaf_304_clk;
 wire clknet_leaf_305_clk;
 wire clknet_leaf_306_clk;
 wire clknet_leaf_307_clk;
 wire clknet_leaf_308_clk;
 wire clknet_leaf_309_clk;
 wire clknet_leaf_310_clk;
 wire clknet_leaf_311_clk;
 wire clknet_leaf_312_clk;
 wire clknet_leaf_313_clk;
 wire clknet_leaf_314_clk;
 wire clknet_leaf_315_clk;
 wire clknet_leaf_316_clk;
 wire clknet_leaf_317_clk;
 wire clknet_leaf_318_clk;
 wire clknet_leaf_319_clk;
 wire clknet_leaf_320_clk;
 wire clknet_leaf_321_clk;
 wire clknet_leaf_322_clk;
 wire clknet_leaf_323_clk;
 wire clknet_leaf_324_clk;
 wire clknet_leaf_325_clk;
 wire clknet_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire clknet_5_0_0_clk;
 wire clknet_5_1_0_clk;
 wire clknet_5_2_0_clk;
 wire clknet_5_3_0_clk;
 wire clknet_5_4_0_clk;
 wire clknet_5_5_0_clk;
 wire clknet_5_6_0_clk;
 wire clknet_5_7_0_clk;
 wire clknet_5_8_0_clk;
 wire clknet_5_9_0_clk;
 wire clknet_5_10_0_clk;
 wire clknet_5_11_0_clk;
 wire clknet_5_12_0_clk;
 wire clknet_5_13_0_clk;
 wire clknet_5_14_0_clk;
 wire clknet_5_15_0_clk;
 wire clknet_5_16_0_clk;
 wire clknet_5_17_0_clk;
 wire clknet_5_18_0_clk;
 wire clknet_5_19_0_clk;
 wire clknet_5_20_0_clk;
 wire clknet_5_21_0_clk;
 wire clknet_5_22_0_clk;
 wire clknet_5_23_0_clk;
 wire clknet_5_24_0_clk;
 wire clknet_5_25_0_clk;
 wire clknet_5_26_0_clk;
 wire clknet_5_27_0_clk;
 wire clknet_5_28_0_clk;
 wire clknet_5_29_0_clk;
 wire clknet_5_30_0_clk;
 wire clknet_5_31_0_clk;
 wire clknet_6_0__leaf_clk;
 wire clknet_6_1__leaf_clk;
 wire clknet_6_2__leaf_clk;
 wire clknet_6_3__leaf_clk;
 wire clknet_6_4__leaf_clk;
 wire clknet_6_5__leaf_clk;
 wire clknet_6_6__leaf_clk;
 wire clknet_6_7__leaf_clk;
 wire clknet_6_8__leaf_clk;
 wire clknet_6_9__leaf_clk;
 wire clknet_6_10__leaf_clk;
 wire clknet_6_11__leaf_clk;
 wire clknet_6_12__leaf_clk;
 wire clknet_6_13__leaf_clk;
 wire clknet_6_14__leaf_clk;
 wire clknet_6_15__leaf_clk;
 wire clknet_6_16__leaf_clk;
 wire clknet_6_17__leaf_clk;
 wire clknet_6_18__leaf_clk;
 wire clknet_6_19__leaf_clk;
 wire clknet_6_20__leaf_clk;
 wire clknet_6_21__leaf_clk;
 wire clknet_6_22__leaf_clk;
 wire clknet_6_23__leaf_clk;
 wire clknet_6_24__leaf_clk;
 wire clknet_6_25__leaf_clk;
 wire clknet_6_26__leaf_clk;
 wire clknet_6_27__leaf_clk;
 wire clknet_6_28__leaf_clk;
 wire clknet_6_29__leaf_clk;
 wire clknet_6_30__leaf_clk;
 wire clknet_6_31__leaf_clk;
 wire clknet_6_32__leaf_clk;
 wire clknet_6_33__leaf_clk;
 wire clknet_6_34__leaf_clk;
 wire clknet_6_35__leaf_clk;
 wire clknet_6_36__leaf_clk;
 wire clknet_6_37__leaf_clk;
 wire clknet_6_38__leaf_clk;
 wire clknet_6_39__leaf_clk;
 wire clknet_6_40__leaf_clk;
 wire clknet_6_41__leaf_clk;
 wire clknet_6_42__leaf_clk;
 wire clknet_6_43__leaf_clk;
 wire clknet_6_44__leaf_clk;
 wire clknet_6_45__leaf_clk;
 wire clknet_6_46__leaf_clk;
 wire clknet_6_47__leaf_clk;
 wire clknet_6_48__leaf_clk;
 wire clknet_6_49__leaf_clk;
 wire clknet_6_50__leaf_clk;
 wire clknet_6_51__leaf_clk;
 wire clknet_6_52__leaf_clk;
 wire clknet_6_53__leaf_clk;
 wire clknet_6_54__leaf_clk;
 wire clknet_6_55__leaf_clk;
 wire clknet_6_56__leaf_clk;
 wire clknet_6_57__leaf_clk;
 wire clknet_6_58__leaf_clk;
 wire clknet_6_59__leaf_clk;
 wire clknet_6_60__leaf_clk;
 wire clknet_6_61__leaf_clk;
 wire clknet_6_62__leaf_clk;
 wire clknet_6_63__leaf_clk;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3654;
 wire net3655;
 wire net3656;
 wire net3657;
 wire net3658;
 wire net3659;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3677;
 wire net3678;
 wire net3679;
 wire net3680;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net3750;
 wire net3751;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3764;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3773;
 wire net3774;
 wire net3775;
 wire net3776;
 wire net3777;
 wire net3778;
 wire net3779;
 wire net3780;
 wire net3781;
 wire net3782;
 wire net3783;
 wire net3784;
 wire net3785;
 wire net3786;
 wire net3787;
 wire net3788;
 wire net3789;
 wire net3790;
 wire net3791;
 wire net3792;
 wire net3793;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net3799;
 wire net3800;
 wire net3801;
 wire net3802;
 wire net3803;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3807;
 wire net3808;
 wire net3809;
 wire net3810;
 wire net3811;
 wire net3812;
 wire net3813;
 wire net3814;
 wire net3815;
 wire net3816;
 wire net3817;
 wire net3818;
 wire net3819;
 wire net3820;
 wire net3821;
 wire net3822;
 wire net3823;
 wire net3824;
 wire net3825;
 wire net3826;
 wire net3827;
 wire net3828;
 wire net3829;
 wire net3830;
 wire net3831;
 wire net3832;
 wire net3833;
 wire net3834;
 wire net3835;
 wire net3836;
 wire net3837;
 wire net3838;
 wire net3839;
 wire net3840;
 wire net3841;
 wire net3842;
 wire net3843;
 wire net3844;
 wire net3845;
 wire net3846;
 wire net3847;
 wire net3848;
 wire net3849;
 wire net3850;
 wire net3851;
 wire net3852;
 wire net3853;
 wire net3854;
 wire net3855;
 wire net3856;
 wire net3857;
 wire net3858;
 wire net3859;
 wire net3860;
 wire net3861;
 wire net3862;
 wire net3863;
 wire net3864;
 wire net3865;
 wire net3866;
 wire net3867;
 wire net3868;
 wire net3869;
 wire net3870;
 wire net3871;
 wire net3872;
 wire net3873;
 wire net3874;
 wire net3875;
 wire net3876;
 wire net3877;
 wire net3878;
 wire net3879;
 wire net3880;
 wire net3881;
 wire net3882;
 wire net3883;
 wire net3884;
 wire net3885;
 wire net3886;
 wire net3887;
 wire net3888;
 wire net3889;
 wire net3890;
 wire net3891;
 wire net3892;
 wire net3893;
 wire net3894;
 wire net3895;
 wire net3896;
 wire net3897;
 wire net3898;
 wire net3899;
 wire net3900;
 wire net3901;
 wire net3902;
 wire net3903;
 wire net3904;
 wire net3905;
 wire net3906;
 wire net3907;
 wire net3908;
 wire net3909;
 wire net3910;
 wire net3911;
 wire net3912;
 wire net3913;
 wire net3914;
 wire net3915;
 wire net3916;
 wire net3917;
 wire net3918;
 wire net3919;
 wire net3920;
 wire net3921;
 wire net3922;
 wire net3923;
 wire net3924;
 wire net3925;
 wire net3926;
 wire net3927;
 wire net3928;
 wire net3929;
 wire net3930;
 wire net3931;
 wire net3932;
 wire net3933;
 wire net3934;
 wire net3935;
 wire net3936;
 wire net3937;
 wire net3938;
 wire net3939;
 wire net3940;
 wire net3941;
 wire net3942;
 wire net3943;
 wire net3944;
 wire net3945;
 wire net3946;
 wire net3947;
 wire net3948;
 wire net3949;
 wire net3950;
 wire net3951;
 wire net3952;
 wire net3953;
 wire net3954;
 wire net3955;
 wire net3956;
 wire net3957;
 wire net3958;
 wire net3959;
 wire net3960;
 wire net3961;
 wire net3962;
 wire net3963;
 wire net3964;
 wire net3965;
 wire net3966;
 wire net3967;
 wire net3968;
 wire net3969;
 wire net3970;
 wire net3971;
 wire net3972;
 wire net3973;
 wire net3974;
 wire net3975;
 wire net3976;
 wire net3977;
 wire net3978;
 wire net3979;
 wire net3980;
 wire net3981;
 wire net3982;
 wire net3983;
 wire net3984;
 wire net3985;
 wire net3986;
 wire net3987;
 wire net3988;
 wire net3989;
 wire net3990;
 wire net3991;
 wire net3992;
 wire net3993;
 wire net3994;
 wire net3995;
 wire net3996;
 wire net3997;
 wire net3998;
 wire net3999;
 wire net4000;
 wire net4001;
 wire net4002;
 wire net4003;
 wire net4004;
 wire net4005;
 wire net4006;
 wire net4007;
 wire net4008;
 wire net4009;
 wire net4010;
 wire net4011;
 wire net4012;
 wire net4013;
 wire net4014;
 wire net4015;
 wire net4016;
 wire net4017;
 wire net4018;
 wire net4019;
 wire net4020;
 wire net4021;
 wire net4022;
 wire net4023;
 wire net4024;
 wire net4025;
 wire net4026;
 wire net4027;
 wire net4028;
 wire net4029;
 wire net4030;
 wire net4031;
 wire net4032;
 wire net4033;
 wire net4034;
 wire net4035;
 wire net4036;
 wire net4037;
 wire net4038;
 wire net4039;
 wire net4040;
 wire net4041;
 wire net4042;
 wire net4043;
 wire net4044;
 wire net4045;
 wire net4046;
 wire net4047;
 wire net4048;
 wire net4049;
 wire net4050;
 wire net4051;
 wire net4052;
 wire net4053;
 wire net4054;
 wire net4055;
 wire net4056;
 wire net4057;
 wire net4058;
 wire net4059;
 wire net4060;
 wire net4061;
 wire net4062;
 wire net4063;
 wire net4064;
 wire net4065;
 wire net4066;
 wire net4067;
 wire net4068;
 wire net4069;
 wire net4070;
 wire net4071;
 wire net4072;
 wire net4073;
 wire net4074;
 wire net4075;
 wire net4076;
 wire net4077;
 wire net4078;
 wire net4079;
 wire net4080;
 wire net4081;
 wire net4082;
 wire net4083;
 wire net4084;
 wire net4085;
 wire net4086;
 wire net4087;
 wire net4088;
 wire net4089;
 wire net4090;
 wire net4091;
 wire net4092;
 wire net4093;
 wire net4094;
 wire net4095;
 wire net4096;
 wire net4097;
 wire net4098;
 wire net4099;
 wire net4100;
 wire net4101;
 wire net4102;
 wire net4103;
 wire net4104;
 wire net4105;
 wire net4106;
 wire net4107;
 wire net4108;
 wire net4109;
 wire net4110;
 wire net4111;
 wire net4112;
 wire net4113;
 wire net4114;
 wire net4115;
 wire net4116;
 wire net4117;
 wire net4118;
 wire net4119;
 wire net4120;
 wire net4121;
 wire net4122;
 wire net4123;
 wire net4124;
 wire net4125;
 wire net4126;
 wire net4127;
 wire net4128;
 wire net4129;
 wire net4130;
 wire net4131;
 wire net4132;
 wire net4133;
 wire net4134;
 wire net4135;
 wire net4136;
 wire net4137;
 wire net4138;
 wire net4139;
 wire net4140;
 wire net4141;
 wire net4142;
 wire net4143;
 wire net4144;
 wire net4145;
 wire net4146;
 wire net4147;
 wire net4148;
 wire net4149;
 wire net4150;
 wire net4151;
 wire net4152;
 wire net4153;
 wire net4154;
 wire net4155;
 wire net4156;
 wire net4157;
 wire net4158;
 wire net4159;
 wire net4160;
 wire net4161;
 wire net4162;
 wire net4163;
 wire net4164;
 wire net4165;
 wire net4166;
 wire net4167;
 wire net4168;
 wire net4169;
 wire net4170;
 wire net4171;
 wire net4172;
 wire net4173;
 wire net4174;
 wire net4175;
 wire net4176;
 wire net4177;
 wire net4178;
 wire net4179;
 wire net4180;
 wire net4181;
 wire net4182;
 wire net4183;
 wire net4184;
 wire net4185;
 wire net4186;
 wire net4187;
 wire net4188;
 wire net4189;
 wire net4190;
 wire net4191;
 wire net4192;
 wire net4193;
 wire net4194;
 wire net4195;
 wire net4196;
 wire net4197;
 wire net4198;
 wire net4199;
 wire net4200;
 wire net4201;
 wire net4202;
 wire net4203;
 wire net4204;
 wire net4205;
 wire net4206;
 wire net4207;
 wire net4208;
 wire net4209;
 wire net4210;
 wire net4211;
 wire net4212;
 wire net4213;
 wire net4214;
 wire net4215;
 wire net4216;
 wire net4217;
 wire net4218;
 wire net4219;
 wire net4220;
 wire net4221;
 wire net4222;
 wire net4223;
 wire net4224;
 wire net4225;
 wire net4226;
 wire net4227;
 wire net4228;
 wire net4229;
 wire net4230;
 wire net4231;
 wire net4232;
 wire net4233;
 wire net4234;
 wire net4235;
 wire net4236;
 wire net4237;
 wire net4238;
 wire net4239;
 wire net4240;
 wire net4241;
 wire net4242;
 wire net4243;
 wire net4244;
 wire net4245;
 wire net4246;
 wire net4247;
 wire net4248;
 wire net4249;
 wire net4250;
 wire net4251;
 wire net4252;
 wire net4253;
 wire net4254;
 wire net4255;
 wire net4256;
 wire net4257;
 wire net4258;
 wire net4259;
 wire net4260;
 wire net4261;
 wire net4262;
 wire net4263;
 wire net4264;
 wire net4265;
 wire net4266;
 wire net4267;
 wire net4268;
 wire net4269;
 wire net4270;
 wire net4271;
 wire net4272;
 wire net4273;
 wire net4274;
 wire net4275;
 wire net4276;
 wire net4277;
 wire net4278;
 wire net4279;
 wire net4280;
 wire net4281;
 wire net4282;
 wire net4283;
 wire net4284;
 wire net4285;
 wire net4286;
 wire net4287;
 wire net4288;
 wire net4289;
 wire net4290;
 wire net4291;
 wire net4292;
 wire net4293;
 wire net4294;
 wire net4295;
 wire net4296;
 wire net4297;
 wire net4298;
 wire net4299;
 wire net4300;
 wire net4301;
 wire net4302;
 wire net4303;
 wire net4304;
 wire net4305;
 wire net4306;
 wire net4307;
 wire net4308;
 wire net4309;
 wire net4310;
 wire net4311;
 wire net4312;
 wire net4313;
 wire net4314;
 wire net4315;
 wire net4316;
 wire net4317;
 wire net4318;
 wire net4319;
 wire net4320;
 wire net4321;
 wire net4322;
 wire net4323;
 wire net4324;
 wire net4325;
 wire net4326;
 wire net4327;
 wire net4328;
 wire net4329;
 wire net4330;
 wire net4331;
 wire net4332;
 wire net4333;
 wire net4334;
 wire net4335;
 wire net4336;
 wire net4337;
 wire net4338;
 wire net4339;
 wire net4340;
 wire net4341;
 wire net4342;
 wire net4343;
 wire net4344;
 wire net4345;
 wire net4346;
 wire net4347;
 wire net4348;
 wire net4349;
 wire net4350;
 wire net4351;
 wire net4352;
 wire net4353;
 wire net4354;
 wire net4355;
 wire net4356;
 wire net4357;
 wire net4358;
 wire net4359;
 wire net4360;
 wire net4361;
 wire net4362;
 wire net4363;
 wire net4364;
 wire net4365;
 wire net4366;
 wire net4367;
 wire net4368;
 wire net4369;
 wire net4370;
 wire net4371;
 wire net4372;
 wire net4373;
 wire net4374;
 wire net4375;
 wire net4376;
 wire net4377;
 wire net4378;
 wire net4379;
 wire net4380;
 wire net4381;
 wire net4382;
 wire net4383;
 wire net4384;
 wire net4385;
 wire net4386;
 wire net4387;
 wire net4388;
 wire net4389;
 wire net4390;
 wire net4391;
 wire net4392;
 wire net4393;
 wire net4394;
 wire net4395;
 wire net4396;
 wire net4397;
 wire net4398;
 wire net4399;
 wire net4400;
 wire net4401;
 wire net4402;
 wire net4403;
 wire net4404;
 wire net4405;
 wire net4406;
 wire net4407;
 wire net4408;
 wire net4409;
 wire net4410;
 wire net4411;
 wire net4412;
 wire net4413;
 wire net4414;
 wire net4415;
 wire net4416;
 wire net4417;
 wire net4418;
 wire net4419;
 wire net4420;
 wire net4421;
 wire net4422;
 wire net4423;
 wire net4424;
 wire net4425;
 wire net4426;
 wire net4427;
 wire net4428;
 wire net4429;
 wire net4430;
 wire net4431;
 wire net4432;
 wire net4433;
 wire net4434;
 wire net4435;
 wire net4436;
 wire net4437;
 wire net4438;
 wire net4439;
 wire net4440;
 wire net4441;
 wire net4442;
 wire net4443;
 wire net4444;
 wire net4445;
 wire net4446;
 wire net4447;
 wire net4448;
 wire net4449;
 wire net4450;
 wire net4451;
 wire net4452;
 wire net4453;
 wire net4454;
 wire net4455;
 wire net4456;
 wire net4457;
 wire net4458;
 wire net4459;
 wire net4460;
 wire net4461;
 wire net4462;
 wire net4463;
 wire net4464;
 wire net4465;
 wire net4466;
 wire net4467;
 wire net4468;
 wire net4469;
 wire net4470;
 wire net4471;
 wire net4472;
 wire net4473;
 wire net4474;
 wire net4475;
 wire net4476;
 wire net4477;
 wire net4478;
 wire net4479;
 wire net4480;
 wire net4481;
 wire net4482;
 wire net4483;
 wire net4484;
 wire net4485;
 wire net4486;
 wire net4487;
 wire net4488;
 wire net4489;
 wire net4490;
 wire net4491;
 wire net4492;
 wire net4493;
 wire net4494;
 wire net4495;
 wire net4496;
 wire net4497;
 wire net4498;
 wire net4499;
 wire net4500;
 wire net4501;
 wire net4502;
 wire net4503;
 wire net4504;
 wire net4505;
 wire net4506;
 wire net4507;
 wire net4508;
 wire net4509;
 wire net4510;
 wire net4511;
 wire net4512;
 wire net4513;
 wire net4514;
 wire net4515;
 wire net4516;
 wire net4517;
 wire net4518;
 wire net4519;
 wire net4520;
 wire net4521;
 wire net4522;
 wire net4523;
 wire net4524;
 wire net4525;
 wire net4526;
 wire net4527;
 wire net4528;
 wire net4529;
 wire net4530;
 wire net4531;
 wire net4532;
 wire net4533;
 wire net4534;
 wire net4535;
 wire net4536;
 wire net4537;
 wire net4538;
 wire net4539;
 wire net4540;
 wire net4541;
 wire net4542;
 wire net4543;
 wire net4544;
 wire net4545;
 wire net4546;
 wire net4547;
 wire net4548;
 wire net4549;
 wire net4550;
 wire net4551;
 wire net4552;
 wire net4553;
 wire net4554;
 wire net4555;
 wire net4556;
 wire net4557;
 wire net4558;
 wire net4559;
 wire net4560;
 wire net4561;
 wire net4562;
 wire net4563;
 wire net4564;
 wire net4565;
 wire net4566;
 wire net4567;
 wire net4568;
 wire net4569;
 wire net4570;
 wire net4571;
 wire net4572;
 wire net4573;
 wire net4574;
 wire net4575;
 wire net4576;
 wire net4577;
 wire net4578;
 wire net4579;
 wire net4580;
 wire net4581;
 wire net4582;
 wire net4583;
 wire net4584;
 wire net4585;
 wire net4586;
 wire net4587;
 wire net4588;
 wire net4589;
 wire net4590;
 wire net4591;
 wire net4592;
 wire net4593;
 wire net4594;
 wire net4595;
 wire net4596;
 wire net4597;
 wire net4598;
 wire net4599;
 wire net4600;
 wire net4601;
 wire net4602;
 wire net4603;
 wire net4604;
 wire net4605;
 wire net4606;
 wire net4607;
 wire net4608;
 wire net4609;
 wire net4610;
 wire net4611;
 wire net4612;
 wire net4613;
 wire net4614;
 wire net4615;
 wire net4616;
 wire net4617;
 wire net4618;
 wire net4619;
 wire net4620;
 wire net4621;
 wire net4622;
 wire net4623;
 wire net4624;
 wire net4625;
 wire net4626;
 wire net4627;
 wire net4628;
 wire net4629;
 wire net4630;
 wire net4631;
 wire net4632;
 wire net4633;
 wire net4634;
 wire net4635;
 wire net4636;
 wire net4637;
 wire net4638;
 wire net4639;
 wire net4640;
 wire net4641;
 wire net4642;
 wire net4643;
 wire net4644;
 wire net4645;
 wire net4646;
 wire net4647;
 wire net4648;
 wire net4649;
 wire net4650;
 wire net4651;
 wire net4652;
 wire net4653;
 wire net4654;
 wire net4655;
 wire net4656;
 wire net4657;
 wire net4658;
 wire net4659;
 wire net4660;
 wire net4661;
 wire net4662;
 wire net4663;
 wire net4664;
 wire net4665;
 wire net4666;
 wire net4667;
 wire net4668;
 wire net4669;
 wire net4670;
 wire net4671;
 wire net4672;
 wire net4673;
 wire net4674;
 wire net4675;
 wire net4676;
 wire net4677;
 wire net4678;
 wire net4679;
 wire net4680;
 wire net4681;
 wire net4682;
 wire net4683;
 wire net4684;
 wire net4685;
 wire net4686;
 wire net4687;
 wire net4688;
 wire net4689;
 wire net4690;
 wire net4691;
 wire net4692;
 wire net4693;
 wire net4694;
 wire net4695;
 wire net4696;
 wire net4697;
 wire net4698;
 wire net4699;
 wire net4700;
 wire net4701;
 wire net4702;
 wire net4703;
 wire net4704;
 wire net4705;
 wire net4706;
 wire net4707;
 wire net4708;
 wire net4709;
 wire net4710;
 wire net4711;
 wire net4712;
 wire net4713;
 wire net4714;
 wire net4715;
 wire net4716;
 wire net4717;
 wire net4718;
 wire net4719;
 wire net4720;
 wire net4721;
 wire net4722;
 wire net4723;
 wire net4724;
 wire net4725;
 wire net4726;
 wire net4727;
 wire net4728;
 wire net4729;
 wire net4730;
 wire net4731;
 wire net4732;
 wire net4733;
 wire net4734;
 wire net4735;
 wire net4736;
 wire net4737;
 wire net4738;
 wire net4739;
 wire net4740;
 wire net4741;
 wire net4742;
 wire net4743;
 wire net4744;
 wire net4745;
 wire net4746;
 wire net4747;
 wire net4748;
 wire net4749;
 wire net4750;
 wire net4751;
 wire net4752;
 wire net4753;
 wire net4754;
 wire net4755;
 wire net4756;
 wire net4757;
 wire net4758;
 wire net4759;
 wire net4760;
 wire net4761;
 wire net4762;
 wire net4763;
 wire net4764;
 wire net4765;
 wire net4766;
 wire net4767;
 wire net4768;
 wire net4769;
 wire net4770;
 wire net4771;
 wire net4772;
 wire net4773;
 wire net4774;
 wire net4775;
 wire net4776;
 wire net4777;
 wire net4778;
 wire net4779;
 wire net4780;
 wire net4781;
 wire net4782;
 wire net4783;
 wire net4784;
 wire net4785;
 wire net4786;
 wire net4787;
 wire net4788;
 wire net4789;
 wire net4790;
 wire net4791;
 wire net4792;
 wire net4793;
 wire net4794;
 wire net4795;
 wire net4796;
 wire net4797;
 wire net4798;
 wire net4799;
 wire net4800;
 wire net4801;
 wire net4802;
 wire net4803;
 wire net4804;
 wire net4805;
 wire net4806;
 wire net4807;
 wire net4808;
 wire net4809;
 wire net4810;
 wire net4811;
 wire net4812;
 wire net4813;
 wire net4814;
 wire net4815;
 wire net4816;
 wire net4817;
 wire net4818;
 wire net4819;
 wire net4820;
 wire net4821;
 wire net4822;
 wire net4823;
 wire net4824;
 wire net4825;
 wire net4826;
 wire net4827;
 wire net4828;
 wire net4829;
 wire net4830;
 wire net4831;
 wire net4832;
 wire net4833;
 wire net4834;
 wire net4835;
 wire net4836;
 wire net4837;
 wire net4838;
 wire net4839;
 wire net4840;
 wire net4841;
 wire net4842;
 wire net4843;
 wire net4844;
 wire net4845;
 wire net4846;
 wire net4847;
 wire net4848;
 wire net4849;
 wire net4850;
 wire net4851;
 wire net4852;
 wire net4853;
 wire net4854;
 wire net4855;
 wire net4856;
 wire net4857;
 wire net4858;
 wire net4859;
 wire net4860;
 wire net4861;
 wire net4862;
 wire net4863;
 wire net4864;
 wire net4865;
 wire net4866;
 wire net4867;
 wire net4868;
 wire net4869;
 wire net4870;
 wire net4871;
 wire net4872;
 wire net4873;
 wire net4874;
 wire net4875;
 wire net4876;
 wire net4877;
 wire net4878;
 wire net4879;
 wire net4880;
 wire net4881;
 wire net4882;
 wire net4883;
 wire net4884;
 wire net4885;
 wire net4886;
 wire net4887;
 wire net4888;
 wire net4889;
 wire net4890;
 wire net4891;
 wire net4892;
 wire net4893;
 wire net4894;
 wire net4895;
 wire net4896;
 wire net4897;
 wire net4898;
 wire net4899;
 wire net4900;
 wire net4901;
 wire net4902;
 wire net4903;
 wire net4904;
 wire net4905;
 wire net4906;
 wire net4907;
 wire net4908;
 wire net4909;
 wire net4910;
 wire net4911;
 wire net4912;
 wire net4913;
 wire net4914;
 wire net4915;
 wire net4916;
 wire net4917;
 wire net4918;
 wire net4919;
 wire net4920;
 wire net4921;
 wire net4922;
 wire net4923;
 wire net4924;
 wire net4925;
 wire net4926;
 wire net4927;
 wire net4928;
 wire net4929;
 wire net4930;
 wire net4931;
 wire net4932;
 wire net4933;
 wire net4934;
 wire net4935;
 wire net4936;
 wire net4937;
 wire net4938;
 wire net4939;
 wire net4940;
 wire net4941;
 wire net4942;
 wire net4943;
 wire net4944;
 wire net4945;
 wire net4946;
 wire net4947;
 wire net4948;
 wire net4949;
 wire net4950;
 wire net4951;
 wire net4952;
 wire net4953;
 wire net4954;
 wire net4955;
 wire net4956;
 wire net4957;
 wire net4958;
 wire net4959;
 wire net4960;
 wire net4961;
 wire net4962;
 wire net4963;
 wire net4964;
 wire net4965;
 wire net4966;
 wire net4967;
 wire net4968;
 wire net4969;
 wire net4970;
 wire net4971;
 wire net4972;
 wire net4973;
 wire net4974;
 wire net4975;
 wire net4976;
 wire net4977;
 wire net4978;
 wire net4979;
 wire net4980;
 wire net4981;
 wire net4982;
 wire net4983;
 wire net4984;
 wire net4985;
 wire net4986;
 wire net4987;
 wire net4988;
 wire net4989;
 wire net4990;
 wire net4991;
 wire net4992;
 wire net4993;
 wire net4994;
 wire net4995;
 wire net4996;
 wire net4997;
 wire net4998;
 wire net4999;
 wire net5000;
 wire net5001;
 wire net5002;
 wire net5003;
 wire net5004;
 wire net5005;
 wire net5006;
 wire net5007;
 wire net5008;
 wire net5009;
 wire net5010;
 wire net5011;
 wire net5012;
 wire net5013;
 wire net5014;
 wire net5015;
 wire net5016;
 wire net5017;
 wire net5018;
 wire net5019;
 wire net5020;
 wire net5021;
 wire net5022;
 wire net5023;
 wire net5024;
 wire net5025;
 wire net5026;
 wire net5027;
 wire net5028;
 wire net5029;
 wire net5030;
 wire net5031;
 wire net5032;
 wire net5033;
 wire net5034;
 wire net5035;
 wire net5036;
 wire net5037;
 wire net5038;
 wire net5039;
 wire net5040;
 wire net5041;
 wire net5042;
 wire net5043;
 wire net5044;
 wire net5045;
 wire net5046;
 wire net5047;
 wire net5048;
 wire net5049;
 wire net5050;
 wire net5051;
 wire net5052;
 wire net5053;
 wire net5054;
 wire net5055;
 wire net5056;
 wire net5057;
 wire net5058;
 wire net5059;
 wire net5060;
 wire net5061;
 wire net5062;
 wire net5063;
 wire net5064;
 wire net5065;
 wire net5066;
 wire net5067;
 wire net5068;
 wire net5069;
 wire net5070;
 wire net5071;
 wire net5072;
 wire net5073;
 wire net5074;
 wire net5075;
 wire net5076;
 wire net5077;
 wire net5078;
 wire net5079;
 wire net5080;
 wire net5081;
 wire net5082;
 wire net5083;
 wire net5084;
 wire net5085;
 wire net5086;
 wire net5087;
 wire net5088;
 wire net5089;
 wire net5090;
 wire net5091;
 wire net5092;
 wire net5093;
 wire net5094;
 wire net5095;
 wire net5096;
 wire net5097;
 wire net5098;
 wire net5099;
 wire net5100;
 wire net5101;
 wire net5102;
 wire net5103;
 wire net5104;
 wire net5105;
 wire net5106;
 wire net5107;
 wire net5108;
 wire net5109;
 wire net5110;
 wire net5111;
 wire net5112;
 wire net5113;
 wire net5114;
 wire net5115;
 wire net5116;
 wire net5117;
 wire net5118;
 wire net5119;
 wire net5120;
 wire net5121;
 wire net5122;
 wire net5123;
 wire net5124;
 wire net5125;
 wire net5126;
 wire net5127;
 wire net5128;
 wire net5129;
 wire net5130;
 wire net5131;
 wire net5132;
 wire net5133;
 wire net5134;
 wire net5135;
 wire net5136;
 wire net5137;
 wire net5138;
 wire net5139;
 wire net5140;
 wire net5141;
 wire net5142;
 wire net5143;
 wire net5144;
 wire net5145;
 wire net5146;
 wire net5147;
 wire net5148;
 wire net5149;
 wire net5150;
 wire net5151;
 wire net5152;
 wire net5153;
 wire net5154;
 wire net5155;
 wire net5156;
 wire net5157;
 wire net5158;
 wire net5159;
 wire net5160;
 wire net5161;
 wire net5162;
 wire net5163;
 wire net5164;
 wire net5165;
 wire net5166;
 wire net5167;
 wire net5168;
 wire net5169;
 wire net5170;
 wire net5171;
 wire net5172;
 wire net5173;
 wire net5174;
 wire net5175;
 wire net5176;
 wire net5177;
 wire net5178;
 wire net5179;
 wire net5180;
 wire net5181;
 wire net5182;
 wire net5183;
 wire net5184;
 wire net5185;
 wire net5186;
 wire net5187;
 wire net5188;
 wire net5189;
 wire net5190;
 wire net5191;
 wire net5192;
 wire net5193;
 wire net5194;
 wire net5195;
 wire net5196;
 wire net5197;
 wire net5198;
 wire net5199;
 wire net5200;
 wire net5201;
 wire net5202;
 wire net5203;
 wire net5204;
 wire net5205;
 wire net5206;
 wire net5207;
 wire net5208;
 wire net5209;
 wire net5210;
 wire net5211;
 wire net5212;
 wire net5213;
 wire net5214;
 wire net5215;
 wire net5216;
 wire net5217;
 wire net5218;
 wire net5219;
 wire net5220;
 wire net5221;
 wire net5222;
 wire net5223;
 wire net5224;
 wire net5225;
 wire net5226;
 wire net5227;
 wire net5228;
 wire net5229;
 wire net5230;
 wire net5231;
 wire net5232;
 wire net5233;
 wire net5234;
 wire net5235;
 wire net5236;
 wire net5237;
 wire net5238;
 wire net5239;
 wire net5240;
 wire net5241;
 wire net5242;
 wire net5243;
 wire net5244;
 wire net5245;
 wire net5246;
 wire net5247;
 wire net5248;
 wire net5249;
 wire net5250;
 wire net5251;
 wire net5252;
 wire net5253;
 wire net5254;
 wire net5255;
 wire net5256;
 wire net5257;
 wire net5258;
 wire net5259;
 wire net5260;
 wire net5261;
 wire net5262;
 wire net5263;
 wire net5264;
 wire net5265;
 wire net5266;
 wire net5267;
 wire net5268;
 wire net5269;
 wire net5270;
 wire net5271;
 wire net5272;
 wire net5273;
 wire net5274;
 wire net5275;
 wire net5276;
 wire net5277;
 wire net5278;
 wire net5279;
 wire net5280;
 wire net5281;
 wire net5282;
 wire net5283;
 wire net5284;
 wire net5285;
 wire net5286;
 wire net5287;
 wire net5288;
 wire net5289;
 wire net5290;
 wire net5291;
 wire net5292;
 wire net5293;
 wire net5294;
 wire net5295;
 wire net5296;
 wire net5297;
 wire net5298;
 wire net5299;
 wire net5300;
 wire net5301;
 wire net5302;
 wire net5303;
 wire net5304;
 wire net5305;
 wire net5306;
 wire net5307;
 wire net5308;
 wire net5309;
 wire net5310;
 wire net5311;
 wire net5312;
 wire net5313;
 wire net5314;
 wire net5315;
 wire net5316;
 wire net5317;
 wire net5318;
 wire net5319;
 wire net5320;
 wire net5321;
 wire net5322;
 wire net5323;
 wire net5324;
 wire net5325;
 wire net5326;
 wire net5327;
 wire net5328;
 wire net5329;
 wire net5330;
 wire net5331;
 wire net5332;
 wire net5333;
 wire net5334;
 wire net5335;
 wire net5336;
 wire net5337;
 wire net5338;
 wire net5339;
 wire net5340;
 wire net5341;
 wire net5342;
 wire net5343;
 wire net5344;
 wire net5345;
 wire net5346;
 wire net5347;
 wire net5348;
 wire net5349;
 wire net5350;
 wire net5351;
 wire net5352;
 wire net5353;
 wire net5354;
 wire net5355;
 wire net5356;
 wire net5357;
 wire net5358;
 wire net5359;
 wire net5360;
 wire net5361;
 wire net5362;
 wire net5363;
 wire net5364;
 wire net5365;
 wire net5366;
 wire net5367;
 wire net5368;
 wire net5369;
 wire net5370;
 wire net5371;
 wire net5372;
 wire net5373;
 wire net5374;
 wire net5375;
 wire net5376;
 wire net5377;
 wire net5378;
 wire net5379;
 wire net5380;
 wire net5381;
 wire net5382;
 wire net5383;
 wire net5384;
 wire net5385;
 wire net5386;
 wire net5387;
 wire net5388;
 wire net5389;
 wire net5390;
 wire net5391;
 wire net5392;
 wire net5393;
 wire net5394;
 wire net5395;
 wire net5396;
 wire net5397;
 wire net5398;
 wire net5399;
 wire net5400;
 wire net5401;
 wire net5402;
 wire net5403;
 wire net5404;
 wire net5405;
 wire net5406;
 wire net5407;
 wire net5408;
 wire net5409;
 wire net5410;
 wire net5411;
 wire net5412;
 wire net5413;
 wire net5414;
 wire net5415;
 wire net5416;
 wire net5417;
 wire net5418;
 wire net5419;
 wire net5420;
 wire net5421;
 wire net5422;
 wire net5423;
 wire net5424;
 wire net5425;
 wire net5426;
 wire net5427;
 wire net5428;
 wire net5429;
 wire net5430;
 wire net5431;
 wire net5432;
 wire net5433;
 wire net5434;
 wire net5435;
 wire net5436;
 wire net5437;
 wire net5438;
 wire net5439;
 wire net5440;
 wire net5441;
 wire net5442;
 wire net5443;
 wire net5444;
 wire net5445;
 wire net5446;
 wire net5447;
 wire net5448;
 wire net5449;
 wire net5450;
 wire net5451;
 wire net5452;
 wire net5453;
 wire net5454;
 wire net5455;
 wire net5456;
 wire net5457;
 wire net5458;
 wire net5459;
 wire net5460;
 wire net5461;
 wire net5462;
 wire net5463;
 wire net5464;
 wire net5465;
 wire net5466;
 wire net5467;
 wire net5468;
 wire net5469;
 wire net5470;
 wire net5471;
 wire net5472;
 wire net5473;
 wire net5474;
 wire net5475;
 wire net5476;
 wire net5477;
 wire net5478;
 wire net5479;
 wire net5480;
 wire net5481;
 wire net5482;
 wire net5483;
 wire net5484;
 wire net5485;
 wire net5486;
 wire net5487;
 wire net5488;
 wire net5489;
 wire net5490;
 wire net5491;
 wire net5492;
 wire net5493;
 wire net5494;
 wire net5495;
 wire net5496;
 wire net5497;
 wire net5498;
 wire net5499;
 wire net5500;
 wire net5501;
 wire net5502;
 wire net5503;
 wire net5504;
 wire net5505;
 wire net5506;
 wire net5507;
 wire net5508;
 wire net5509;
 wire net5510;
 wire net5511;
 wire net5512;
 wire net5513;
 wire net5514;
 wire net5515;
 wire net5516;
 wire net5517;
 wire net5518;
 wire net5519;
 wire net5520;
 wire net5521;
 wire net5522;
 wire net5523;
 wire net5524;
 wire net5525;
 wire net5526;
 wire net5527;
 wire net5528;
 wire net5529;
 wire net5530;
 wire net5531;
 wire net5532;
 wire net5533;
 wire net5534;
 wire net5535;
 wire net5536;
 wire net5537;
 wire net5538;
 wire net5539;
 wire net5540;
 wire net5541;
 wire net5542;
 wire net5543;
 wire net5544;
 wire net5545;
 wire net5546;
 wire net5547;
 wire net5548;
 wire net5549;
 wire net5550;
 wire net5551;
 wire net5552;
 wire net5553;
 wire net5554;
 wire net5555;
 wire net5556;
 wire net5557;
 wire net5558;
 wire net5559;
 wire net5560;
 wire net5561;
 wire net5562;
 wire net5563;
 wire net5564;
 wire net5565;
 wire net5566;
 wire net5567;
 wire net5568;
 wire net5569;
 wire net5570;
 wire net5571;
 wire net5572;
 wire net5573;
 wire net5574;
 wire net5575;
 wire net5576;
 wire net5577;
 wire net5578;
 wire net5579;
 wire net5580;

 sg13g2_inv_1 _19337_ (.Y(_10375_),
    .A(net5462));
 sg13g2_inv_1 _19338_ (.Y(_10376_),
    .A(\soc_I.qqspi_I.spi_buf[24] ));
 sg13g2_inv_1 _19339_ (.Y(_10377_),
    .A(sclk));
 sg13g2_inv_1 _19340_ (.Y(_10378_),
    .A(net3705));
 sg13g2_inv_1 _19341_ (.Y(_10379_),
    .A(net4645));
 sg13g2_inv_1 _19342_ (.Y(_10380_),
    .A(net4102));
 sg13g2_inv_1 _19343_ (.Y(_10381_),
    .A(net4008));
 sg13g2_inv_1 _19344_ (.Y(_10382_),
    .A(net4316));
 sg13g2_inv_1 _19345_ (.Y(_10383_),
    .A(net3947));
 sg13g2_inv_1 _19346_ (.Y(_10384_),
    .A(net3719));
 sg13g2_inv_1 _19347_ (.Y(_10385_),
    .A(\soc_I.spi0_I.spi_buf[0] ));
 sg13g2_inv_1 _19348_ (.Y(_10386_),
    .A(\soc_I.tx_uart_i.tx_data_reg[6] ));
 sg13g2_inv_1 _19349_ (.Y(_10387_),
    .A(net2608));
 sg13g2_inv_2 _19350_ (.Y(_10388_),
    .A(\soc_I.tx_uart_i.ready ));
 sg13g2_inv_1 _19351_ (.Y(_10389_),
    .A(net3147));
 sg13g2_inv_1 _19352_ (.Y(_10390_),
    .A(net2606));
 sg13g2_inv_1 _19353_ (.Y(_10391_),
    .A(\soc_I.rx_uart_i.fifo_i.wr_ptr[1] ));
 sg13g2_inv_1 _19354_ (.Y(_10392_),
    .A(net2604));
 sg13g2_inv_1 _19355_ (.Y(_10393_),
    .A(net4545));
 sg13g2_inv_1 _19356_ (.Y(_10394_),
    .A(net3095));
 sg13g2_inv_1 _19357_ (.Y(_10395_),
    .A(net3400));
 sg13g2_inv_2 _19358_ (.Y(_10396_),
    .A(\soc_I.rx_uart_i.fifo_i.din[0] ));
 sg13g2_inv_1 _19359_ (.Y(_10397_),
    .A(net5215));
 sg13g2_inv_1 _19360_ (.Y(_10398_),
    .A(net2839));
 sg13g2_inv_1 _19361_ (.Y(_10399_),
    .A(net4776));
 sg13g2_inv_2 _19362_ (.Y(_10400_),
    .A(net4564));
 sg13g2_inv_1 _19363_ (.Y(_10401_),
    .A(\soc_I.clint_I.mtime[61] ));
 sg13g2_inv_1 _19364_ (.Y(_10402_),
    .A(\soc_I.clint_I.mtime[60] ));
 sg13g2_inv_1 _19365_ (.Y(_10403_),
    .A(\soc_I.clint_I.mtime[59] ));
 sg13g2_inv_1 _19366_ (.Y(_10404_),
    .A(net4268));
 sg13g2_inv_1 _19367_ (.Y(_10405_),
    .A(net5113));
 sg13g2_inv_1 _19368_ (.Y(_10406_),
    .A(net4274));
 sg13g2_inv_1 _19369_ (.Y(_10407_),
    .A(net4946));
 sg13g2_inv_1 _19370_ (.Y(_10408_),
    .A(\soc_I.clint_I.mtime[52] ));
 sg13g2_inv_1 _19371_ (.Y(_10409_),
    .A(\soc_I.clint_I.mtime[48] ));
 sg13g2_inv_2 _19372_ (.Y(_10410_),
    .A(net4001));
 sg13g2_inv_1 _19373_ (.Y(_10411_),
    .A(net5552));
 sg13g2_inv_2 _19374_ (.Y(_10412_),
    .A(net5498));
 sg13g2_inv_1 _19375_ (.Y(_10413_),
    .A(\soc_I.clint_I.mtime[44] ));
 sg13g2_inv_1 _19376_ (.Y(_10414_),
    .A(\soc_I.clint_I.mtime[39] ));
 sg13g2_inv_2 _19377_ (.Y(_10415_),
    .A(net5482));
 sg13g2_inv_1 _19378_ (.Y(_10416_),
    .A(net5166));
 sg13g2_inv_1 _19379_ (.Y(_10417_),
    .A(net5546));
 sg13g2_inv_1 _19380_ (.Y(_10418_),
    .A(\soc_I.clint_I.mtime[35] ));
 sg13g2_inv_1 _19381_ (.Y(_10419_),
    .A(\soc_I.clint_I.mtime[34] ));
 sg13g2_inv_1 _19382_ (.Y(_10420_),
    .A(net4996));
 sg13g2_inv_1 _19383_ (.Y(_10421_),
    .A(net5509));
 sg13g2_inv_1 _19384_ (.Y(_10422_),
    .A(\soc_I.clint_I.mtime[30] ));
 sg13g2_inv_1 _19385_ (.Y(_10423_),
    .A(net4555));
 sg13g2_inv_1 _19386_ (.Y(_10424_),
    .A(net5194));
 sg13g2_inv_1 _19387_ (.Y(_10425_),
    .A(\soc_I.clint_I.mtime[25] ));
 sg13g2_inv_2 _19388_ (.Y(_10426_),
    .A(net5297));
 sg13g2_inv_1 _19389_ (.Y(_10427_),
    .A(\soc_I.clint_I.mtime[23] ));
 sg13g2_inv_1 _19390_ (.Y(_10428_),
    .A(net5119));
 sg13g2_inv_1 _19391_ (.Y(_10429_),
    .A(\soc_I.clint_I.mtime[19] ));
 sg13g2_inv_2 _19392_ (.Y(_10430_),
    .A(net5390));
 sg13g2_inv_1 _19393_ (.Y(_10431_),
    .A(\soc_I.clint_I.mtime[17] ));
 sg13g2_inv_1 _19394_ (.Y(_10432_),
    .A(\soc_I.clint_I.mtime[15] ));
 sg13g2_inv_1 _19395_ (.Y(_10433_),
    .A(net5243));
 sg13g2_inv_1 _19396_ (.Y(_10434_),
    .A(\soc_I.clint_I.mtime[13] ));
 sg13g2_inv_1 _19397_ (.Y(_10435_),
    .A(\soc_I.clint_I.mtime[11] ));
 sg13g2_inv_1 _19398_ (.Y(_10436_),
    .A(\soc_I.clint_I.mtime[10] ));
 sg13g2_inv_1 _19399_ (.Y(_10437_),
    .A(\soc_I.clint_I.mtime[9] ));
 sg13g2_inv_1 _19400_ (.Y(_10438_),
    .A(net5087));
 sg13g2_inv_1 _19401_ (.Y(_10439_),
    .A(\soc_I.clint_I.mtime[7] ));
 sg13g2_inv_1 _19402_ (.Y(_10440_),
    .A(net3799));
 sg13g2_inv_1 _19403_ (.Y(_10441_),
    .A(net3593));
 sg13g2_inv_2 _19404_ (.Y(_10442_),
    .A(net4489));
 sg13g2_inv_1 _19405_ (.Y(_10443_),
    .A(\soc_I.clint_I.mtime[3] ));
 sg13g2_inv_1 _19406_ (.Y(_10444_),
    .A(\soc_I.clint_I.mtime[1] ));
 sg13g2_inv_1 _19407_ (.Y(_10445_),
    .A(\soc_I.clint_I.mtime[0] ));
 sg13g2_inv_1 _19408_ (.Y(_10446_),
    .A(\soc_I.clint_I.mtimecmp[36] ));
 sg13g2_inv_1 _19409_ (.Y(_10447_),
    .A(\soc_I.clint_I.mtimecmp[35] ));
 sg13g2_inv_1 _19410_ (.Y(_10448_),
    .A(\soc_I.clint_I.mtimecmp[34] ));
 sg13g2_inv_1 _19411_ (.Y(_10449_),
    .A(\soc_I.clint_I.mtimecmp[33] ));
 sg13g2_inv_1 _19412_ (.Y(_10450_),
    .A(net4981));
 sg13g2_inv_1 _19413_ (.Y(_10451_),
    .A(net4242));
 sg13g2_inv_1 _19414_ (.Y(_10452_),
    .A(net4353));
 sg13g2_inv_1 _19415_ (.Y(_10453_),
    .A(\soc_I.PC[20] ));
 sg13g2_inv_2 _19416_ (.Y(_10454_),
    .A(net5308));
 sg13g2_inv_2 _19417_ (.Y(_10455_),
    .A(net5370));
 sg13g2_inv_2 _19418_ (.Y(_10456_),
    .A(net5211));
 sg13g2_inv_2 _19419_ (.Y(_10457_),
    .A(net5226));
 sg13g2_inv_1 _19420_ (.Y(_10458_),
    .A(net9431));
 sg13g2_inv_4 _19421_ (.A(net9499),
    .Y(_10459_));
 sg13g2_inv_4 _19422_ (.A(net9537),
    .Y(_10460_));
 sg13g2_inv_8 _19423_ (.Y(_10461_),
    .A(net9550));
 sg13g2_inv_8 _19424_ (.Y(_10462_),
    .A(net9555));
 sg13g2_inv_8 _19425_ (.Y(_10463_),
    .A(net9573));
 sg13g2_inv_8 _19426_ (.Y(_10464_),
    .A(net9684));
 sg13g2_inv_2 _19427_ (.Y(_10465_),
    .A(net9705));
 sg13g2_inv_1 _19428_ (.Y(_10466_),
    .A(net9709));
 sg13g2_inv_1 _19429_ (.Y(_10467_),
    .A(\soc_I.kianv_I.Instr[8] ));
 sg13g2_inv_1 _19430_ (.Y(_10468_),
    .A(net5557));
 sg13g2_inv_1 _19431_ (.Y(_10469_),
    .A(net9715));
 sg13g2_inv_1 _19432_ (.Y(_10470_),
    .A(\soc_I.kianv_I.Instr[2] ));
 sg13g2_inv_1 _19433_ (.Y(_10471_),
    .A(net4118));
 sg13g2_inv_1 _19434_ (.Y(_10472_),
    .A(net4300));
 sg13g2_inv_2 _19435_ (.Y(_10473_),
    .A(net5024));
 sg13g2_inv_1 _19436_ (.Y(_10474_),
    .A(net4783));
 sg13g2_inv_1 _19437_ (.Y(_10475_),
    .A(net5089));
 sg13g2_inv_1 _19438_ (.Y(_10476_),
    .A(net5311));
 sg13g2_inv_1 _19439_ (.Y(_10477_),
    .A(net5152));
 sg13g2_inv_1 _19440_ (.Y(_10478_),
    .A(net4588));
 sg13g2_inv_1 _19441_ (.Y(_10479_),
    .A(net5127));
 sg13g2_inv_1 _19442_ (.Y(_10480_),
    .A(net4785));
 sg13g2_inv_1 _19443_ (.Y(_10481_),
    .A(net4226));
 sg13g2_inv_1 _19444_ (.Y(_10482_),
    .A(net5063));
 sg13g2_inv_1 _19445_ (.Y(_10483_),
    .A(net5541));
 sg13g2_inv_1 _19446_ (.Y(_10484_),
    .A(net5439));
 sg13g2_inv_1 _19447_ (.Y(_10485_),
    .A(net4330));
 sg13g2_inv_1 _19448_ (.Y(_10486_),
    .A(net4797));
 sg13g2_inv_1 _19449_ (.Y(_10487_),
    .A(net5450));
 sg13g2_inv_1 _19450_ (.Y(_10488_),
    .A(net5328));
 sg13g2_inv_1 _19451_ (.Y(_10489_),
    .A(net4526));
 sg13g2_inv_1 _19452_ (.Y(_10490_),
    .A(net5157));
 sg13g2_inv_1 _19453_ (.Y(_10491_),
    .A(net5241));
 sg13g2_inv_2 _19454_ (.Y(_10492_),
    .A(net4972));
 sg13g2_inv_1 _19455_ (.Y(_10493_),
    .A(net4452));
 sg13g2_inv_2 _19456_ (.Y(_10494_),
    .A(net4590));
 sg13g2_inv_1 _19457_ (.Y(_10495_),
    .A(net4541));
 sg13g2_inv_1 _19458_ (.Y(_10496_),
    .A(net3999));
 sg13g2_inv_1 _19459_ (.Y(_10497_),
    .A(net2664));
 sg13g2_inv_1 _19460_ (.Y(_10498_),
    .A(net2726));
 sg13g2_inv_1 _19461_ (.Y(_10499_),
    .A(net2755));
 sg13g2_inv_1 _19462_ (.Y(_10500_),
    .A(net2683));
 sg13g2_inv_1 _19463_ (.Y(_10501_),
    .A(net4188));
 sg13g2_inv_1 _19464_ (.Y(_10502_),
    .A(net2815));
 sg13g2_inv_1 _19465_ (.Y(_10503_),
    .A(net2854));
 sg13g2_inv_1 _19466_ (.Y(_10504_),
    .A(net2736));
 sg13g2_inv_1 _19467_ (.Y(_10505_),
    .A(net2663));
 sg13g2_inv_1 _19468_ (.Y(_10506_),
    .A(net2751));
 sg13g2_inv_1 _19469_ (.Y(_10507_),
    .A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[31] ));
 sg13g2_inv_1 _19470_ (.Y(_10508_),
    .A(net9222));
 sg13g2_inv_1 _19471_ (.Y(_10509_),
    .A(net9722));
 sg13g2_inv_1 _19472_ (.Y(_10510_),
    .A(net9734));
 sg13g2_inv_1 _19473_ (.Y(_10511_),
    .A(net9743));
 sg13g2_inv_1 _19474_ (.Y(_10512_),
    .A(net9756));
 sg13g2_inv_1 _19475_ (.Y(_10513_),
    .A(net9237));
 sg13g2_inv_1 _19476_ (.Y(_10514_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[30] ));
 sg13g2_inv_2 _19477_ (.Y(_10515_),
    .A(net3964));
 sg13g2_inv_2 _19478_ (.Y(_10516_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[1] ));
 sg13g2_inv_2 _19479_ (.Y(_10517_),
    .A(net4684));
 sg13g2_inv_1 _19480_ (.Y(_10518_),
    .A(net4028));
 sg13g2_inv_1 _19481_ (.Y(_10519_),
    .A(net3193));
 sg13g2_inv_1 _19482_ (.Y(_10520_),
    .A(net5363));
 sg13g2_inv_1 _19483_ (.Y(_10521_),
    .A(net5086));
 sg13g2_inv_1 _19484_ (.Y(_10522_),
    .A(net5034));
 sg13g2_inv_1 _19485_ (.Y(_10523_),
    .A(net4511));
 sg13g2_inv_1 _19486_ (.Y(_10524_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[55] ));
 sg13g2_inv_1 _19487_ (.Y(_10525_),
    .A(net4647));
 sg13g2_inv_1 _19488_ (.Y(_10526_),
    .A(net5549));
 sg13g2_inv_1 _19489_ (.Y(_10527_),
    .A(net5093));
 sg13g2_inv_1 _19490_ (.Y(_10528_),
    .A(net5481));
 sg13g2_inv_1 _19491_ (.Y(_10529_),
    .A(net5489));
 sg13g2_inv_1 _19492_ (.Y(_10530_),
    .A(net3791));
 sg13g2_inv_1 _19493_ (.Y(_10531_),
    .A(net4058));
 sg13g2_inv_1 _19494_ (.Y(_10532_),
    .A(net5344));
 sg13g2_inv_2 _19495_ (.Y(_10533_),
    .A(net5453));
 sg13g2_inv_1 _19496_ (.Y(_10534_),
    .A(net5199));
 sg13g2_inv_1 _19497_ (.Y(_10535_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[36] ));
 sg13g2_inv_1 _19498_ (.Y(_10536_),
    .A(net5314));
 sg13g2_inv_1 _19499_ (.Y(_10537_),
    .A(net5341));
 sg13g2_inv_1 _19500_ (.Y(_10538_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[32] ));
 sg13g2_inv_1 _19501_ (.Y(_10539_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[31] ));
 sg13g2_inv_1 _19502_ (.Y(_10540_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[30] ));
 sg13g2_inv_1 _19503_ (.Y(_10541_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[27] ));
 sg13g2_inv_1 _19504_ (.Y(_10542_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[23] ));
 sg13g2_inv_1 _19505_ (.Y(_10543_),
    .A(net5524));
 sg13g2_inv_1 _19506_ (.Y(_10544_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[13] ));
 sg13g2_inv_1 _19507_ (.Y(_10545_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[12] ));
 sg13g2_inv_1 _19508_ (.Y(_10546_),
    .A(net5346));
 sg13g2_inv_1 _19509_ (.Y(_10547_),
    .A(net3098));
 sg13g2_inv_1 _19510_ (.Y(_10548_),
    .A(net4920));
 sg13g2_inv_1 _19511_ (.Y(_10549_),
    .A(net5495));
 sg13g2_inv_1 _19512_ (.Y(_10550_),
    .A(net5540));
 sg13g2_inv_1 _19513_ (.Y(_10551_),
    .A(net5366));
 sg13g2_inv_1 _19514_ (.Y(_10552_),
    .A(net4129));
 sg13g2_inv_1 _19515_ (.Y(_10553_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[0] ));
 sg13g2_inv_1 _19516_ (.Y(_10554_),
    .A(net4221));
 sg13g2_inv_1 _19517_ (.Y(_10555_),
    .A(net4144));
 sg13g2_inv_1 _19518_ (.Y(_10556_),
    .A(net4477));
 sg13g2_inv_1 _19519_ (.Y(_10557_),
    .A(net4704));
 sg13g2_inv_1 _19520_ (.Y(_10558_),
    .A(\soc_I.clint_I.mtimecmp[31] ));
 sg13g2_inv_1 _19521_ (.Y(_10559_),
    .A(\soc_I.clint_I.mtimecmp[30] ));
 sg13g2_inv_1 _19522_ (.Y(_10560_),
    .A(\soc_I.clint_I.mtimecmp[29] ));
 sg13g2_inv_2 _19523_ (.Y(_10561_),
    .A(net5295));
 sg13g2_inv_1 _19524_ (.Y(_10562_),
    .A(\soc_I.clint_I.mtimecmp[22] ));
 sg13g2_inv_1 _19525_ (.Y(_10563_),
    .A(\soc_I.clint_I.mtimecmp[21] ));
 sg13g2_inv_1 _19526_ (.Y(_10564_),
    .A(\soc_I.clint_I.mtimecmp[20] ));
 sg13g2_inv_1 _19527_ (.Y(_10565_),
    .A(\soc_I.clint_I.mtimecmp[13] ));
 sg13g2_inv_1 _19528_ (.Y(_10566_),
    .A(\soc_I.clint_I.mtimecmp[12] ));
 sg13g2_inv_1 _19529_ (.Y(_10567_),
    .A(\soc_I.clint_I.mtimecmp[11] ));
 sg13g2_inv_1 _19530_ (.Y(_10568_),
    .A(\soc_I.clint_I.mtimecmp[10] ));
 sg13g2_inv_1 _19531_ (.Y(_10569_),
    .A(\soc_I.clint_I.mtimecmp[9] ));
 sg13g2_inv_1 _19532_ (.Y(_10570_),
    .A(\soc_I.clint_I.mtimecmp[8] ));
 sg13g2_inv_1 _19533_ (.Y(_10571_),
    .A(net4856));
 sg13g2_inv_1 _19534_ (.Y(_10572_),
    .A(\soc_I.clint_I.mtimecmp[63] ));
 sg13g2_inv_1 _19535_ (.Y(_10573_),
    .A(\soc_I.clint_I.mtimecmp[59] ));
 sg13g2_inv_1 _19536_ (.Y(_10574_),
    .A(\soc_I.clint_I.mtimecmp[58] ));
 sg13g2_inv_1 _19537_ (.Y(_10575_),
    .A(\soc_I.clint_I.mtimecmp[57] ));
 sg13g2_inv_1 _19538_ (.Y(_10576_),
    .A(\soc_I.clint_I.mtimecmp[56] ));
 sg13g2_inv_1 _19539_ (.Y(_10577_),
    .A(\soc_I.clint_I.mtimecmp[54] ));
 sg13g2_inv_1 _19540_ (.Y(_10578_),
    .A(\soc_I.clint_I.mtimecmp[53] ));
 sg13g2_inv_1 _19541_ (.Y(_10579_),
    .A(\soc_I.clint_I.mtimecmp[49] ));
 sg13g2_inv_1 _19542_ (.Y(_10580_),
    .A(\soc_I.clint_I.mtimecmp[48] ));
 sg13g2_inv_1 _19543_ (.Y(_10581_),
    .A(\soc_I.clint_I.mtimecmp[46] ));
 sg13g2_inv_1 _19544_ (.Y(_10582_),
    .A(\soc_I.clint_I.mtimecmp[45] ));
 sg13g2_inv_1 _19545_ (.Y(_10583_),
    .A(\soc_I.clint_I.mtimecmp[43] ));
 sg13g2_inv_1 _19546_ (.Y(_10584_),
    .A(\soc_I.clint_I.mtimecmp[42] ));
 sg13g2_inv_1 _19547_ (.Y(_10585_),
    .A(\soc_I.clint_I.mtimecmp[41] ));
 sg13g2_inv_1 _19548_ (.Y(_10586_),
    .A(\soc_I.clint_I.mtimecmp[40] ));
 sg13g2_inv_1 _19549_ (.Y(_10587_),
    .A(_00188_));
 sg13g2_inv_1 _19550_ (.Y(_10588_),
    .A(_00189_));
 sg13g2_inv_1 _19551_ (.Y(_10589_),
    .A(\soc_I.tx_uart_i.wait_states[0] ));
 sg13g2_inv_1 _19552_ (.Y(_10590_),
    .A(_00216_));
 sg13g2_inv_1 _19553_ (.Y(_10591_),
    .A(\soc_I.kianv_I.datapath_unit_I.A2[16] ));
 sg13g2_inv_1 _19554_ (.Y(_10592_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.div_state[0] ));
 sg13g2_inv_1 _19555_ (.Y(_10593_),
    .A(net9342));
 sg13g2_inv_2 _19556_ (.Y(_10594_),
    .A(\soc_I.qqspi_I.state[5] ));
 sg13g2_inv_1 _19557_ (.Y(_10595_),
    .A(_00242_));
 sg13g2_inv_4 _19558_ (.A(_00244_),
    .Y(_10596_));
 sg13g2_inv_1 _19559_ (.Y(_10597_),
    .A(_00246_));
 sg13g2_inv_1 _19560_ (.Y(_10598_),
    .A(_00247_));
 sg13g2_inv_1 _19561_ (.Y(_10599_),
    .A(_00248_));
 sg13g2_inv_1 _19562_ (.Y(_10600_),
    .A(\soc_I.clint_I.tick_cnt[12] ));
 sg13g2_inv_1 _19563_ (.Y(_10601_),
    .A(\soc_I.clint_I.tick_cnt[15] ));
 sg13g2_inv_2 _19564_ (.Y(_10602_),
    .A(net9296));
 sg13g2_inv_1 _19565_ (.Y(_10603_),
    .A(net9254));
 sg13g2_inv_4 _19566_ (.A(\soc_I.spi_div_ready ),
    .Y(_10604_));
 sg13g2_inv_2 _19567_ (.Y(_10605_),
    .A(net9291));
 sg13g2_inv_2 _19568_ (.Y(_10606_),
    .A(net9212));
 sg13g2_inv_1 _19569_ (.Y(_10607_),
    .A(net9716));
 sg13g2_inv_1 _19570_ (.Y(_10608_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[4] ));
 sg13g2_inv_1 _19571_ (.Y(_10609_),
    .A(net4039));
 sg13g2_inv_1 _19572_ (.Y(_10610_),
    .A(net3993));
 sg13g2_inv_1 _19573_ (.Y(_10611_),
    .A(net3219));
 sg13g2_inv_1 _19574_ (.Y(_10612_),
    .A(net3374));
 sg13g2_inv_1 _19575_ (.Y(_10613_),
    .A(net3236));
 sg13g2_inv_1 _19576_ (.Y(_10614_),
    .A(net3643));
 sg13g2_inv_1 _19577_ (.Y(_10615_),
    .A(net4808));
 sg13g2_inv_1 _19578_ (.Y(_10616_),
    .A(net4948));
 sg13g2_inv_1 _19579_ (.Y(_10617_),
    .A(net3673));
 sg13g2_inv_1 _19580_ (.Y(_10618_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[0] ));
 sg13g2_inv_1 _19581_ (.Y(_10619_),
    .A(net5066));
 sg13g2_inv_1 _19582_ (.Y(_10620_),
    .A(net5201));
 sg13g2_inv_1 _19583_ (.Y(_10621_),
    .A(net5214));
 sg13g2_inv_1 _19584_ (.Y(_10622_),
    .A(net5069));
 sg13g2_inv_1 _19585_ (.Y(_10623_),
    .A(net4713));
 sg13g2_inv_1 _19586_ (.Y(_10624_),
    .A(net4929));
 sg13g2_inv_1 _19587_ (.Y(_10625_),
    .A(net5083));
 sg13g2_inv_1 _19588_ (.Y(_10626_),
    .A(net5425));
 sg13g2_inv_1 _19589_ (.Y(_10627_),
    .A(net5236));
 sg13g2_inv_1 _19590_ (.Y(_10628_),
    .A(net5264));
 sg13g2_inv_1 _19591_ (.Y(_10629_),
    .A(net5396));
 sg13g2_inv_1 _19592_ (.Y(_10630_),
    .A(net5350));
 sg13g2_inv_1 _19593_ (.Y(_10631_),
    .A(net5378));
 sg13g2_inv_2 _19594_ (.Y(_10632_),
    .A(net5427));
 sg13g2_inv_1 _19595_ (.Y(_10633_),
    .A(net4068));
 sg13g2_inv_2 _19596_ (.Y(_10634_),
    .A(net5335));
 sg13g2_inv_1 _19597_ (.Y(_10635_),
    .A(net5431));
 sg13g2_inv_1 _19598_ (.Y(_10636_),
    .A(net5554));
 sg13g2_inv_1 _19599_ (.Y(_10637_),
    .A(net5533));
 sg13g2_inv_1 _19600_ (.Y(_10638_),
    .A(net5340));
 sg13g2_inv_1 _19601_ (.Y(_10639_),
    .A(net5401));
 sg13g2_inv_1 _19602_ (.Y(_10640_),
    .A(net5408));
 sg13g2_inv_1 _19603_ (.Y(_10641_),
    .A(net5357));
 sg13g2_inv_1 _19604_ (.Y(_10642_),
    .A(net5111));
 sg13g2_inv_1 _19605_ (.Y(_10643_),
    .A(net5132));
 sg13g2_inv_1 _19606_ (.Y(_10644_),
    .A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mip[7] ));
 sg13g2_inv_1 _19607_ (.Y(_10645_),
    .A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mip[3] ));
 sg13g2_inv_1 _19608_ (.Y(_10646_),
    .A(\soc_I.kianv_I.datapath_unit_I.ADDR_I.q[0] ));
 sg13g2_inv_2 _19609_ (.Y(_10647_),
    .A(net9422));
 sg13g2_inv_1 _19610_ (.Y(_10648_),
    .A(net4426));
 sg13g2_inv_1 _19611_ (.Y(_10649_),
    .A(net4259));
 sg13g2_inv_1 _19612_ (.Y(_10650_),
    .A(\soc_I.rx_uart_i.fifo_i.cnt[2] ));
 sg13g2_inv_1 _19613_ (.Y(_10651_),
    .A(net5293));
 sg13g2_inv_1 _19614_ (.Y(_10652_),
    .A(net5265));
 sg13g2_inv_1 _19615_ (.Y(_10653_),
    .A(net3670));
 sg13g2_inv_1 _19616_ (.Y(_10654_),
    .A(_00014_));
 sg13g2_inv_1 _19617_ (.Y(_10655_),
    .A(_00017_));
 sg13g2_inv_1 _19618_ (.Y(_10656_),
    .A(net3092));
 sg13g2_inv_1 _19619_ (.Y(_10657_),
    .A(_00021_));
 sg13g2_inv_1 _19620_ (.Y(_10658_),
    .A(_00025_));
 sg13g2_inv_1 _19621_ (.Y(_10659_),
    .A(_00030_));
 sg13g2_inv_1 _19622_ (.Y(_10660_),
    .A(_00037_));
 sg13g2_inv_1 _19623_ (.Y(_10661_),
    .A(_00041_));
 sg13g2_inv_1 _19624_ (.Y(_10662_),
    .A(_00045_));
 sg13g2_inv_1 _19625_ (.Y(_10663_),
    .A(_00047_));
 sg13g2_inv_1 _19626_ (.Y(_10664_),
    .A(_00052_));
 sg13g2_inv_1 _19627_ (.Y(_10665_),
    .A(_00055_));
 sg13g2_inv_1 _19628_ (.Y(_10666_),
    .A(net4725));
 sg13g2_inv_1 _19629_ (.Y(_10667_),
    .A(_00063_));
 sg13g2_inv_1 _19630_ (.Y(_10668_),
    .A(_00062_));
 sg13g2_inv_1 _19631_ (.Y(_10669_),
    .A(_00066_));
 sg13g2_inv_1 _19632_ (.Y(_10670_),
    .A(net4382));
 sg13g2_inv_1 _19633_ (.Y(_10671_),
    .A(_00071_));
 sg13g2_inv_1 _19634_ (.Y(_10672_),
    .A(_00074_));
 sg13g2_inv_1 _19635_ (.Y(_10673_),
    .A(_00076_));
 sg13g2_inv_1 _19636_ (.Y(_10674_),
    .A(net9179));
 sg13g2_inv_1 _19637_ (.Y(_10675_),
    .A(\soc_I.rx_uart_i.fifo_i.ram[13][0] ));
 sg13g2_inv_2 _19638_ (.Y(_10676_),
    .A(net9174));
 sg13g2_inv_1 _19639_ (.Y(_10677_),
    .A(\soc_I.rx_uart_i.fifo_i.ram[13][1] ));
 sg13g2_inv_1 _19640_ (.Y(_10678_),
    .A(\soc_I.rx_uart_i.fifo_i.ram[13][3] ));
 sg13g2_inv_1 _19641_ (.Y(_10679_),
    .A(\soc_I.rx_uart_i.fifo_i.ram[13][4] ));
 sg13g2_inv_1 _19642_ (.Y(_10680_),
    .A(\soc_I.rx_uart_i.fifo_i.ram[13][6] ));
 sg13g2_inv_1 _19643_ (.Y(_10681_),
    .A(\soc_I.rx_uart_i.fifo_i.ram[13][7] ));
 sg13g2_inv_1 _19644_ (.Y(_10682_),
    .A(_00081_));
 sg13g2_inv_1 _19645_ (.Y(_10683_),
    .A(_00085_));
 sg13g2_inv_1 _19646_ (.Y(_10684_),
    .A(_00103_));
 sg13g2_inv_1 _19647_ (.Y(_10685_),
    .A(_00121_));
 sg13g2_inv_1 _19648_ (.Y(_10686_),
    .A(_00120_));
 sg13g2_inv_1 _19649_ (.Y(_10687_),
    .A(_00126_));
 sg13g2_inv_1 _19650_ (.Y(_10688_),
    .A(_00131_));
 sg13g2_inv_1 _19651_ (.Y(_10689_),
    .A(_00130_));
 sg13g2_inv_1 _19652_ (.Y(_10690_),
    .A(_00141_));
 sg13g2_inv_1 _19653_ (.Y(_10691_),
    .A(_00140_));
 sg13g2_inv_1 _19654_ (.Y(_10692_),
    .A(_00145_));
 sg13g2_inv_1 _19655_ (.Y(_10693_),
    .A(_00148_));
 sg13g2_inv_1 _19656_ (.Y(_10694_),
    .A(_00151_));
 sg13g2_inv_1 _19657_ (.Y(_10695_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][0] ));
 sg13g2_inv_1 _19658_ (.Y(_10696_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][0] ));
 sg13g2_inv_1 _19659_ (.Y(_10697_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][0] ));
 sg13g2_inv_1 _19660_ (.Y(_10698_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][0] ));
 sg13g2_inv_1 _19661_ (.Y(_10699_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][1] ));
 sg13g2_inv_1 _19662_ (.Y(_10700_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][1] ));
 sg13g2_inv_1 _19663_ (.Y(_10701_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][1] ));
 sg13g2_inv_1 _19664_ (.Y(_10702_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][1] ));
 sg13g2_inv_1 _19665_ (.Y(_10703_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][2] ));
 sg13g2_inv_1 _19666_ (.Y(_10704_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][2] ));
 sg13g2_inv_1 _19667_ (.Y(_10705_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][2] ));
 sg13g2_inv_1 _19668_ (.Y(_10706_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][2] ));
 sg13g2_inv_1 _19669_ (.Y(_10707_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][3] ));
 sg13g2_inv_1 _19670_ (.Y(_10708_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][3] ));
 sg13g2_inv_1 _19671_ (.Y(_10709_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][3] ));
 sg13g2_inv_1 _19672_ (.Y(_10710_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][4] ));
 sg13g2_inv_1 _19673_ (.Y(_10711_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][4] ));
 sg13g2_inv_1 _19674_ (.Y(_10712_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][4] ));
 sg13g2_inv_1 _19675_ (.Y(_10713_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][5] ));
 sg13g2_inv_1 _19676_ (.Y(_10714_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][5] ));
 sg13g2_inv_1 _19677_ (.Y(_10715_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][6] ));
 sg13g2_inv_1 _19678_ (.Y(_10716_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][6] ));
 sg13g2_inv_1 _19679_ (.Y(_10717_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][6] ));
 sg13g2_inv_1 _19680_ (.Y(_10718_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][7] ));
 sg13g2_inv_1 _19681_ (.Y(_10719_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][7] ));
 sg13g2_inv_1 _19682_ (.Y(_10720_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][7] ));
 sg13g2_inv_1 _19683_ (.Y(_10721_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][7] ));
 sg13g2_inv_1 _19684_ (.Y(_10722_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][8] ));
 sg13g2_inv_1 _19685_ (.Y(_10723_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][8] ));
 sg13g2_inv_1 _19686_ (.Y(_10724_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][8] ));
 sg13g2_inv_1 _19687_ (.Y(_10725_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][8] ));
 sg13g2_inv_1 _19688_ (.Y(_10726_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][8] ));
 sg13g2_inv_1 _19689_ (.Y(_10727_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][8] ));
 sg13g2_inv_1 _19690_ (.Y(_10728_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][9] ));
 sg13g2_inv_1 _19691_ (.Y(_10729_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][9] ));
 sg13g2_inv_1 _19692_ (.Y(_10730_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][9] ));
 sg13g2_inv_1 _19693_ (.Y(_10731_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][9] ));
 sg13g2_inv_1 _19694_ (.Y(_10732_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][10] ));
 sg13g2_inv_1 _19695_ (.Y(_10733_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][10] ));
 sg13g2_inv_1 _19696_ (.Y(_10734_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][10] ));
 sg13g2_inv_1 _19697_ (.Y(_10735_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][10] ));
 sg13g2_inv_1 _19698_ (.Y(_10736_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][10] ));
 sg13g2_inv_1 _19699_ (.Y(_10737_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][11] ));
 sg13g2_inv_1 _19700_ (.Y(_10738_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][11] ));
 sg13g2_inv_1 _19701_ (.Y(_10739_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][11] ));
 sg13g2_inv_1 _19702_ (.Y(_10740_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][12] ));
 sg13g2_inv_1 _19703_ (.Y(_10741_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][12] ));
 sg13g2_inv_1 _19704_ (.Y(_10742_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][12] ));
 sg13g2_inv_1 _19705_ (.Y(_10743_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][12] ));
 sg13g2_inv_1 _19706_ (.Y(_10744_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][13] ));
 sg13g2_inv_1 _19707_ (.Y(_10745_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][13] ));
 sg13g2_inv_1 _19708_ (.Y(_10746_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][13] ));
 sg13g2_inv_1 _19709_ (.Y(_10747_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][13] ));
 sg13g2_inv_1 _19710_ (.Y(_10748_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][14] ));
 sg13g2_inv_1 _19711_ (.Y(_10749_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][14] ));
 sg13g2_inv_1 _19712_ (.Y(_10750_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][14] ));
 sg13g2_inv_1 _19713_ (.Y(_10751_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][14] ));
 sg13g2_inv_1 _19714_ (.Y(_10752_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][14] ));
 sg13g2_inv_1 _19715_ (.Y(_10753_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][15] ));
 sg13g2_inv_1 _19716_ (.Y(_10754_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][15] ));
 sg13g2_inv_1 _19717_ (.Y(_10755_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][15] ));
 sg13g2_inv_1 _19718_ (.Y(_10756_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][16] ));
 sg13g2_inv_1 _19719_ (.Y(_10757_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][16] ));
 sg13g2_inv_1 _19720_ (.Y(_10758_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][16] ));
 sg13g2_inv_1 _19721_ (.Y(_10759_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][16] ));
 sg13g2_inv_1 _19722_ (.Y(_10760_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][17] ));
 sg13g2_inv_1 _19723_ (.Y(_10761_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][17] ));
 sg13g2_inv_1 _19724_ (.Y(_10762_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][17] ));
 sg13g2_inv_1 _19725_ (.Y(_10763_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][17] ));
 sg13g2_inv_1 _19726_ (.Y(_10764_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][18] ));
 sg13g2_inv_1 _19727_ (.Y(_10765_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][18] ));
 sg13g2_inv_1 _19728_ (.Y(_10766_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][19] ));
 sg13g2_inv_1 _19729_ (.Y(_10767_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][19] ));
 sg13g2_inv_1 _19730_ (.Y(_10768_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][19] ));
 sg13g2_inv_1 _19731_ (.Y(_10769_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][19] ));
 sg13g2_inv_1 _19732_ (.Y(_10770_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][19] ));
 sg13g2_inv_1 _19733_ (.Y(_10771_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][20] ));
 sg13g2_inv_1 _19734_ (.Y(_10772_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][20] ));
 sg13g2_inv_1 _19735_ (.Y(_10773_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][20] ));
 sg13g2_inv_1 _19736_ (.Y(_10774_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][20] ));
 sg13g2_inv_1 _19737_ (.Y(_10775_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][21] ));
 sg13g2_inv_1 _19738_ (.Y(_10776_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][21] ));
 sg13g2_inv_1 _19739_ (.Y(_10777_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][21] ));
 sg13g2_inv_1 _19740_ (.Y(_10778_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][21] ));
 sg13g2_inv_1 _19741_ (.Y(_10779_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][22] ));
 sg13g2_inv_1 _19742_ (.Y(_10780_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][22] ));
 sg13g2_inv_1 _19743_ (.Y(_10781_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][22] ));
 sg13g2_inv_1 _19744_ (.Y(_10782_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][22] ));
 sg13g2_inv_1 _19745_ (.Y(_10783_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][22] ));
 sg13g2_inv_1 _19746_ (.Y(_10784_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][23] ));
 sg13g2_inv_1 _19747_ (.Y(_10785_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][23] ));
 sg13g2_inv_1 _19748_ (.Y(_10786_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][23] ));
 sg13g2_inv_1 _19749_ (.Y(_10787_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][23] ));
 sg13g2_inv_1 _19750_ (.Y(_10788_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][24] ));
 sg13g2_inv_1 _19751_ (.Y(_10789_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][24] ));
 sg13g2_inv_1 _19752_ (.Y(_10790_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][24] ));
 sg13g2_inv_1 _19753_ (.Y(_10791_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][25] ));
 sg13g2_inv_1 _19754_ (.Y(_10792_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][25] ));
 sg13g2_inv_1 _19755_ (.Y(_10793_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][25] ));
 sg13g2_inv_1 _19756_ (.Y(_10794_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][26] ));
 sg13g2_inv_1 _19757_ (.Y(_10795_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][26] ));
 sg13g2_inv_1 _19758_ (.Y(_10796_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][26] ));
 sg13g2_inv_1 _19759_ (.Y(_10797_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][26] ));
 sg13g2_inv_1 _19760_ (.Y(_10798_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][26] ));
 sg13g2_inv_1 _19761_ (.Y(_10799_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][27] ));
 sg13g2_inv_1 _19762_ (.Y(_10800_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][27] ));
 sg13g2_inv_1 _19763_ (.Y(_10801_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][27] ));
 sg13g2_inv_1 _19764_ (.Y(_10802_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][28] ));
 sg13g2_inv_1 _19765_ (.Y(_10803_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][28] ));
 sg13g2_inv_1 _19766_ (.Y(_10804_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][28] ));
 sg13g2_inv_1 _19767_ (.Y(_10805_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][28] ));
 sg13g2_inv_1 _19768_ (.Y(_10806_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][28] ));
 sg13g2_inv_1 _19769_ (.Y(_10807_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][29] ));
 sg13g2_inv_1 _19770_ (.Y(_10808_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][29] ));
 sg13g2_inv_1 _19771_ (.Y(_10809_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][29] ));
 sg13g2_inv_1 _19772_ (.Y(_10810_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][29] ));
 sg13g2_inv_1 _19773_ (.Y(_10811_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][30] ));
 sg13g2_inv_1 _19774_ (.Y(_10812_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][30] ));
 sg13g2_inv_1 _19775_ (.Y(_10813_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][30] ));
 sg13g2_inv_1 _19776_ (.Y(_10814_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][31] ));
 sg13g2_inv_1 _19777_ (.Y(_10815_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][31] ));
 sg13g2_inv_1 _19778_ (.Y(_10816_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][31] ));
 sg13g2_inv_1 _19779_ (.Y(_10817_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][31] ));
 sg13g2_inv_1 _19780_ (.Y(_10818_),
    .A(_00168_));
 sg13g2_inv_1 _19781_ (.Y(_10819_),
    .A(_00169_));
 sg13g2_inv_1 _19782_ (.Y(_10820_),
    .A(_00170_));
 sg13g2_inv_1 _19783_ (.Y(_10821_),
    .A(_00171_));
 sg13g2_inv_1 _19784_ (.Y(_10822_),
    .A(_00172_));
 sg13g2_inv_1 _19785_ (.Y(_10823_),
    .A(_00173_));
 sg13g2_inv_1 _19786_ (.Y(_10824_),
    .A(_00174_));
 sg13g2_inv_1 _19787_ (.Y(_10825_),
    .A(_00176_));
 sg13g2_inv_1 _19788_ (.Y(_10826_),
    .A(_00177_));
 sg13g2_inv_1 _19789_ (.Y(_10827_),
    .A(net5361));
 sg13g2_inv_1 _19790_ (.Y(_10828_),
    .A(_00180_));
 sg13g2_inv_1 _19791_ (.Y(_10829_),
    .A(_00181_));
 sg13g2_inv_1 _19792_ (.Y(_10830_),
    .A(_00182_));
 sg13g2_inv_1 _19793_ (.Y(_10831_),
    .A(_00183_));
 sg13g2_nor2b_2 _19794_ (.A(net9201),
    .B_N(net9200),
    .Y(_10832_));
 sg13g2_nor2b_1 _19795_ (.A(net9197),
    .B_N(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[0] ),
    .Y(_10833_));
 sg13g2_nand2_2 _19796_ (.Y(_10834_),
    .A(_10832_),
    .B(_10833_));
 sg13g2_nor2_1 _19797_ (.A(net9202),
    .B(net9204),
    .Y(_10835_));
 sg13g2_or2_2 _19798_ (.X(_10836_),
    .B(net9203),
    .A(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[4] ));
 sg13g2_nor2_2 _19799_ (.A(_10834_),
    .B(_10836_),
    .Y(_10837_));
 sg13g2_nor2b_2 _19800_ (.A(net9203),
    .B_N(net9202),
    .Y(_10838_));
 sg13g2_nand2b_2 _19801_ (.Y(_10839_),
    .B(net9202),
    .A_N(net9203));
 sg13g2_nor2_1 _19802_ (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[0] ),
    .B(net9197),
    .Y(_10840_));
 sg13g2_nand2_2 _19803_ (.Y(_10841_),
    .A(net9199),
    .B(net9201));
 sg13g2_nor3_2 _19804_ (.A(net9196),
    .B(net9197),
    .C(_10841_),
    .Y(_10842_));
 sg13g2_nand3_1 _19805_ (.B(net9201),
    .C(net8976),
    .A(net9199),
    .Y(_10843_));
 sg13g2_nor2_1 _19806_ (.A(_10839_),
    .B(_10843_),
    .Y(_10844_));
 sg13g2_nand2_2 _19807_ (.Y(_10845_),
    .A(net8978),
    .B(_10842_));
 sg13g2_nand2b_2 _19808_ (.Y(_10846_),
    .B(net8738),
    .A_N(_10837_));
 sg13g2_nand2_2 _19809_ (.Y(_10847_),
    .A(net9196),
    .B(net9197));
 sg13g2_nor2_1 _19810_ (.A(net9199),
    .B(net9201),
    .Y(_10848_));
 sg13g2_or2_2 _19811_ (.X(_10849_),
    .B(net9201),
    .A(net9200));
 sg13g2_nor3_2 _19812_ (.A(net9204),
    .B(_10847_),
    .C(_10849_),
    .Y(_10850_));
 sg13g2_nor2_2 _19813_ (.A(_10834_),
    .B(net8977),
    .Y(_10851_));
 sg13g2_inv_1 _19814_ (.Y(_10852_),
    .A(_10851_));
 sg13g2_nor2b_1 _19815_ (.A(net9199),
    .B_N(net9201),
    .Y(_10853_));
 sg13g2_and3_1 _19816_ (.X(_10854_),
    .A(net8978),
    .B(net8975),
    .C(net8973));
 sg13g2_nand3_1 _19817_ (.B(net8975),
    .C(net8973),
    .A(net8978),
    .Y(_10855_));
 sg13g2_nor2_2 _19818_ (.A(_10846_),
    .B(_10851_),
    .Y(_10856_));
 sg13g2_o21ai_1 _19819_ (.B1(net8738),
    .Y(_10857_),
    .A1(net9204),
    .A2(_10834_));
 sg13g2_nor3_2 _19820_ (.A(_10850_),
    .B(net8859),
    .C(net8667),
    .Y(_10858_));
 sg13g2_or3_2 _19821_ (.A(_10850_),
    .B(net8859),
    .C(net8667),
    .X(_10859_));
 sg13g2_nor2b_2 _19822_ (.A(net9196),
    .B_N(net9198),
    .Y(_10860_));
 sg13g2_nand2b_2 _19823_ (.Y(_10861_),
    .B(net9197),
    .A_N(net9196));
 sg13g2_and2_1 _19824_ (.A(net8973),
    .B(_10860_),
    .X(_10862_));
 sg13g2_nand2_2 _19825_ (.Y(_10863_),
    .A(_10853_),
    .B(_10860_));
 sg13g2_nor2_1 _19826_ (.A(_10839_),
    .B(_10863_),
    .Y(_10864_));
 sg13g2_nand2_2 _19827_ (.Y(_10865_),
    .A(net8978),
    .B(_10862_));
 sg13g2_nand2_2 _19828_ (.Y(_10866_),
    .A(net8976),
    .B(_10848_));
 sg13g2_nor2_2 _19829_ (.A(_10836_),
    .B(_10866_),
    .Y(_10867_));
 sg13g2_nor2_1 _19830_ (.A(net8724),
    .B(_10867_),
    .Y(_10868_));
 sg13g2_or2_2 _19831_ (.X(_10869_),
    .B(_10867_),
    .A(net8724));
 sg13g2_nand3_1 _19832_ (.B(net8975),
    .C(net8973),
    .A(net8979),
    .Y(_10870_));
 sg13g2_nand2_1 _19833_ (.Y(_10871_),
    .A(net8979),
    .B(_10860_));
 sg13g2_nand3_1 _19834_ (.B(net8979),
    .C(_10860_),
    .A(_10832_),
    .Y(_10872_));
 sg13g2_nand2_2 _19835_ (.Y(_10873_),
    .A(_10870_),
    .B(_10872_));
 sg13g2_nand2b_2 _19836_ (.Y(_10874_),
    .B(net9703),
    .A_N(net9698));
 sg13g2_nand2b_1 _19837_ (.Y(_10875_),
    .B(_10873_),
    .A_N(_10874_));
 sg13g2_nor2_2 _19838_ (.A(_10836_),
    .B(_10863_),
    .Y(_10876_));
 sg13g2_nand2_1 _19839_ (.Y(_10877_),
    .A(_10835_),
    .B(_10862_));
 sg13g2_nand2_2 _19840_ (.Y(_10878_),
    .A(net9698),
    .B(net9702));
 sg13g2_nand2_1 _19841_ (.Y(_10879_),
    .A(_10876_),
    .B(_10878_));
 sg13g2_nor2_2 _19842_ (.A(_10836_),
    .B(_10843_),
    .Y(_10880_));
 sg13g2_nand4_1 _19843_ (.B(net9201),
    .C(net8979),
    .A(net9199),
    .Y(_10881_),
    .D(net8976));
 sg13g2_a221oi_1 _19844_ (.B2(_10878_),
    .C1(net9196),
    .B1(_10876_),
    .A1(_10835_),
    .Y(_10882_),
    .A2(_10842_));
 sg13g2_nand2_1 _19845_ (.Y(_10883_),
    .A(net9201),
    .B(net8980));
 sg13g2_nand3_1 _19846_ (.B(net8980),
    .C(net8979),
    .A(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[3] ),
    .Y(_10884_));
 sg13g2_nand4_1 _19847_ (.B(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[3] ),
    .C(net8980),
    .A(net9199),
    .Y(_10885_),
    .D(_10835_));
 sg13g2_o21ai_1 _19848_ (.B1(_10885_),
    .Y(_10886_),
    .A1(net9204),
    .A2(_10863_));
 sg13g2_nor2_1 _19849_ (.A(_10873_),
    .B(_10880_),
    .Y(_10887_));
 sg13g2_nor3_1 _19850_ (.A(_10873_),
    .B(_10880_),
    .C(_10886_),
    .Y(_10888_));
 sg13g2_a21oi_2 _19851_ (.B1(_10888_),
    .Y(_10889_),
    .A2(_10882_),
    .A1(_10875_));
 sg13g2_a21o_2 _19852_ (.A2(_10882_),
    .A1(_10875_),
    .B1(_10888_),
    .X(_10890_));
 sg13g2_nor2_2 _19853_ (.A(net9430),
    .B(net9431),
    .Y(_10891_));
 sg13g2_nand4_1 _19854_ (.B(net9428),
    .C(_00189_),
    .A(net9425),
    .Y(_10892_),
    .D(_10891_));
 sg13g2_nor2b_1 _19855_ (.A(net9425),
    .B_N(net9428),
    .Y(_10893_));
 sg13g2_nand3_1 _19856_ (.B(_10891_),
    .C(_10893_),
    .A(_00189_),
    .Y(_10894_));
 sg13g2_nor2_2 _19857_ (.A(net9425),
    .B(net9428),
    .Y(_10895_));
 sg13g2_nand3_1 _19858_ (.B(_10891_),
    .C(_10895_),
    .A(net9424),
    .Y(_10896_));
 sg13g2_nor2b_1 _19859_ (.A(net9428),
    .B_N(net9425),
    .Y(_10897_));
 sg13g2_nor2_1 _19860_ (.A(net9427),
    .B(net9430),
    .Y(_10898_));
 sg13g2_and2_1 _19861_ (.A(_10891_),
    .B(_10897_),
    .X(_10899_));
 sg13g2_nand3b_1 _19862_ (.B(_10891_),
    .C(_10897_),
    .Y(_10900_),
    .A_N(net9423));
 sg13g2_and4_2 _19863_ (.A(_10892_),
    .B(_10894_),
    .C(_10896_),
    .D(_10900_),
    .X(_10901_));
 sg13g2_nor2_1 _19864_ (.A(net9423),
    .B(\soc_I.kianv_I.Instr[27] ),
    .Y(_10902_));
 sg13g2_nand3_1 _19865_ (.B(_10895_),
    .C(_10902_),
    .A(net9430),
    .Y(_10903_));
 sg13g2_and2_1 _19866_ (.A(net9431),
    .B(_00189_),
    .X(_10904_));
 sg13g2_nand3_1 _19867_ (.B(_10895_),
    .C(_10904_),
    .A(net9430),
    .Y(_10905_));
 sg13g2_nor3_2 _19868_ (.A(net9425),
    .B(net9427),
    .C(net9430),
    .Y(_10906_));
 sg13g2_nand2_1 _19869_ (.Y(_10907_),
    .A(_00189_),
    .B(_10906_));
 sg13g2_and3_1 _19870_ (.X(_10908_),
    .A(_10903_),
    .B(_10905_),
    .C(_10907_));
 sg13g2_and2_1 _19871_ (.A(_10901_),
    .B(_10908_),
    .X(_10909_));
 sg13g2_nand3_1 _19872_ (.B(_10891_),
    .C(_10893_),
    .A(net9423),
    .Y(_10910_));
 sg13g2_nand3_1 _19873_ (.B(_10908_),
    .C(_10910_),
    .A(_10901_),
    .Y(_10911_));
 sg13g2_a21oi_2 _19874_ (.B1(_10865_),
    .Y(_10912_),
    .A2(_10911_),
    .A1(_10892_));
 sg13g2_nor2b_1 _19875_ (.A(net9703),
    .B_N(net9698),
    .Y(_10913_));
 sg13g2_nand2_1 _19876_ (.Y(_10914_),
    .A(net9706),
    .B(net8972));
 sg13g2_nor2b_2 _19877_ (.A(net9701),
    .B_N(net9707),
    .Y(_10915_));
 sg13g2_nand2b_2 _19878_ (.Y(_10916_),
    .B(net9707),
    .A_N(net9701));
 sg13g2_nand2_1 _19879_ (.Y(_10917_),
    .A(_00188_),
    .B(net8962));
 sg13g2_nand2_1 _19880_ (.Y(_10918_),
    .A(_10914_),
    .B(_10917_));
 sg13g2_nand2_2 _19881_ (.Y(_10919_),
    .A(net9702),
    .B(net9706));
 sg13g2_nand2b_1 _19882_ (.Y(_10920_),
    .B(_10587_),
    .A_N(_10919_));
 sg13g2_nand3_1 _19883_ (.B(_10917_),
    .C(_10920_),
    .A(_10914_),
    .Y(_10921_));
 sg13g2_nor2_1 _19884_ (.A(net9702),
    .B(_00212_),
    .Y(_10922_));
 sg13g2_or2_1 _19885_ (.X(_10923_),
    .B(_00212_),
    .A(net9702));
 sg13g2_nor2_2 _19886_ (.A(net9699),
    .B(net9703),
    .Y(_10924_));
 sg13g2_or2_2 _19887_ (.X(_10925_),
    .B(net9704),
    .A(net9698));
 sg13g2_o21ai_1 _19888_ (.B1(_10923_),
    .Y(_10926_),
    .A1(_10915_),
    .A2(_10924_));
 sg13g2_nand3_1 _19889_ (.B(_10921_),
    .C(_10926_),
    .A(_10873_),
    .Y(_10927_));
 sg13g2_nand2_2 _19890_ (.Y(_10928_),
    .A(_10879_),
    .B(_10927_));
 sg13g2_or2_1 _19891_ (.X(_10929_),
    .B(_10928_),
    .A(_10912_));
 sg13g2_o21ai_1 _19892_ (.B1(_10889_),
    .Y(_10930_),
    .A1(_10912_),
    .A2(_10928_));
 sg13g2_nor2_1 _19893_ (.A(net9431),
    .B(_10907_),
    .Y(_10931_));
 sg13g2_nor2_1 _19894_ (.A(_10901_),
    .B(_10931_),
    .Y(_10932_));
 sg13g2_and2_1 _19895_ (.A(_00189_),
    .B(_10899_),
    .X(_10933_));
 sg13g2_nand2_1 _19896_ (.Y(_10934_),
    .A(_00189_),
    .B(_10899_));
 sg13g2_nand3_1 _19897_ (.B(_10891_),
    .C(_10897_),
    .A(net9423),
    .Y(_10935_));
 sg13g2_and4_1 _19898_ (.A(_10892_),
    .B(_10907_),
    .C(_10910_),
    .D(_10935_),
    .X(_10936_));
 sg13g2_nor2_1 _19899_ (.A(_10458_),
    .B(_10907_),
    .Y(_10937_));
 sg13g2_a21oi_1 _19900_ (.A1(_10904_),
    .A2(_10906_),
    .Y(_10938_),
    .B1(net9425));
 sg13g2_or3_1 _19901_ (.A(_10933_),
    .B(_10936_),
    .C(_10938_),
    .X(_10939_));
 sg13g2_nand3_1 _19902_ (.B(_10932_),
    .C(_10939_),
    .A(net8727),
    .Y(_10940_));
 sg13g2_nand2b_1 _19903_ (.Y(_10941_),
    .B(_10919_),
    .A_N(net9699));
 sg13g2_nand3_1 _19904_ (.B(net9708),
    .C(_10923_),
    .A(net9698),
    .Y(_10942_));
 sg13g2_nand3_1 _19905_ (.B(_10941_),
    .C(_10942_),
    .A(_10873_),
    .Y(_10943_));
 sg13g2_or2_1 _19906_ (.X(_10944_),
    .B(_10910_),
    .A(_10865_));
 sg13g2_a21oi_1 _19907_ (.A1(_10876_),
    .A2(net8972),
    .Y(_10945_),
    .B1(_10880_));
 sg13g2_and3_1 _19908_ (.X(_10946_),
    .A(_10943_),
    .B(_10944_),
    .C(_10945_));
 sg13g2_and2_2 _19909_ (.A(_10940_),
    .B(_10946_),
    .X(_10947_));
 sg13g2_inv_2 _19910_ (.Y(_10948_),
    .A(_10947_));
 sg13g2_a21oi_1 _19911_ (.A1(_10901_),
    .A2(_10908_),
    .Y(_10949_),
    .B1(net9425));
 sg13g2_nand3b_1 _19912_ (.B(net8727),
    .C(_10939_),
    .Y(_10950_),
    .A_N(_10949_));
 sg13g2_nand3_1 _19913_ (.B(_10876_),
    .C(_10921_),
    .A(_10874_),
    .Y(_10951_));
 sg13g2_a21oi_2 _19914_ (.B1(net9706),
    .Y(_10952_),
    .A2(net9702),
    .A1(net9699));
 sg13g2_a21oi_1 _19915_ (.A1(net9706),
    .A2(_10587_),
    .Y(_10953_),
    .B1(_10952_));
 sg13g2_nand3b_1 _19916_ (.B(\soc_I.kianv_I.Instr[1] ),
    .C(\soc_I.kianv_I.Instr[0] ),
    .Y(_10954_),
    .A_N(\soc_I.kianv_I.Instr[3] ));
 sg13g2_nor2_1 _19917_ (.A(_10470_),
    .B(_10954_),
    .Y(_10955_));
 sg13g2_nand3b_1 _19918_ (.B(\soc_I.kianv_I.Instr[4] ),
    .C(_00214_),
    .Y(_10956_),
    .A_N(net9713));
 sg13g2_nor3_2 _19919_ (.A(_10470_),
    .B(_10954_),
    .C(_10956_),
    .Y(_10957_));
 sg13g2_nand3b_1 _19920_ (.B(net8972),
    .C(net9706),
    .Y(_10958_),
    .A_N(_00213_));
 sg13g2_a21oi_1 _19921_ (.A1(_10926_),
    .A2(_10958_),
    .Y(_10959_),
    .B1(_10957_));
 sg13g2_a221oi_1 _19922_ (.B2(_10925_),
    .C1(_10922_),
    .B1(_10916_),
    .A1(net9426),
    .Y(_10960_),
    .A2(net9713));
 sg13g2_a21oi_1 _19923_ (.A1(_10870_),
    .A2(_10872_),
    .Y(_10961_),
    .B1(_10960_));
 sg13g2_o21ai_1 _19924_ (.B1(_10961_),
    .Y(_10962_),
    .A1(_10953_),
    .A2(_10959_));
 sg13g2_and3_2 _19925_ (.X(_10963_),
    .A(_10885_),
    .B(_10951_),
    .C(_10962_));
 sg13g2_and2_2 _19926_ (.A(_10950_),
    .B(_10963_),
    .X(_10964_));
 sg13g2_nand2_2 _19927_ (.Y(_10965_),
    .A(_10950_),
    .B(_10963_));
 sg13g2_nand2_2 _19928_ (.Y(_10966_),
    .A(_10947_),
    .B(net8529));
 sg13g2_nor2_1 _19929_ (.A(_10930_),
    .B(_10966_),
    .Y(_10967_));
 sg13g2_nand4_1 _19930_ (.B(net9197),
    .C(net8979),
    .A(net9196),
    .Y(_10968_),
    .D(net8973));
 sg13g2_nor2_1 _19931_ (.A(net8977),
    .B(_10866_),
    .Y(_10969_));
 sg13g2_nand3_1 _19932_ (.B(net8975),
    .C(net8974),
    .A(net8978),
    .Y(_10970_));
 sg13g2_nand3_1 _19933_ (.B(net8974),
    .C(_10860_),
    .A(net8979),
    .Y(_10971_));
 sg13g2_nand4_1 _19934_ (.B(_10968_),
    .C(_10970_),
    .A(_10870_),
    .Y(_10972_),
    .D(_10971_));
 sg13g2_nor3_1 _19935_ (.A(net8977),
    .B(_10849_),
    .C(_10861_),
    .Y(_10973_));
 sg13g2_nand3_1 _19936_ (.B(net8974),
    .C(_10860_),
    .A(_10838_),
    .Y(_10974_));
 sg13g2_nand4_1 _19937_ (.B(net9197),
    .C(net8978),
    .A(net9196),
    .Y(_10975_),
    .D(net8973));
 sg13g2_nand2_2 _19938_ (.Y(_10976_),
    .A(net8842),
    .B(_10975_));
 sg13g2_nor2_1 _19939_ (.A(_10972_),
    .B(_10976_),
    .Y(_10977_));
 sg13g2_o21ai_1 _19940_ (.B1(_10977_),
    .Y(_10978_),
    .A1(net8974),
    .A2(_10871_));
 sg13g2_nand2_1 _19941_ (.Y(_10979_),
    .A(net8980),
    .B(_10848_));
 sg13g2_nor2_1 _19942_ (.A(_10836_),
    .B(_10979_),
    .Y(_10980_));
 sg13g2_nand3_1 _19943_ (.B(net8979),
    .C(net8974),
    .A(net8980),
    .Y(_10981_));
 sg13g2_and2_1 _19944_ (.A(_10884_),
    .B(_10981_),
    .X(_10982_));
 sg13g2_nand2_1 _19945_ (.Y(_10983_),
    .A(_10884_),
    .B(_10981_));
 sg13g2_nor3_2 _19946_ (.A(net9199),
    .B(_10839_),
    .C(_10883_),
    .Y(_10984_));
 sg13g2_nand3_1 _19947_ (.B(net8978),
    .C(net8973),
    .A(net8980),
    .Y(_10985_));
 sg13g2_o21ai_1 _19948_ (.B1(_10985_),
    .Y(_10986_),
    .A1(_10865_),
    .A2(_10937_));
 sg13g2_a22oi_1 _19949_ (.Y(_10987_),
    .B1(net8650),
    .B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[31] ),
    .A2(net8564),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[31] ));
 sg13g2_nor2_1 _19950_ (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[31] ),
    .B(net8717),
    .Y(_10988_));
 sg13g2_nor4_2 _19951_ (.A(net8728),
    .B(net8569),
    .C(net8715),
    .Y(_10989_),
    .D(_10984_));
 sg13g2_a21oi_1 _19952_ (.A1(net8717),
    .A2(_10987_),
    .Y(_10990_),
    .B1(_10988_));
 sg13g2_nand2_1 _19953_ (.Y(_10991_),
    .A(\soc_I.PC[31] ),
    .B(net8525));
 sg13g2_nor2b_2 _19954_ (.A(_10990_),
    .B_N(_10991_),
    .Y(_10992_));
 sg13g2_nand2b_2 _19955_ (.Y(_10993_),
    .B(_10991_),
    .A_N(_10990_));
 sg13g2_nand4_1 _19956_ (.B(_10885_),
    .C(_10981_),
    .A(_10881_),
    .Y(_10994_),
    .D(_10985_));
 sg13g2_nor3_2 _19957_ (.A(_10972_),
    .B(_10976_),
    .C(_10994_),
    .Y(_10995_));
 sg13g2_or3_1 _19958_ (.A(_10972_),
    .B(_10976_),
    .C(_10994_),
    .X(_10996_));
 sg13g2_nor2_2 _19959_ (.A(\soc_I.kianv_I.Instr[2] ),
    .B(_10954_),
    .Y(_10997_));
 sg13g2_nand2_1 _19960_ (.Y(_10998_),
    .A(net9713),
    .B(net9715));
 sg13g2_nor3_1 _19961_ (.A(\soc_I.kianv_I.Instr[2] ),
    .B(_10954_),
    .C(_10998_),
    .Y(_10999_));
 sg13g2_nand3_1 _19962_ (.B(net9715),
    .C(_10997_),
    .A(net9713),
    .Y(_11000_));
 sg13g2_nand2_1 _19963_ (.Y(_11001_),
    .A(net9702),
    .B(_00188_));
 sg13g2_o21ai_1 _19964_ (.B1(net9704),
    .Y(_11002_),
    .A1(net9699),
    .A2(_00188_));
 sg13g2_a21oi_1 _19965_ (.A1(_10952_),
    .A2(_11001_),
    .Y(_11003_),
    .B1(_00214_));
 sg13g2_and2_1 _19966_ (.A(_10999_),
    .B(_11003_),
    .X(_11004_));
 sg13g2_nand2b_1 _19967_ (.Y(_11005_),
    .B(net9713),
    .A_N(net9715));
 sg13g2_nor2_2 _19968_ (.A(_00214_),
    .B(_11005_),
    .Y(_11006_));
 sg13g2_nor3_1 _19969_ (.A(\soc_I.kianv_I.Instr[2] ),
    .B(_10954_),
    .C(_10956_),
    .Y(_11007_));
 sg13g2_a221oi_1 _19970_ (.B2(_10955_),
    .C1(_11007_),
    .B1(_11006_),
    .A1(_10999_),
    .Y(_11008_),
    .A2(_11003_));
 sg13g2_nor2_1 _19971_ (.A(net9712),
    .B(net9715),
    .Y(_11009_));
 sg13g2_nor4_2 _19972_ (.A(net9712),
    .B(net9715),
    .C(\soc_I.kianv_I.Instr[2] ),
    .Y(_11010_),
    .D(_10954_));
 sg13g2_nand2_2 _19973_ (.Y(_11011_),
    .A(_10997_),
    .B(_11009_));
 sg13g2_nand2b_2 _19974_ (.Y(_11012_),
    .B(_11010_),
    .A_N(net9713));
 sg13g2_nand2_1 _19975_ (.Y(_11013_),
    .A(_11008_),
    .B(_11012_));
 sg13g2_a21o_1 _19976_ (.A2(_11012_),
    .A1(_11008_),
    .B1(_00189_),
    .X(_11014_));
 sg13g2_nand3_1 _19977_ (.B(_11008_),
    .C(_11012_),
    .A(net9424),
    .Y(_11015_));
 sg13g2_nand3_1 _19978_ (.B(_11014_),
    .C(_11015_),
    .A(net8643),
    .Y(_11016_));
 sg13g2_nor2_1 _19979_ (.A(net9199),
    .B(_10884_),
    .Y(_11017_));
 sg13g2_nor4_1 _19980_ (.A(_10867_),
    .B(_10976_),
    .C(_10984_),
    .D(_11017_),
    .Y(_11018_));
 sg13g2_or4_1 _19981_ (.A(_10867_),
    .B(_10976_),
    .C(_10984_),
    .D(_11017_),
    .X(_11019_));
 sg13g2_a21oi_2 _19982_ (.B1(net8636),
    .Y(_11020_),
    .A2(net8644),
    .A1(_00217_));
 sg13g2_and2_2 _19983_ (.A(_11016_),
    .B(_11020_),
    .X(_11021_));
 sg13g2_nand2_2 _19984_ (.Y(_11022_),
    .A(_11016_),
    .B(_11020_));
 sg13g2_and4_1 _19985_ (.A(_10940_),
    .B(_10946_),
    .C(_10950_),
    .D(_10963_),
    .X(_11023_));
 sg13g2_nand2_2 _19986_ (.Y(_11024_),
    .A(_10947_),
    .B(_10964_));
 sg13g2_nor4_1 _19987_ (.A(net9426),
    .B(net9427),
    .C(_10901_),
    .D(_10931_),
    .Y(_11025_));
 sg13g2_o21ai_1 _19988_ (.B1(net8727),
    .Y(_11026_),
    .A1(_10909_),
    .A2(_11025_));
 sg13g2_or2_2 _19989_ (.X(_11027_),
    .B(_10878_),
    .A(_10877_));
 sg13g2_nand2_2 _19990_ (.Y(_11028_),
    .A(_11026_),
    .B(_11027_));
 sg13g2_nor3_2 _19991_ (.A(_10889_),
    .B(_10912_),
    .C(_10928_),
    .Y(_11029_));
 sg13g2_nand2b_1 _19992_ (.Y(_11030_),
    .B(_10890_),
    .A_N(_10929_));
 sg13g2_nand2_2 _19993_ (.Y(_11031_),
    .A(_11028_),
    .B(_11029_));
 sg13g2_nor2_1 _19994_ (.A(_11024_),
    .B(_11031_),
    .Y(_11032_));
 sg13g2_nand3_1 _19995_ (.B(_11028_),
    .C(_11029_),
    .A(_11023_),
    .Y(_11033_));
 sg13g2_a22oi_1 _19996_ (.Y(_11034_),
    .B1(_10950_),
    .B2(_10963_),
    .A2(_10946_),
    .A1(_10940_));
 sg13g2_nand2_1 _19997_ (.Y(_11035_),
    .A(_10948_),
    .B(net8529));
 sg13g2_nor3_2 _19998_ (.A(_10890_),
    .B(_10912_),
    .C(_10928_),
    .Y(_11036_));
 sg13g2_and2_1 _19999_ (.A(_11023_),
    .B(_11036_),
    .X(_11037_));
 sg13g2_o21ai_1 _20000_ (.B1(_11036_),
    .Y(_11038_),
    .A1(_11023_),
    .A2(_11034_));
 sg13g2_nand3_1 _20001_ (.B(net8529),
    .C(_11029_),
    .A(_10947_),
    .Y(_11039_));
 sg13g2_and2_1 _20002_ (.A(_10930_),
    .B(_11026_),
    .X(_11040_));
 sg13g2_nor2_1 _20003_ (.A(_10890_),
    .B(net8529),
    .Y(_11041_));
 sg13g2_and4_2 _20004_ (.A(_11033_),
    .B(_11038_),
    .C(_11039_),
    .D(_11040_),
    .X(_11042_));
 sg13g2_nand4_1 _20005_ (.B(_11038_),
    .C(_11039_),
    .A(_11033_),
    .Y(_11043_),
    .D(_11040_));
 sg13g2_xnor2_1 _20006_ (.Y(_11044_),
    .A(_11022_),
    .B(net8313));
 sg13g2_nand2_1 _20007_ (.Y(_11045_),
    .A(net8314),
    .B(_11044_));
 sg13g2_nor2_1 _20008_ (.A(net8314),
    .B(_11044_),
    .Y(_11046_));
 sg13g2_xnor2_1 _20009_ (.Y(_11047_),
    .A(net8314),
    .B(_11044_));
 sg13g2_a22oi_1 _20010_ (.Y(_11048_),
    .B1(net8651),
    .B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[30] ),
    .A2(net8565),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[30] ));
 sg13g2_nor2_1 _20011_ (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[30] ),
    .B(net8719),
    .Y(_11049_));
 sg13g2_a21oi_1 _20012_ (.A1(net8719),
    .A2(_11048_),
    .Y(_11050_),
    .B1(_11049_));
 sg13g2_nand2_1 _20013_ (.Y(_11051_),
    .A(\soc_I.PC[30] ),
    .B(net8525));
 sg13g2_nor2b_2 _20014_ (.A(_11050_),
    .B_N(_11051_),
    .Y(_11052_));
 sg13g2_nand2b_2 _20015_ (.Y(_11053_),
    .B(_11051_),
    .A_N(_11050_));
 sg13g2_nand2_1 _20016_ (.Y(_11054_),
    .A(net9714),
    .B(_11009_));
 sg13g2_and2_2 _20017_ (.A(net9713),
    .B(_11010_),
    .X(_11055_));
 sg13g2_and2_1 _20018_ (.A(_10997_),
    .B(_11006_),
    .X(_11056_));
 sg13g2_nand2_1 _20019_ (.Y(_11057_),
    .A(_10997_),
    .B(_11006_));
 sg13g2_and3_1 _20020_ (.X(_11058_),
    .A(_11008_),
    .B(_11011_),
    .C(_11056_));
 sg13g2_or2_1 _20021_ (.X(_11059_),
    .B(_11058_),
    .A(_11055_));
 sg13g2_a221oi_1 _20022_ (.B2(net9423),
    .C1(net8649),
    .B1(_11059_),
    .A1(_10588_),
    .Y(_11060_),
    .A2(_11013_));
 sg13g2_inv_1 _20023_ (.Y(_11061_),
    .A(net8523));
 sg13g2_nor4_2 _20024_ (.A(net9712),
    .B(_10470_),
    .C(_10954_),
    .Y(_11062_),
    .D(_10998_));
 sg13g2_nor2_2 _20025_ (.A(_10957_),
    .B(_11062_),
    .Y(_11063_));
 sg13g2_or2_1 _20026_ (.X(_11064_),
    .B(_11062_),
    .A(_10957_));
 sg13g2_nand2_1 _20027_ (.Y(_11065_),
    .A(_11057_),
    .B(net8711));
 sg13g2_and4_2 _20028_ (.A(_11008_),
    .B(_11011_),
    .C(_11057_),
    .D(net8711),
    .X(_11066_));
 sg13g2_nand4_1 _20029_ (.B(_11011_),
    .C(_11057_),
    .A(_11008_),
    .Y(_11067_),
    .D(net8711));
 sg13g2_a21oi_2 _20030_ (.B1(_11061_),
    .Y(_11068_),
    .A2(_11066_),
    .A1(net9423));
 sg13g2_nand2_1 _20031_ (.Y(_11069_),
    .A(net9426),
    .B(net8709));
 sg13g2_a221oi_1 _20032_ (.B2(_11069_),
    .C1(net8637),
    .B1(net8309),
    .A1(_00218_),
    .Y(_11070_),
    .A2(net8649));
 sg13g2_xnor2_1 _20033_ (.Y(_11071_),
    .A(net8311),
    .B(net8008));
 sg13g2_nor2_1 _20034_ (.A(_11052_),
    .B(_11071_),
    .Y(_11072_));
 sg13g2_xnor2_1 _20035_ (.Y(_11073_),
    .A(_11052_),
    .B(_11071_));
 sg13g2_inv_1 _20036_ (.Y(_11074_),
    .A(_11073_));
 sg13g2_a22oi_1 _20037_ (.Y(_11075_),
    .B1(net8654),
    .B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[29] ),
    .A2(net8568),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[29] ));
 sg13g2_nor2_1 _20038_ (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[29] ),
    .B(net8718),
    .Y(_11076_));
 sg13g2_a21oi_1 _20039_ (.A1(net8718),
    .A2(_11075_),
    .Y(_11077_),
    .B1(_11076_));
 sg13g2_a21oi_1 _20040_ (.A1(\soc_I.PC[29] ),
    .A2(net8524),
    .Y(_11078_),
    .B1(_11077_));
 sg13g2_nand2_1 _20041_ (.Y(_11079_),
    .A(net9429),
    .B(net8710));
 sg13g2_a221oi_1 _20042_ (.B2(_11079_),
    .C1(net8635),
    .B1(net8309),
    .A1(_00219_),
    .Y(_11080_),
    .A2(net8644));
 sg13g2_xnor2_1 _20043_ (.Y(_11081_),
    .A(net8311),
    .B(net8007));
 sg13g2_and2_1 _20044_ (.A(net8307),
    .B(_11081_),
    .X(_11082_));
 sg13g2_a221oi_1 _20045_ (.B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[7] ),
    .C1(net8712),
    .B1(net8650),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[7] ),
    .Y(_11083_),
    .A2(net8564));
 sg13g2_nor2_1 _20046_ (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[7] ),
    .B(net8719),
    .Y(_11084_));
 sg13g2_nand2_1 _20047_ (.Y(_11085_),
    .A(\soc_I.PC[7] ),
    .B(net8524));
 sg13g2_o21ai_1 _20048_ (.B1(_11085_),
    .Y(_11086_),
    .A1(_11083_),
    .A2(_11084_));
 sg13g2_inv_2 _20049_ (.Y(_11087_),
    .A(_11086_));
 sg13g2_nand2_2 _20050_ (.Y(_11088_),
    .A(net9431),
    .B(net8711));
 sg13g2_a21o_1 _20051_ (.A2(net8649),
    .A1(_00235_),
    .B1(net8637),
    .X(_11089_));
 sg13g2_a21oi_2 _20052_ (.B1(_11089_),
    .Y(_11090_),
    .A2(_11088_),
    .A1(net8643));
 sg13g2_xnor2_1 _20053_ (.Y(_11091_),
    .A(net8312),
    .B(net8522));
 sg13g2_nor2_1 _20054_ (.A(_11087_),
    .B(_11091_),
    .Y(_11092_));
 sg13g2_a221oi_1 _20055_ (.B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[6] ),
    .C1(net8713),
    .B1(net8652),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[6] ),
    .Y(_11093_),
    .A2(net8566));
 sg13g2_nor2_1 _20056_ (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[6] ),
    .B(net8720),
    .Y(_11094_));
 sg13g2_nand2_1 _20057_ (.Y(_11095_),
    .A(\soc_I.PC[6] ),
    .B(net8526));
 sg13g2_o21ai_1 _20058_ (.B1(_11095_),
    .Y(_11096_),
    .A1(_11093_),
    .A2(_11094_));
 sg13g2_inv_2 _20059_ (.Y(_11097_),
    .A(_11096_));
 sg13g2_nand2_2 _20060_ (.Y(_11098_),
    .A(\soc_I.kianv_I.Instr[26] ),
    .B(net8711));
 sg13g2_a21o_1 _20061_ (.A2(net8647),
    .A1(_00187_),
    .B1(net8637),
    .X(_11099_));
 sg13g2_a21oi_2 _20062_ (.B1(_11099_),
    .Y(_11100_),
    .A2(_11098_),
    .A1(net8642));
 sg13g2_xnor2_1 _20063_ (.Y(_11101_),
    .A(net8310),
    .B(net8521));
 sg13g2_or2_1 _20064_ (.X(_11102_),
    .B(_11101_),
    .A(_11097_));
 sg13g2_a221oi_1 _20065_ (.B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[5] ),
    .C1(net8713),
    .B1(net8652),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[5] ),
    .Y(_11103_),
    .A2(net8566));
 sg13g2_nor2_1 _20066_ (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[5] ),
    .B(net8721),
    .Y(_11104_));
 sg13g2_nand2_1 _20067_ (.Y(_11105_),
    .A(\soc_I.PC[5] ),
    .B(net8526));
 sg13g2_o21ai_1 _20068_ (.B1(_11105_),
    .Y(_11106_),
    .A1(_11103_),
    .A2(_11104_));
 sg13g2_a21oi_1 _20069_ (.A1(\soc_I.kianv_I.Instr[25] ),
    .A2(_11063_),
    .Y(_11107_),
    .B1(net8646));
 sg13g2_a21oi_1 _20070_ (.A1(_00193_),
    .A2(net8647),
    .Y(_11108_),
    .B1(net8636));
 sg13g2_nor2b_1 _20071_ (.A(_11107_),
    .B_N(_11108_),
    .Y(_11109_));
 sg13g2_xnor2_1 _20072_ (.Y(_11110_),
    .A(net8313),
    .B(net8520));
 sg13g2_nand2_1 _20073_ (.Y(_11111_),
    .A(net8304),
    .B(_11110_));
 sg13g2_inv_1 _20074_ (.Y(_11112_),
    .A(_11111_));
 sg13g2_nor2_1 _20075_ (.A(net8304),
    .B(_11110_),
    .Y(_11113_));
 sg13g2_a221oi_1 _20076_ (.B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[4] ),
    .C1(net8713),
    .B1(net8652),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[4] ),
    .Y(_11114_),
    .A2(net8566));
 sg13g2_a21oi_1 _20077_ (.A1(_10492_),
    .A2(net8713),
    .Y(_11115_),
    .B1(_11114_));
 sg13g2_nand2_1 _20078_ (.Y(_11116_),
    .A(\soc_I.PC[4] ),
    .B(net8526));
 sg13g2_nor2b_2 _20079_ (.A(_11115_),
    .B_N(_11116_),
    .Y(_11117_));
 sg13g2_nand2b_2 _20080_ (.Y(_11118_),
    .B(_11116_),
    .A_N(_11115_));
 sg13g2_nor2_1 _20081_ (.A(_00236_),
    .B(_11067_),
    .Y(_11119_));
 sg13g2_a22oi_1 _20082_ (.Y(_11120_),
    .B1(_11059_),
    .B2(\soc_I.kianv_I.Instr[11] ),
    .A2(net8641),
    .A1(net9434));
 sg13g2_a221oi_1 _20083_ (.B2(net9709),
    .C1(_11119_),
    .B1(_11059_),
    .A1(net9434),
    .Y(_11121_),
    .A2(net8641));
 sg13g2_nand2b_1 _20084_ (.Y(_11122_),
    .B(_11120_),
    .A_N(_11119_));
 sg13g2_a21o_1 _20085_ (.A2(net8647),
    .A1(_00197_),
    .B1(net8637),
    .X(_11123_));
 sg13g2_a21oi_2 _20086_ (.B1(_11123_),
    .Y(_11124_),
    .A2(_11121_),
    .A1(net8643));
 sg13g2_a21o_1 _20087_ (.A2(_11121_),
    .A1(net8642),
    .B1(_11123_),
    .X(_11125_));
 sg13g2_xnor2_1 _20088_ (.Y(_11126_),
    .A(net8310),
    .B(net8449));
 sg13g2_nor2_1 _20089_ (.A(net8303),
    .B(_11126_),
    .Y(_11127_));
 sg13g2_xnor2_1 _20090_ (.Y(_11128_),
    .A(net8303),
    .B(_11126_));
 sg13g2_a221oi_1 _20091_ (.B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[3] ),
    .C1(net8714),
    .B1(net8653),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[3] ),
    .Y(_11129_),
    .A2(net8567));
 sg13g2_nor2_1 _20092_ (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[3] ),
    .B(net8719),
    .Y(_11130_));
 sg13g2_nand2_1 _20093_ (.Y(_11131_),
    .A(\soc_I.PC[3] ),
    .B(net8525));
 sg13g2_o21ai_1 _20094_ (.B1(_11131_),
    .Y(_11132_),
    .A1(_11129_),
    .A2(_11130_));
 sg13g2_nor2_1 _20095_ (.A(_00238_),
    .B(_11067_),
    .Y(_11133_));
 sg13g2_a221oi_1 _20096_ (.B2(\soc_I.kianv_I.Instr[10] ),
    .C1(_11133_),
    .B1(_11059_),
    .A1(net9442),
    .Y(_11134_),
    .A2(net8641));
 sg13g2_a21o_1 _20097_ (.A2(net8647),
    .A1(_00237_),
    .B1(net8636),
    .X(_11135_));
 sg13g2_a21oi_1 _20098_ (.A1(net8642),
    .A2(_11134_),
    .Y(_11136_),
    .B1(_11135_));
 sg13g2_a21o_1 _20099_ (.A2(_11134_),
    .A1(net8642),
    .B1(_11135_),
    .X(_11137_));
 sg13g2_xnor2_1 _20100_ (.Y(_11138_),
    .A(net8313),
    .B(net8438));
 sg13g2_nor2_1 _20101_ (.A(net8301),
    .B(_11138_),
    .Y(_11139_));
 sg13g2_a221oi_1 _20102_ (.B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[2] ),
    .C1(net8713),
    .B1(net8652),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[2] ),
    .Y(_11140_),
    .A2(net8566));
 sg13g2_a21oi_1 _20103_ (.A1(_10494_),
    .A2(net8713),
    .Y(_11141_),
    .B1(_11140_));
 sg13g2_nand2_1 _20104_ (.Y(_11142_),
    .A(\soc_I.PC[2] ),
    .B(net8526));
 sg13g2_nor2b_2 _20105_ (.A(_11141_),
    .B_N(_11142_),
    .Y(_11143_));
 sg13g2_nand2b_2 _20106_ (.Y(_11144_),
    .B(_11142_),
    .A_N(_11141_));
 sg13g2_a21oi_1 _20107_ (.A1(_00201_),
    .A2(net8639),
    .Y(_11145_),
    .B1(net8642));
 sg13g2_o21ai_1 _20108_ (.B1(\soc_I.kianv_I.Instr[9] ),
    .Y(_11146_),
    .A1(_11055_),
    .A2(_11058_));
 sg13g2_nand2b_1 _20109_ (.Y(_11147_),
    .B(_11066_),
    .A_N(_00215_));
 sg13g2_nand2_1 _20110_ (.Y(_11148_),
    .A(net9458),
    .B(net8641));
 sg13g2_and3_1 _20111_ (.X(_11149_),
    .A(_11146_),
    .B(_11147_),
    .C(_11148_));
 sg13g2_nand3_1 _20112_ (.B(_11147_),
    .C(_11148_),
    .A(_11146_),
    .Y(_11150_));
 sg13g2_nor2_1 _20113_ (.A(net8647),
    .B(net8636),
    .Y(_11151_));
 sg13g2_a21oi_2 _20114_ (.B1(_11145_),
    .Y(_11152_),
    .A2(_11151_),
    .A1(_11150_));
 sg13g2_a21o_1 _20115_ (.A2(_11151_),
    .A1(_11150_),
    .B1(_11145_),
    .X(_11153_));
 sg13g2_xnor2_1 _20116_ (.Y(_11154_),
    .A(net8310),
    .B(net8427));
 sg13g2_and2_1 _20117_ (.A(_11144_),
    .B(_11154_),
    .X(_11155_));
 sg13g2_a221oi_1 _20118_ (.B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[1] ),
    .C1(net8716),
    .B1(_10986_),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[1] ),
    .Y(_11156_),
    .A2(net8569));
 sg13g2_nor2_1 _20119_ (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[1] ),
    .B(net8722),
    .Y(_11157_));
 sg13g2_nand2_1 _20120_ (.Y(_11158_),
    .A(\soc_I.PC[1] ),
    .B(net8528));
 sg13g2_o21ai_1 _20121_ (.B1(_11158_),
    .Y(_11159_),
    .A1(_11156_),
    .A2(_11157_));
 sg13g2_inv_1 _20122_ (.Y(_11160_),
    .A(net8299));
 sg13g2_o21ai_1 _20123_ (.B1(\soc_I.kianv_I.Instr[8] ),
    .Y(_11161_),
    .A1(_11055_),
    .A2(_11058_));
 sg13g2_a22oi_1 _20124_ (.Y(_11162_),
    .B1(_11066_),
    .B2(_10590_),
    .A2(net8641),
    .A1(net9487));
 sg13g2_and2_2 _20125_ (.A(_11161_),
    .B(_11162_),
    .X(_11163_));
 sg13g2_nand2_2 _20126_ (.Y(_11164_),
    .A(_11161_),
    .B(_11162_));
 sg13g2_nand3_1 _20127_ (.B(_11161_),
    .C(_11162_),
    .A(net8643),
    .Y(_11165_));
 sg13g2_a21oi_2 _20128_ (.B1(net8636),
    .Y(_11166_),
    .A2(net8647),
    .A1(_00205_));
 sg13g2_a21o_1 _20129_ (.A2(net8646),
    .A1(_00205_),
    .B1(net8635),
    .X(_11167_));
 sg13g2_and2_1 _20130_ (.A(_11165_),
    .B(_11166_),
    .X(_11168_));
 sg13g2_nand2_1 _20131_ (.Y(_11169_),
    .A(_11165_),
    .B(_11166_));
 sg13g2_xnor2_1 _20132_ (.Y(_11170_),
    .A(net8310),
    .B(net8400));
 sg13g2_or2_1 _20133_ (.X(_11171_),
    .B(_11170_),
    .A(_11160_));
 sg13g2_xnor2_1 _20134_ (.Y(_11172_),
    .A(_11160_),
    .B(_11170_));
 sg13g2_and2_1 _20135_ (.A(\soc_I.kianv_I.Instr[7] ),
    .B(_11055_),
    .X(_11173_));
 sg13g2_a21oi_2 _20136_ (.B1(_11173_),
    .Y(_11174_),
    .A2(net8641),
    .A1(net9522));
 sg13g2_a21o_1 _20137_ (.A2(net8641),
    .A1(net9522),
    .B1(_11173_),
    .X(_11175_));
 sg13g2_nand2_1 _20138_ (.Y(_11176_),
    .A(net8642),
    .B(net8562));
 sg13g2_nand2b_1 _20139_ (.Y(_11177_),
    .B(net8647),
    .A_N(_00209_));
 sg13g2_and2_1 _20140_ (.A(_00209_),
    .B(net8644),
    .X(_11178_));
 sg13g2_a221oi_1 _20141_ (.B2(\soc_I.kianv_I.Instr[7] ),
    .C1(net8649),
    .B1(_11055_),
    .A1(net9522),
    .Y(_11179_),
    .A2(net8641));
 sg13g2_nor2_1 _20142_ (.A(_11178_),
    .B(_11179_),
    .Y(_11180_));
 sg13g2_nor3_1 _20143_ (.A(net8635),
    .B(_11178_),
    .C(_11179_),
    .Y(_11181_));
 sg13g2_nand2_1 _20144_ (.Y(_11182_),
    .A(net8639),
    .B(_11180_));
 sg13g2_a221oi_1 _20145_ (.B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[0] ),
    .C1(net8716),
    .B1(net8651),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[0] ),
    .Y(_11183_),
    .A2(net8565));
 sg13g2_a21oi_1 _20146_ (.A1(_10496_),
    .A2(net8712),
    .Y(_11184_),
    .B1(_11183_));
 sg13g2_a21oi_2 _20147_ (.B1(_11184_),
    .Y(_11185_),
    .A2(net8525),
    .A1(\soc_I.PC[0] ));
 sg13g2_inv_1 _20148_ (.Y(_11186_),
    .A(net8298));
 sg13g2_nand2_1 _20149_ (.Y(_11187_),
    .A(net8510),
    .B(_11185_));
 sg13g2_o21ai_1 _20150_ (.B1(_11187_),
    .Y(_11188_),
    .A1(net8312),
    .A2(net8510));
 sg13g2_o21ai_1 _20151_ (.B1(_11171_),
    .Y(_11189_),
    .A1(_11172_),
    .A2(_11188_));
 sg13g2_xnor2_1 _20152_ (.Y(_11190_),
    .A(_11144_),
    .B(_11154_));
 sg13g2_inv_1 _20153_ (.Y(_11191_),
    .A(_11190_));
 sg13g2_a21oi_1 _20154_ (.A1(_11189_),
    .A2(_11191_),
    .Y(_11192_),
    .B1(_11155_));
 sg13g2_a221oi_1 _20155_ (.B2(_11191_),
    .C1(_11155_),
    .B1(_11189_),
    .A1(net8301),
    .Y(_11193_),
    .A2(_11138_));
 sg13g2_nor3_2 _20156_ (.A(_11128_),
    .B(_11139_),
    .C(_11193_),
    .Y(_11194_));
 sg13g2_nor2_1 _20157_ (.A(_11127_),
    .B(_11194_),
    .Y(_11195_));
 sg13g2_nor3_1 _20158_ (.A(_11112_),
    .B(_11127_),
    .C(_11194_),
    .Y(_11196_));
 sg13g2_nor2_1 _20159_ (.A(_11113_),
    .B(_11196_),
    .Y(_11197_));
 sg13g2_o21ai_1 _20160_ (.B1(_11102_),
    .Y(_11198_),
    .A1(_11113_),
    .A2(_11196_));
 sg13g2_nand2_1 _20161_ (.Y(_11199_),
    .A(_11087_),
    .B(_11091_));
 sg13g2_nand2_1 _20162_ (.Y(_11200_),
    .A(_11097_),
    .B(_11101_));
 sg13g2_and2_1 _20163_ (.A(_11199_),
    .B(_11200_),
    .X(_11201_));
 sg13g2_a21o_2 _20164_ (.A2(_11201_),
    .A1(_11198_),
    .B1(_11092_),
    .X(_11202_));
 sg13g2_a22oi_1 _20165_ (.Y(_11203_),
    .B1(net8652),
    .B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[8] ),
    .A2(net8566),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[8] ));
 sg13g2_nor2_1 _20166_ (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[8] ),
    .B(net8720),
    .Y(_11204_));
 sg13g2_a21oi_1 _20167_ (.A1(net8720),
    .A2(_11203_),
    .Y(_11205_),
    .B1(_11204_));
 sg13g2_nand2_1 _20168_ (.Y(_11206_),
    .A(\soc_I.PC[8] ),
    .B(net8526));
 sg13g2_nor2b_2 _20169_ (.A(_11205_),
    .B_N(_11206_),
    .Y(_11207_));
 sg13g2_nand2b_2 _20170_ (.Y(_11208_),
    .B(_11206_),
    .A_N(_11205_));
 sg13g2_nand2_2 _20171_ (.Y(_11209_),
    .A(net9430),
    .B(net8711));
 sg13g2_inv_1 _20172_ (.Y(_11210_),
    .A(_11209_));
 sg13g2_a21o_1 _20173_ (.A2(net8646),
    .A1(_00211_),
    .B1(net8637),
    .X(_11211_));
 sg13g2_a21oi_2 _20174_ (.B1(_11211_),
    .Y(_11212_),
    .A2(_11209_),
    .A1(net8642));
 sg13g2_xnor2_1 _20175_ (.Y(_11213_),
    .A(net8312),
    .B(net8507));
 sg13g2_nor2_1 _20176_ (.A(_11207_),
    .B(_11213_),
    .Y(_11214_));
 sg13g2_xnor2_1 _20177_ (.Y(_11215_),
    .A(_11208_),
    .B(_11213_));
 sg13g2_inv_1 _20178_ (.Y(_11216_),
    .A(_11215_));
 sg13g2_a22oi_1 _20179_ (.Y(_11217_),
    .B1(net8652),
    .B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[10] ),
    .A2(net8566),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[10] ));
 sg13g2_nor2_1 _20180_ (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[10] ),
    .B(net8720),
    .Y(_11218_));
 sg13g2_a21oi_1 _20181_ (.A1(net8720),
    .A2(_11217_),
    .Y(_11219_),
    .B1(_11218_));
 sg13g2_nand2_1 _20182_ (.Y(_11220_),
    .A(\soc_I.PC[10] ),
    .B(net8526));
 sg13g2_nor2b_2 _20183_ (.A(_11219_),
    .B_N(_11220_),
    .Y(_11221_));
 sg13g2_nand2b_2 _20184_ (.Y(_11222_),
    .B(_11220_),
    .A_N(_11219_));
 sg13g2_o21ai_1 _20185_ (.B1(net8643),
    .Y(_11223_),
    .A1(_00213_),
    .A2(net8709));
 sg13g2_a21oi_1 _20186_ (.A1(_00203_),
    .A2(net8647),
    .Y(_11224_),
    .B1(net8635));
 sg13g2_and2_1 _20187_ (.A(_11223_),
    .B(_11224_),
    .X(_11225_));
 sg13g2_xnor2_1 _20188_ (.Y(_11226_),
    .A(net8310),
    .B(net8506));
 sg13g2_nor2_1 _20189_ (.A(_11221_),
    .B(_11226_),
    .Y(_11227_));
 sg13g2_or2_1 _20190_ (.X(_11228_),
    .B(_11226_),
    .A(_11221_));
 sg13g2_xnor2_1 _20191_ (.Y(_11229_),
    .A(_11221_),
    .B(_11226_));
 sg13g2_inv_1 _20192_ (.Y(_11230_),
    .A(_11229_));
 sg13g2_a221oi_1 _20193_ (.B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[11] ),
    .C1(net8712),
    .B1(net8650),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[11] ),
    .Y(_11231_),
    .A2(net8564));
 sg13g2_nor2_1 _20194_ (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[11] ),
    .B(net8719),
    .Y(_11232_));
 sg13g2_nand2_1 _20195_ (.Y(_11233_),
    .A(\soc_I.PC[11] ),
    .B(net8524));
 sg13g2_o21ai_1 _20196_ (.B1(_11233_),
    .Y(_11234_),
    .A1(_11231_),
    .A2(_11232_));
 sg13g2_o21ai_1 _20197_ (.B1(_11014_),
    .Y(_11235_),
    .A1(net9132),
    .A2(_11067_));
 sg13g2_a221oi_1 _20198_ (.B2(\soc_I.kianv_I.Instr[7] ),
    .C1(_11235_),
    .B1(_11058_),
    .A1(net9424),
    .Y(_11236_),
    .A2(_11055_));
 sg13g2_a21o_1 _20199_ (.A2(net8649),
    .A1(_00234_),
    .B1(net8637),
    .X(_11237_));
 sg13g2_a21oi_2 _20200_ (.B1(_11237_),
    .Y(_11238_),
    .A2(_11236_),
    .A1(net8643));
 sg13g2_xnor2_1 _20201_ (.Y(_11239_),
    .A(net8313),
    .B(net8382));
 sg13g2_nor2_1 _20202_ (.A(net8296),
    .B(_11239_),
    .Y(_11240_));
 sg13g2_xnor2_1 _20203_ (.Y(_11241_),
    .A(net8296),
    .B(_11239_));
 sg13g2_a22oi_1 _20204_ (.Y(_11242_),
    .B1(net8653),
    .B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[9] ),
    .A2(net8567),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[9] ));
 sg13g2_nor2_1 _20205_ (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[9] ),
    .B(net8720),
    .Y(_11243_));
 sg13g2_a21oi_1 _20206_ (.A1(net8720),
    .A2(_11242_),
    .Y(_11244_),
    .B1(_11243_));
 sg13g2_nand2_1 _20207_ (.Y(_11245_),
    .A(\soc_I.PC[9] ),
    .B(net8526));
 sg13g2_nor2b_2 _20208_ (.A(_11244_),
    .B_N(_11245_),
    .Y(_11246_));
 sg13g2_nand2b_2 _20209_ (.Y(_11247_),
    .B(_11245_),
    .A_N(_11244_));
 sg13g2_a21oi_1 _20210_ (.A1(net9429),
    .A2(_11063_),
    .Y(_11248_),
    .B1(net8646));
 sg13g2_a21oi_1 _20211_ (.A1(_00207_),
    .A2(net8646),
    .Y(_11249_),
    .B1(net8635));
 sg13g2_nor2b_1 _20212_ (.A(_11248_),
    .B_N(_11249_),
    .Y(_11250_));
 sg13g2_xnor2_1 _20213_ (.Y(_11251_),
    .A(net8310),
    .B(net8505));
 sg13g2_nand2_1 _20214_ (.Y(_11252_),
    .A(_11246_),
    .B(_11251_));
 sg13g2_or2_1 _20215_ (.X(_11253_),
    .B(_11251_),
    .A(_11246_));
 sg13g2_nand2_1 _20216_ (.Y(_11254_),
    .A(_11252_),
    .B(_11253_));
 sg13g2_nor4_2 _20217_ (.A(_11216_),
    .B(_11229_),
    .C(_11241_),
    .Y(_11255_),
    .D(_11254_));
 sg13g2_nand2b_1 _20218_ (.Y(_11256_),
    .B(_11253_),
    .A_N(_11214_));
 sg13g2_nand2_1 _20219_ (.Y(_11257_),
    .A(_11252_),
    .B(_11256_));
 sg13g2_nor3_1 _20220_ (.A(_11229_),
    .B(_11241_),
    .C(_11257_),
    .Y(_11258_));
 sg13g2_a21oi_1 _20221_ (.A1(net8296),
    .A2(_11239_),
    .Y(_11259_),
    .B1(_11258_));
 sg13g2_o21ai_1 _20222_ (.B1(_11259_),
    .Y(_11260_),
    .A1(_11228_),
    .A2(_11240_));
 sg13g2_a21oi_2 _20223_ (.B1(_11260_),
    .Y(_11261_),
    .A2(_11255_),
    .A1(_11202_));
 sg13g2_a21o_1 _20224_ (.A2(_11255_),
    .A1(_11202_),
    .B1(_11260_),
    .X(_11262_));
 sg13g2_a22oi_1 _20225_ (.Y(_11263_),
    .B1(net8651),
    .B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[14] ),
    .A2(net8565),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[14] ));
 sg13g2_nor2_1 _20226_ (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[14] ),
    .B(net8718),
    .Y(_11264_));
 sg13g2_a21oi_1 _20227_ (.A1(net8719),
    .A2(_11263_),
    .Y(_11265_),
    .B1(_11264_));
 sg13g2_nand2_1 _20228_ (.Y(_11266_),
    .A(\soc_I.PC[14] ),
    .B(net8525));
 sg13g2_nor2b_2 _20229_ (.A(_11265_),
    .B_N(_11266_),
    .Y(_11267_));
 sg13g2_nand2b_2 _20230_ (.Y(_11268_),
    .B(_11266_),
    .A_N(_11265_));
 sg13g2_nand2_2 _20231_ (.Y(_11269_),
    .A(_11063_),
    .B(_11067_));
 sg13g2_nand2_1 _20232_ (.Y(_11270_),
    .A(net9698),
    .B(_11269_));
 sg13g2_a22oi_1 _20233_ (.Y(_11271_),
    .B1(net8523),
    .B2(_11270_),
    .A2(net8645),
    .A1(_00191_));
 sg13g2_and2_2 _20234_ (.A(net8639),
    .B(_11271_),
    .X(_11272_));
 sg13g2_nand2_2 _20235_ (.Y(_11273_),
    .A(net8638),
    .B(_11271_));
 sg13g2_xnor2_1 _20236_ (.Y(_11274_),
    .A(net8311),
    .B(_11272_));
 sg13g2_nor2_1 _20237_ (.A(_11267_),
    .B(_11274_),
    .Y(_11275_));
 sg13g2_xnor2_1 _20238_ (.Y(_11276_),
    .A(net8295),
    .B(_11274_));
 sg13g2_a221oi_1 _20239_ (.B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[15] ),
    .C1(net8712),
    .B1(net8650),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[15] ),
    .Y(_11277_),
    .A2(net8564));
 sg13g2_nor2_1 _20240_ (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[15] ),
    .B(net8717),
    .Y(_11278_));
 sg13g2_nand2_1 _20241_ (.Y(_11279_),
    .A(\soc_I.PC[15] ),
    .B(net8525));
 sg13g2_o21ai_1 _20242_ (.B1(_11279_),
    .Y(_11280_),
    .A1(_11277_),
    .A2(_11278_));
 sg13g2_nand2_1 _20243_ (.Y(_11281_),
    .A(net9663),
    .B(_11269_));
 sg13g2_a221oi_1 _20244_ (.B2(_11281_),
    .C1(net8635),
    .B1(net8523),
    .A1(_00233_),
    .Y(_11282_),
    .A2(net8645));
 sg13g2_xnor2_1 _20245_ (.Y(_11283_),
    .A(net8313),
    .B(net8381));
 sg13g2_nand2_1 _20246_ (.Y(_11284_),
    .A(net8293),
    .B(_11283_));
 sg13g2_or2_1 _20247_ (.X(_11285_),
    .B(_11283_),
    .A(net8293));
 sg13g2_nand2_1 _20248_ (.Y(_11286_),
    .A(_11284_),
    .B(_11285_));
 sg13g2_nor2_1 _20249_ (.A(_11276_),
    .B(_11286_),
    .Y(_11287_));
 sg13g2_a221oi_1 _20250_ (.B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[12] ),
    .C1(net8713),
    .B1(net8652),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[12] ),
    .Y(_11288_),
    .A2(net8566));
 sg13g2_nor2_1 _20251_ (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[12] ),
    .B(net8720),
    .Y(_11289_));
 sg13g2_nand2_1 _20252_ (.Y(_11290_),
    .A(\soc_I.PC[12] ),
    .B(net8526));
 sg13g2_o21ai_1 _20253_ (.B1(_11290_),
    .Y(_11291_),
    .A1(_11288_),
    .A2(_11289_));
 sg13g2_inv_2 _20254_ (.Y(_11292_),
    .A(net8292));
 sg13g2_nand2_1 _20255_ (.Y(_11293_),
    .A(net9706),
    .B(_11269_));
 sg13g2_a221oi_1 _20256_ (.B2(_11293_),
    .C1(net8636),
    .B1(net8523),
    .A1(_00199_),
    .Y(_11294_),
    .A2(net8644));
 sg13g2_xnor2_1 _20257_ (.Y(_11295_),
    .A(net8310),
    .B(net8380));
 sg13g2_or2_1 _20258_ (.X(_11296_),
    .B(_11295_),
    .A(_11292_));
 sg13g2_xnor2_1 _20259_ (.Y(_11297_),
    .A(_11292_),
    .B(_11295_));
 sg13g2_inv_1 _20260_ (.Y(_11298_),
    .A(_11297_));
 sg13g2_a22oi_1 _20261_ (.Y(_11299_),
    .B1(net8654),
    .B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[13] ),
    .A2(net8568),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[13] ));
 sg13g2_nor2_1 _20262_ (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[13] ),
    .B(net8721),
    .Y(_11300_));
 sg13g2_a21oi_1 _20263_ (.A1(net8722),
    .A2(_11299_),
    .Y(_11301_),
    .B1(_11300_));
 sg13g2_nand2_1 _20264_ (.Y(_11302_),
    .A(\soc_I.PC[13] ),
    .B(net8527));
 sg13g2_nor2b_2 _20265_ (.A(_11301_),
    .B_N(_11302_),
    .Y(_11303_));
 sg13g2_nand2b_2 _20266_ (.Y(_11304_),
    .B(_11302_),
    .A_N(_11301_));
 sg13g2_nand2_1 _20267_ (.Y(_11305_),
    .A(net9703),
    .B(_11269_));
 sg13g2_a22oi_1 _20268_ (.Y(_11306_),
    .B1(net8523),
    .B2(_11305_),
    .A2(net8645),
    .A1(_00195_));
 sg13g2_nand2_2 _20269_ (.Y(_11307_),
    .A(net8640),
    .B(_11306_));
 sg13g2_inv_2 _20270_ (.Y(_11308_),
    .A(net8290));
 sg13g2_xnor2_1 _20271_ (.Y(_11309_),
    .A(net8310),
    .B(net8290));
 sg13g2_or2_1 _20272_ (.X(_11310_),
    .B(_11309_),
    .A(_11304_));
 sg13g2_inv_1 _20273_ (.Y(_11311_),
    .A(_11310_));
 sg13g2_nand2_1 _20274_ (.Y(_11312_),
    .A(_11304_),
    .B(_11309_));
 sg13g2_nand2_1 _20275_ (.Y(_11313_),
    .A(_11310_),
    .B(_11312_));
 sg13g2_nand4_1 _20276_ (.B(_11298_),
    .C(_11310_),
    .A(_11287_),
    .Y(_11314_),
    .D(_11312_));
 sg13g2_nand2_1 _20277_ (.Y(_11315_),
    .A(_11296_),
    .B(_11312_));
 sg13g2_nand3_1 _20278_ (.B(_11310_),
    .C(_11315_),
    .A(_11287_),
    .Y(_11316_));
 sg13g2_nand2_1 _20279_ (.Y(_11317_),
    .A(_11275_),
    .B(_11285_));
 sg13g2_and3_1 _20280_ (.X(_11318_),
    .A(_11284_),
    .B(_11316_),
    .C(_11317_));
 sg13g2_o21ai_1 _20281_ (.B1(_11318_),
    .Y(_11319_),
    .A1(_11261_),
    .A2(_11314_));
 sg13g2_a221oi_1 _20282_ (.B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[22] ),
    .C1(net8715),
    .B1(net8654),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[22] ),
    .Y(_11320_),
    .A2(net8568));
 sg13g2_a21oi_1 _20283_ (.A1(_10479_),
    .A2(net8715),
    .Y(_11321_),
    .B1(_11320_));
 sg13g2_a21oi_1 _20284_ (.A1(\soc_I.PC[22] ),
    .A2(net8527),
    .Y(_11322_),
    .B1(_11321_));
 sg13g2_inv_2 _20285_ (.Y(_11323_),
    .A(net8288));
 sg13g2_nand2_1 _20286_ (.Y(_11324_),
    .A(net9462),
    .B(net8710));
 sg13g2_a22oi_1 _20287_ (.Y(_11325_),
    .B1(net8309),
    .B2(_11324_),
    .A2(net8648),
    .A1(_00226_));
 sg13g2_nand2_2 _20288_ (.Y(_11326_),
    .A(net8638),
    .B(_11325_));
 sg13g2_inv_1 _20289_ (.Y(_11327_),
    .A(_11326_));
 sg13g2_xnor2_1 _20290_ (.Y(_11328_),
    .A(_11042_),
    .B(_11326_));
 sg13g2_nor2_1 _20291_ (.A(net8288),
    .B(_11328_),
    .Y(_11329_));
 sg13g2_inv_1 _20292_ (.Y(_11330_),
    .A(_11329_));
 sg13g2_xnor2_1 _20293_ (.Y(_11331_),
    .A(net8288),
    .B(_11328_));
 sg13g2_a221oi_1 _20294_ (.B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[23] ),
    .C1(net8712),
    .B1(net8650),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[23] ),
    .Y(_11332_),
    .A2(net8564));
 sg13g2_nor2_1 _20295_ (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[23] ),
    .B(net8718),
    .Y(_11333_));
 sg13g2_nand2_1 _20296_ (.Y(_11334_),
    .A(\soc_I.PC[23] ),
    .B(net8524));
 sg13g2_o21ai_1 _20297_ (.B1(_11334_),
    .Y(_11335_),
    .A1(_11332_),
    .A2(_11333_));
 sg13g2_inv_1 _20298_ (.Y(_11336_),
    .A(net8287));
 sg13g2_nand2_1 _20299_ (.Y(_11337_),
    .A(net9444),
    .B(net8710));
 sg13g2_a22oi_1 _20300_ (.Y(_11338_),
    .B1(_11068_),
    .B2(_11337_),
    .A2(net8648),
    .A1(_00225_));
 sg13g2_nand2_2 _20301_ (.Y(_11339_),
    .A(net8638),
    .B(_11338_));
 sg13g2_inv_1 _20302_ (.Y(_11340_),
    .A(_11339_));
 sg13g2_xnor2_1 _20303_ (.Y(_11341_),
    .A(net8313),
    .B(_11339_));
 sg13g2_nor2_1 _20304_ (.A(_11336_),
    .B(_11341_),
    .Y(_11342_));
 sg13g2_nand2_1 _20305_ (.Y(_11343_),
    .A(_11336_),
    .B(_11341_));
 sg13g2_nand2b_1 _20306_ (.Y(_11344_),
    .B(_11343_),
    .A_N(_11342_));
 sg13g2_nor2_1 _20307_ (.A(_11331_),
    .B(_11344_),
    .Y(_11345_));
 sg13g2_a22oi_1 _20308_ (.Y(_11346_),
    .B1(net8653),
    .B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[20] ),
    .A2(net8567),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[20] ));
 sg13g2_nor2_1 _20309_ (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[20] ),
    .B(net8721),
    .Y(_11347_));
 sg13g2_a21oi_1 _20310_ (.A1(net8721),
    .A2(_11346_),
    .Y(_11348_),
    .B1(_11347_));
 sg13g2_a21oi_2 _20311_ (.B1(_11348_),
    .Y(_11349_),
    .A2(net8527),
    .A1(\soc_I.PC[20] ));
 sg13g2_inv_2 _20312_ (.Y(_11350_),
    .A(net8286));
 sg13g2_nand2_1 _20313_ (.Y(_11351_),
    .A(net9527),
    .B(net8710));
 sg13g2_a22oi_1 _20314_ (.Y(_11352_),
    .B1(net8309),
    .B2(_11351_),
    .A2(net8648),
    .A1(_00228_));
 sg13g2_and2_2 _20315_ (.A(net8638),
    .B(_11352_),
    .X(_11353_));
 sg13g2_nand2_2 _20316_ (.Y(_11354_),
    .A(net8638),
    .B(_11352_));
 sg13g2_xnor2_1 _20317_ (.Y(_11355_),
    .A(net8312),
    .B(_11353_));
 sg13g2_or2_1 _20318_ (.X(_11356_),
    .B(_11355_),
    .A(net8286));
 sg13g2_xnor2_1 _20319_ (.Y(_11357_),
    .A(_11350_),
    .B(_11355_));
 sg13g2_inv_1 _20320_ (.Y(_11358_),
    .A(_11357_));
 sg13g2_a221oi_1 _20321_ (.B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[21] ),
    .C1(net8714),
    .B1(net8654),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[21] ),
    .Y(_11359_),
    .A2(net8568));
 sg13g2_nor2_1 _20322_ (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[21] ),
    .B(net8721),
    .Y(_11360_));
 sg13g2_nand2_1 _20323_ (.Y(_11361_),
    .A(\soc_I.PC[21] ),
    .B(net8527));
 sg13g2_o21ai_1 _20324_ (.B1(_11361_),
    .Y(_11362_),
    .A1(_11359_),
    .A2(_11360_));
 sg13g2_nand2_1 _20325_ (.Y(_11363_),
    .A(net9491),
    .B(net8710));
 sg13g2_a22oi_1 _20326_ (.Y(_11364_),
    .B1(_11068_),
    .B2(_11363_),
    .A2(net8648),
    .A1(_00227_));
 sg13g2_and2_2 _20327_ (.A(net8639),
    .B(_11364_),
    .X(_11365_));
 sg13g2_nand2_2 _20328_ (.Y(_11366_),
    .A(net8638),
    .B(_11364_));
 sg13g2_xnor2_1 _20329_ (.Y(_11367_),
    .A(net8313),
    .B(_11365_));
 sg13g2_or2_1 _20330_ (.X(_11368_),
    .B(_11367_),
    .A(net8284));
 sg13g2_nand2_1 _20331_ (.Y(_11369_),
    .A(net8284),
    .B(_11367_));
 sg13g2_inv_1 _20332_ (.Y(_11370_),
    .A(_11369_));
 sg13g2_nand2_1 _20333_ (.Y(_11371_),
    .A(_11368_),
    .B(_11369_));
 sg13g2_inv_1 _20334_ (.Y(_11372_),
    .A(_11371_));
 sg13g2_nand3_1 _20335_ (.B(_11357_),
    .C(_11372_),
    .A(_11345_),
    .Y(_11373_));
 sg13g2_a22oi_1 _20336_ (.Y(_11374_),
    .B1(net8650),
    .B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[16] ),
    .A2(net8564),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[16] ));
 sg13g2_nor2_1 _20337_ (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[16] ),
    .B(net8717),
    .Y(_11375_));
 sg13g2_a21oi_1 _20338_ (.A1(net8718),
    .A2(_11374_),
    .Y(_11376_),
    .B1(_11375_));
 sg13g2_nand2_1 _20339_ (.Y(_11377_),
    .A(\led[0] ),
    .B(net8524));
 sg13g2_nor2b_2 _20340_ (.A(_11376_),
    .B_N(_11377_),
    .Y(_11378_));
 sg13g2_nand2b_2 _20341_ (.Y(_11379_),
    .B(_11377_),
    .A_N(_11376_));
 sg13g2_nand2_1 _20342_ (.Y(_11380_),
    .A(net9606),
    .B(_11269_));
 sg13g2_a22oi_1 _20343_ (.Y(_11381_),
    .B1(net8523),
    .B2(_11380_),
    .A2(net8644),
    .A1(_00232_));
 sg13g2_and2_1 _20344_ (.A(net8639),
    .B(_11381_),
    .X(_11382_));
 sg13g2_nand2_2 _20345_ (.Y(_11383_),
    .A(net8639),
    .B(_11381_));
 sg13g2_xnor2_1 _20346_ (.Y(_11384_),
    .A(net8311),
    .B(_11382_));
 sg13g2_nor2_1 _20347_ (.A(_11378_),
    .B(_11384_),
    .Y(_11385_));
 sg13g2_xnor2_1 _20348_ (.Y(_11386_),
    .A(_11379_),
    .B(_11384_));
 sg13g2_xnor2_1 _20349_ (.Y(_11387_),
    .A(net8283),
    .B(_11384_));
 sg13g2_a22oi_1 _20350_ (.Y(_11388_),
    .B1(net8650),
    .B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[18] ),
    .A2(net8564),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[18] ));
 sg13g2_nor2_1 _20351_ (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[18] ),
    .B(net8717),
    .Y(_11389_));
 sg13g2_a21oi_1 _20352_ (.A1(net8717),
    .A2(_11388_),
    .Y(_11390_),
    .B1(_11389_));
 sg13g2_a21oi_1 _20353_ (.A1(\led[2] ),
    .A2(net8524),
    .Y(_11391_),
    .B1(_11390_));
 sg13g2_inv_1 _20354_ (.Y(_11392_),
    .A(net8281));
 sg13g2_nand2_1 _20355_ (.Y(_11393_),
    .A(net9555),
    .B(_11269_));
 sg13g2_a221oi_1 _20356_ (.B2(_11393_),
    .C1(net8635),
    .B1(net8523),
    .A1(_00230_),
    .Y(_11394_),
    .A2(net8644));
 sg13g2_xnor2_1 _20357_ (.Y(_11395_),
    .A(net8312),
    .B(net8379));
 sg13g2_nor2_1 _20358_ (.A(net8281),
    .B(_11395_),
    .Y(_11396_));
 sg13g2_xnor2_1 _20359_ (.Y(_11397_),
    .A(net8281),
    .B(_11395_));
 sg13g2_a221oi_1 _20360_ (.B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[19] ),
    .C1(net8712),
    .B1(net8651),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[19] ),
    .Y(_11398_),
    .A2(net8565));
 sg13g2_nor2_1 _20361_ (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[19] ),
    .B(net8717),
    .Y(_11399_));
 sg13g2_nand2_1 _20362_ (.Y(_11400_),
    .A(\led[3] ),
    .B(net8524));
 sg13g2_o21ai_1 _20363_ (.B1(_11400_),
    .Y(_11401_),
    .A1(_11398_),
    .A2(_11399_));
 sg13g2_inv_1 _20364_ (.Y(_11402_),
    .A(net8279));
 sg13g2_nand2_1 _20365_ (.Y(_11403_),
    .A(net9547),
    .B(_11269_));
 sg13g2_a221oi_1 _20366_ (.B2(_11403_),
    .C1(net8635),
    .B1(net8523),
    .A1(_00229_),
    .Y(_11404_),
    .A2(net8644));
 sg13g2_xnor2_1 _20367_ (.Y(_11405_),
    .A(_11042_),
    .B(_11404_));
 sg13g2_nand2_1 _20368_ (.Y(_11406_),
    .A(net8280),
    .B(_11405_));
 sg13g2_or2_1 _20369_ (.X(_11407_),
    .B(_11405_),
    .A(net8280));
 sg13g2_nand2_1 _20370_ (.Y(_11408_),
    .A(_11406_),
    .B(_11407_));
 sg13g2_nor2_1 _20371_ (.A(_11397_),
    .B(_11408_),
    .Y(_11409_));
 sg13g2_a221oi_1 _20372_ (.B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[17] ),
    .C1(net8712),
    .B1(net8650),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[17] ),
    .Y(_11410_),
    .A2(net8564));
 sg13g2_nor2_1 _20373_ (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[17] ),
    .B(net8717),
    .Y(_11411_));
 sg13g2_nand2_1 _20374_ (.Y(_11412_),
    .A(\led[1] ),
    .B(net8524));
 sg13g2_o21ai_1 _20375_ (.B1(_11412_),
    .Y(_11413_),
    .A1(_11410_),
    .A2(_11411_));
 sg13g2_nand2_1 _20376_ (.Y(_11414_),
    .A(net9568),
    .B(_11269_));
 sg13g2_a22oi_1 _20377_ (.Y(_11415_),
    .B1(_11060_),
    .B2(_11414_),
    .A2(net8644),
    .A1(_00231_));
 sg13g2_nand2_2 _20378_ (.Y(_11416_),
    .A(net8639),
    .B(_11415_));
 sg13g2_inv_1 _20379_ (.Y(_11417_),
    .A(_11416_));
 sg13g2_xnor2_1 _20380_ (.Y(_11418_),
    .A(net8312),
    .B(_11416_));
 sg13g2_nand2_1 _20381_ (.Y(_11419_),
    .A(net8277),
    .B(_11418_));
 sg13g2_nor2_1 _20382_ (.A(net8277),
    .B(_11418_),
    .Y(_11420_));
 sg13g2_or2_1 _20383_ (.X(_11421_),
    .B(_11418_),
    .A(net8276));
 sg13g2_nand2_1 _20384_ (.Y(_11422_),
    .A(_11419_),
    .B(_11421_));
 sg13g2_nor4_1 _20385_ (.A(_11387_),
    .B(_11397_),
    .C(_11408_),
    .D(_11422_),
    .Y(_11423_));
 sg13g2_nor2b_1 _20386_ (.A(_11373_),
    .B_N(_11423_),
    .Y(_11424_));
 sg13g2_nand2b_1 _20387_ (.Y(_11425_),
    .B(_11419_),
    .A_N(_11385_));
 sg13g2_nand3_1 _20388_ (.B(_11421_),
    .C(_11425_),
    .A(_11409_),
    .Y(_11426_));
 sg13g2_nand2_1 _20389_ (.Y(_11427_),
    .A(_11396_),
    .B(_11407_));
 sg13g2_nand3_1 _20390_ (.B(_11426_),
    .C(_11427_),
    .A(_11406_),
    .Y(_11428_));
 sg13g2_nand2b_1 _20391_ (.Y(_11429_),
    .B(_11428_),
    .A_N(_11373_));
 sg13g2_o21ai_1 _20392_ (.B1(_11343_),
    .Y(_11430_),
    .A1(_11329_),
    .A2(_11342_));
 sg13g2_nand2_1 _20393_ (.Y(_11431_),
    .A(_11356_),
    .B(_11369_));
 sg13g2_nand3_1 _20394_ (.B(_11368_),
    .C(_11431_),
    .A(_11345_),
    .Y(_11432_));
 sg13g2_nand3_1 _20395_ (.B(_11430_),
    .C(_11432_),
    .A(_11429_),
    .Y(_11433_));
 sg13g2_a21oi_2 _20396_ (.B1(_11433_),
    .Y(_11434_),
    .A2(_11424_),
    .A1(_11319_));
 sg13g2_a22oi_1 _20397_ (.Y(_11435_),
    .B1(net8654),
    .B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[26] ),
    .A2(net8568),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[26] ));
 sg13g2_nor2_1 _20398_ (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[26] ),
    .B(net8721),
    .Y(_11436_));
 sg13g2_a21oi_1 _20399_ (.A1(net8721),
    .A2(_11435_),
    .Y(_11437_),
    .B1(_11436_));
 sg13g2_nand2_1 _20400_ (.Y(_11438_),
    .A(\soc_I.PC[26] ),
    .B(net8527));
 sg13g2_nor2b_2 _20401_ (.A(_11437_),
    .B_N(_11438_),
    .Y(_11439_));
 sg13g2_nand2b_2 _20402_ (.Y(_11440_),
    .B(_11438_),
    .A_N(_11437_));
 sg13g2_nand2_1 _20403_ (.Y(_11441_),
    .A(\soc_I.kianv_I.Instr[26] ),
    .B(net8709));
 sg13g2_a221oi_1 _20404_ (.B2(_11441_),
    .C1(net8637),
    .B1(net8309),
    .A1(_00222_),
    .Y(_11442_),
    .A2(net8645));
 sg13g2_xnor2_1 _20405_ (.Y(_11443_),
    .A(net8311),
    .B(net8006));
 sg13g2_nor2_1 _20406_ (.A(net8275),
    .B(_11443_),
    .Y(_11444_));
 sg13g2_inv_1 _20407_ (.Y(_11445_),
    .A(_11444_));
 sg13g2_xnor2_1 _20408_ (.Y(_11446_),
    .A(net8275),
    .B(_11443_));
 sg13g2_a221oi_1 _20409_ (.B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[27] ),
    .C1(net8712),
    .B1(net8651),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[27] ),
    .Y(_11447_),
    .A2(net8565));
 sg13g2_nor2_1 _20410_ (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[27] ),
    .B(net8719),
    .Y(_11448_));
 sg13g2_nand2_1 _20411_ (.Y(_11449_),
    .A(\soc_I.PC[27] ),
    .B(net8528));
 sg13g2_o21ai_1 _20412_ (.B1(_11449_),
    .Y(_11450_),
    .A1(_11447_),
    .A2(_11448_));
 sg13g2_nand2_1 _20413_ (.Y(_11451_),
    .A(net9431),
    .B(net8709));
 sg13g2_a22oi_1 _20414_ (.Y(_11452_),
    .B1(net8309),
    .B2(_11451_),
    .A2(net8649),
    .A1(_00221_));
 sg13g2_nand2_2 _20415_ (.Y(_11453_),
    .A(net8640),
    .B(_11452_));
 sg13g2_inv_1 _20416_ (.Y(_11454_),
    .A(_11453_));
 sg13g2_xnor2_1 _20417_ (.Y(_11455_),
    .A(net8311),
    .B(_11453_));
 sg13g2_or2_1 _20418_ (.X(_11456_),
    .B(_11455_),
    .A(net8273));
 sg13g2_nand2_1 _20419_ (.Y(_11457_),
    .A(net8273),
    .B(_11455_));
 sg13g2_nand2_1 _20420_ (.Y(_11458_),
    .A(_11456_),
    .B(_11457_));
 sg13g2_nor2_1 _20421_ (.A(_11446_),
    .B(_11458_),
    .Y(_11459_));
 sg13g2_a221oi_1 _20422_ (.B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[24] ),
    .C1(net8713),
    .B1(net8652),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[24] ),
    .Y(_11460_),
    .A2(net8566));
 sg13g2_a21oi_1 _20423_ (.A1(_10477_),
    .A2(net8715),
    .Y(_11461_),
    .B1(_11460_));
 sg13g2_a21oi_1 _20424_ (.A1(\soc_I.PC[24] ),
    .A2(net8527),
    .Y(_11462_),
    .B1(_11461_));
 sg13g2_inv_4 _20425_ (.A(net8272),
    .Y(_11463_));
 sg13g2_nand2_1 _20426_ (.Y(_11464_),
    .A(net9435),
    .B(net8709));
 sg13g2_a221oi_1 _20427_ (.B2(_11464_),
    .C1(net8636),
    .B1(_11068_),
    .A1(_00224_),
    .Y(_11465_),
    .A2(net8648));
 sg13g2_xnor2_1 _20428_ (.Y(_11466_),
    .A(net8311),
    .B(_11465_));
 sg13g2_or2_1 _20429_ (.X(_11467_),
    .B(_11466_),
    .A(net8271));
 sg13g2_xnor2_1 _20430_ (.Y(_11468_),
    .A(net8271),
    .B(_11466_));
 sg13g2_inv_1 _20431_ (.Y(_11469_),
    .A(_11468_));
 sg13g2_a221oi_1 _20432_ (.B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[25] ),
    .C1(net8715),
    .B1(net8654),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[25] ),
    .Y(_11470_),
    .A2(net8568));
 sg13g2_a21oi_1 _20433_ (.A1(_10476_),
    .A2(net8715),
    .Y(_11471_),
    .B1(_11470_));
 sg13g2_a21oi_2 _20434_ (.B1(_11471_),
    .Y(_11472_),
    .A2(net8527),
    .A1(\soc_I.PC[25] ));
 sg13g2_inv_1 _20435_ (.Y(_11473_),
    .A(_11472_));
 sg13g2_nand2_1 _20436_ (.Y(_11474_),
    .A(\soc_I.kianv_I.Instr[25] ),
    .B(net8710));
 sg13g2_a22oi_1 _20437_ (.Y(_11475_),
    .B1(net8309),
    .B2(_11474_),
    .A2(net8648),
    .A1(_00223_));
 sg13g2_and2_2 _20438_ (.A(net8638),
    .B(_11475_),
    .X(_11476_));
 sg13g2_nand2_2 _20439_ (.Y(_11477_),
    .A(net8638),
    .B(_11475_));
 sg13g2_xnor2_1 _20440_ (.Y(_11478_),
    .A(net8311),
    .B(_11476_));
 sg13g2_nand2_2 _20441_ (.Y(_11479_),
    .A(net8270),
    .B(_11478_));
 sg13g2_or2_1 _20442_ (.X(_11480_),
    .B(_11478_),
    .A(net8270));
 sg13g2_nand2_1 _20443_ (.Y(_11481_),
    .A(_11479_),
    .B(_11480_));
 sg13g2_nand4_1 _20444_ (.B(_11469_),
    .C(_11479_),
    .A(_11459_),
    .Y(_11482_),
    .D(_11480_));
 sg13g2_nand2_1 _20445_ (.Y(_11483_),
    .A(_11467_),
    .B(_11480_));
 sg13g2_inv_1 _20446_ (.Y(_11484_),
    .A(_11483_));
 sg13g2_nand3_1 _20447_ (.B(_11479_),
    .C(_11483_),
    .A(_11459_),
    .Y(_11485_));
 sg13g2_nand2_1 _20448_ (.Y(_11486_),
    .A(_11457_),
    .B(_11485_));
 sg13g2_a21oi_1 _20449_ (.A1(_11444_),
    .A2(_11456_),
    .Y(_11487_),
    .B1(_11486_));
 sg13g2_o21ai_1 _20450_ (.B1(_11487_),
    .Y(_11488_),
    .A1(_11434_),
    .A2(_11482_));
 sg13g2_a221oi_1 _20451_ (.B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[28] ),
    .C1(net8714),
    .B1(net8653),
    .A1(\soc_I.kianv_I.datapath_unit_I.A1[28] ),
    .Y(_11489_),
    .A2(net8567));
 sg13g2_a21oi_1 _20452_ (.A1(_10473_),
    .A2(net8716),
    .Y(_11490_),
    .B1(_11489_));
 sg13g2_a21oi_1 _20453_ (.A1(\soc_I.PC[28] ),
    .A2(net8528),
    .Y(_11491_),
    .B1(_11490_));
 sg13g2_inv_2 _20454_ (.Y(_11492_),
    .A(net8268));
 sg13g2_nand2_1 _20455_ (.Y(_11493_),
    .A(\soc_I.kianv_I.Instr[28] ),
    .B(net8709));
 sg13g2_a22oi_1 _20456_ (.Y(_11494_),
    .B1(net8309),
    .B2(_11493_),
    .A2(net8649),
    .A1(_00220_));
 sg13g2_nand2_2 _20457_ (.Y(_11495_),
    .A(net8640),
    .B(_11494_));
 sg13g2_inv_1 _20458_ (.Y(_11496_),
    .A(_11495_));
 sg13g2_xnor2_1 _20459_ (.Y(_11497_),
    .A(net8313),
    .B(_11495_));
 sg13g2_nor2_1 _20460_ (.A(net8268),
    .B(_11497_),
    .Y(_11498_));
 sg13g2_xnor2_1 _20461_ (.Y(_11499_),
    .A(_11492_),
    .B(_11497_));
 sg13g2_inv_1 _20462_ (.Y(_11500_),
    .A(_11499_));
 sg13g2_nand2_1 _20463_ (.Y(_11501_),
    .A(_11488_),
    .B(_11499_));
 sg13g2_nor2_1 _20464_ (.A(net8307),
    .B(_11081_),
    .Y(_11502_));
 sg13g2_nor2_1 _20465_ (.A(_11498_),
    .B(_11502_),
    .Y(_11503_));
 sg13g2_a21oi_1 _20466_ (.A1(_11501_),
    .A2(_11503_),
    .Y(_11504_),
    .B1(_11082_));
 sg13g2_a21oi_1 _20467_ (.A1(_11074_),
    .A2(_11504_),
    .Y(_11505_),
    .B1(_11072_));
 sg13g2_xor2_1 _20468_ (.B(_11505_),
    .A(_11047_),
    .X(_11506_));
 sg13g2_xnor2_1 _20469_ (.Y(_11507_),
    .A(_11047_),
    .B(_11505_));
 sg13g2_xnor2_1 _20470_ (.Y(_11508_),
    .A(_11074_),
    .B(_11504_));
 sg13g2_o21ai_1 _20471_ (.B1(_11484_),
    .Y(_11509_),
    .A1(_11434_),
    .A2(_11468_));
 sg13g2_nand3b_1 _20472_ (.B(_11479_),
    .C(_11509_),
    .Y(_11510_),
    .A_N(_11446_));
 sg13g2_and4_1 _20473_ (.A(_11445_),
    .B(_11456_),
    .C(_11457_),
    .D(_11510_),
    .X(_11511_));
 sg13g2_a22oi_1 _20474_ (.Y(_11512_),
    .B1(_11510_),
    .B2(_11445_),
    .A2(_11457_),
    .A1(_11456_));
 sg13g2_or2_1 _20475_ (.X(_11513_),
    .B(_11512_),
    .A(_11511_));
 sg13g2_a21o_1 _20476_ (.A2(_11509_),
    .A1(_11479_),
    .B1(_11446_),
    .X(_11514_));
 sg13g2_nand3_1 _20477_ (.B(_11479_),
    .C(_11509_),
    .A(_11446_),
    .Y(_11515_));
 sg13g2_a21oi_1 _20478_ (.A1(_11262_),
    .A2(_11298_),
    .Y(_11516_),
    .B1(_11315_));
 sg13g2_nor3_1 _20479_ (.A(_11276_),
    .B(_11311_),
    .C(_11516_),
    .Y(_11517_));
 sg13g2_nor2_1 _20480_ (.A(_11275_),
    .B(_11517_),
    .Y(_11518_));
 sg13g2_xnor2_1 _20481_ (.Y(_11519_),
    .A(_11286_),
    .B(_11518_));
 sg13g2_a21oi_1 _20482_ (.A1(_11319_),
    .A2(_11423_),
    .Y(_11520_),
    .B1(_11428_));
 sg13g2_xnor2_1 _20483_ (.Y(_11521_),
    .A(_11357_),
    .B(_11520_));
 sg13g2_a21oi_1 _20484_ (.A1(_11319_),
    .A2(_11386_),
    .Y(_11522_),
    .B1(_11425_));
 sg13g2_nor3_1 _20485_ (.A(_11397_),
    .B(_11420_),
    .C(_11522_),
    .Y(_11523_));
 sg13g2_or3_1 _20486_ (.A(_11397_),
    .B(_11420_),
    .C(_11522_),
    .X(_11524_));
 sg13g2_o21ai_1 _20487_ (.B1(_11397_),
    .Y(_11525_),
    .A1(_11420_),
    .A2(_11522_));
 sg13g2_and2_1 _20488_ (.A(_11524_),
    .B(_11525_),
    .X(_11526_));
 sg13g2_a21oi_1 _20489_ (.A1(_11524_),
    .A2(_11525_),
    .Y(_11527_),
    .B1(_11521_));
 sg13g2_nand4_1 _20490_ (.B(_11515_),
    .C(_11519_),
    .A(_11514_),
    .Y(_11528_),
    .D(_11527_));
 sg13g2_o21ai_1 _20491_ (.B1(_11356_),
    .Y(_11529_),
    .A1(_11358_),
    .A2(_11520_));
 sg13g2_xnor2_1 _20492_ (.Y(_11530_),
    .A(_11372_),
    .B(_11529_));
 sg13g2_o21ai_1 _20493_ (.B1(_11408_),
    .Y(_11531_),
    .A1(_11396_),
    .A2(_11523_));
 sg13g2_or3_1 _20494_ (.A(_11396_),
    .B(_11408_),
    .C(_11523_),
    .X(_11532_));
 sg13g2_nand3_1 _20495_ (.B(_11531_),
    .C(_11532_),
    .A(_11530_),
    .Y(_11533_));
 sg13g2_nor4_1 _20496_ (.A(_11511_),
    .B(_11512_),
    .C(_11528_),
    .D(_11533_),
    .Y(_11534_));
 sg13g2_a21oi_1 _20497_ (.A1(_11368_),
    .A2(_11529_),
    .Y(_11535_),
    .B1(_11370_));
 sg13g2_o21ai_1 _20498_ (.B1(_11330_),
    .Y(_11536_),
    .A1(_11331_),
    .A2(_11535_));
 sg13g2_xor2_1 _20499_ (.B(_11536_),
    .A(_11344_),
    .X(_11537_));
 sg13g2_or2_1 _20500_ (.X(_11538_),
    .B(_11502_),
    .A(_11082_));
 sg13g2_a21oi_1 _20501_ (.A1(_11488_),
    .A2(_11499_),
    .Y(_11539_),
    .B1(_11498_));
 sg13g2_xor2_1 _20502_ (.B(_11539_),
    .A(_11538_),
    .X(_11540_));
 sg13g2_xor2_1 _20503_ (.B(_11535_),
    .A(_11331_),
    .X(_11541_));
 sg13g2_o21ai_1 _20504_ (.B1(_11467_),
    .Y(_11542_),
    .A1(_11434_),
    .A2(_11468_));
 sg13g2_xor2_1 _20505_ (.B(_11542_),
    .A(_11481_),
    .X(_11543_));
 sg13g2_xnor2_1 _20506_ (.Y(_11544_),
    .A(_11488_),
    .B(_11499_));
 sg13g2_o21ai_1 _20507_ (.B1(_11276_),
    .Y(_11545_),
    .A1(_11311_),
    .A2(_11516_));
 sg13g2_nor2b_1 _20508_ (.A(_11517_),
    .B_N(_11545_),
    .Y(_11546_));
 sg13g2_xnor2_1 _20509_ (.Y(_11547_),
    .A(_11319_),
    .B(_11387_));
 sg13g2_a21oi_1 _20510_ (.A1(_11202_),
    .A2(_11215_),
    .Y(_11548_),
    .B1(_11256_));
 sg13g2_a21oi_1 _20511_ (.A1(_11246_),
    .A2(_11251_),
    .Y(_11549_),
    .B1(_11548_));
 sg13g2_a21oi_1 _20512_ (.A1(_11230_),
    .A2(_11549_),
    .Y(_11550_),
    .B1(_11227_));
 sg13g2_xor2_1 _20513_ (.B(_11550_),
    .A(_11241_),
    .X(_11551_));
 sg13g2_o21ai_1 _20514_ (.B1(_11296_),
    .Y(_11552_),
    .A1(_11261_),
    .A2(_11297_));
 sg13g2_xor2_1 _20515_ (.B(_11552_),
    .A(_11313_),
    .X(_11553_));
 sg13g2_xnor2_1 _20516_ (.Y(_11554_),
    .A(_11230_),
    .B(_11549_));
 sg13g2_xnor2_1 _20517_ (.Y(_11555_),
    .A(_11262_),
    .B(_11298_));
 sg13g2_a21oi_1 _20518_ (.A1(_11202_),
    .A2(_11215_),
    .Y(_11556_),
    .B1(_11214_));
 sg13g2_xor2_1 _20519_ (.B(_11556_),
    .A(_11254_),
    .X(_11557_));
 sg13g2_xnor2_1 _20520_ (.Y(_11558_),
    .A(_11202_),
    .B(_11216_));
 sg13g2_nor2b_1 _20521_ (.A(_11092_),
    .B_N(_11199_),
    .Y(_11559_));
 sg13g2_nand2_1 _20522_ (.Y(_11560_),
    .A(_11102_),
    .B(_11200_));
 sg13g2_nand2_1 _20523_ (.Y(_11561_),
    .A(_11198_),
    .B(_11200_));
 sg13g2_xor2_1 _20524_ (.B(_11561_),
    .A(_11559_),
    .X(_11562_));
 sg13g2_xor2_1 _20525_ (.B(_11560_),
    .A(_11197_),
    .X(_11563_));
 sg13g2_or2_1 _20526_ (.X(_11564_),
    .B(_11113_),
    .A(_11112_));
 sg13g2_xor2_1 _20527_ (.B(_11564_),
    .A(_11195_),
    .X(_11565_));
 sg13g2_o21ai_1 _20528_ (.B1(_11128_),
    .Y(_11566_),
    .A1(_11139_),
    .A2(_11193_));
 sg13g2_nand2b_1 _20529_ (.Y(_11567_),
    .B(_11566_),
    .A_N(_11194_));
 sg13g2_xor2_1 _20530_ (.B(_11138_),
    .A(net8301),
    .X(_11568_));
 sg13g2_xnor2_1 _20531_ (.Y(_11569_),
    .A(_11192_),
    .B(_11568_));
 sg13g2_xnor2_1 _20532_ (.Y(_11570_),
    .A(_11189_),
    .B(_11190_));
 sg13g2_nor2_1 _20533_ (.A(net8510),
    .B(net8298),
    .Y(_11571_));
 sg13g2_xnor2_1 _20534_ (.Y(_11572_),
    .A(net8519),
    .B(net8298));
 sg13g2_xor2_1 _20535_ (.B(_11188_),
    .A(_11172_),
    .X(_11573_));
 sg13g2_nor4_1 _20536_ (.A(_11569_),
    .B(_11570_),
    .C(_11572_),
    .D(_11573_),
    .Y(_11574_));
 sg13g2_nand4_1 _20537_ (.B(_11563_),
    .C(_11567_),
    .A(_11562_),
    .Y(_11575_),
    .D(_11574_));
 sg13g2_nor4_1 _20538_ (.A(_11557_),
    .B(_11558_),
    .C(_11565_),
    .D(_11575_),
    .Y(_11576_));
 sg13g2_nand4_1 _20539_ (.B(_11554_),
    .C(_11555_),
    .A(_11553_),
    .Y(_11577_),
    .D(_11576_));
 sg13g2_nor4_2 _20540_ (.A(_11546_),
    .B(_11547_),
    .C(_11551_),
    .Y(_11578_),
    .D(_11577_));
 sg13g2_a21oi_1 _20541_ (.A1(_11319_),
    .A2(_11386_),
    .Y(_11579_),
    .B1(_11385_));
 sg13g2_xor2_1 _20542_ (.B(_11579_),
    .A(_11422_),
    .X(_11580_));
 sg13g2_xnor2_1 _20543_ (.Y(_11581_),
    .A(_11434_),
    .B(_11469_));
 sg13g2_nor2_1 _20544_ (.A(_11580_),
    .B(_11581_),
    .Y(_11582_));
 sg13g2_nand4_1 _20545_ (.B(_11544_),
    .C(_11578_),
    .A(_11543_),
    .Y(_11583_),
    .D(_11582_));
 sg13g2_nor3_1 _20546_ (.A(_11540_),
    .B(_11541_),
    .C(_11583_),
    .Y(_11584_));
 sg13g2_nand4_1 _20547_ (.B(_11534_),
    .C(_11537_),
    .A(_11508_),
    .Y(_11585_),
    .D(_11584_));
 sg13g2_nand2b_1 _20548_ (.Y(_11586_),
    .B(_11507_),
    .A_N(_11585_));
 sg13g2_o21ai_1 _20549_ (.B1(_10967_),
    .Y(_11587_),
    .A1(_11506_),
    .A2(_11585_));
 sg13g2_nor2_1 _20550_ (.A(_10930_),
    .B(_11024_),
    .Y(_11588_));
 sg13g2_nand2_1 _20551_ (.Y(_11589_),
    .A(_10948_),
    .B(_10964_));
 sg13g2_nor2_1 _20552_ (.A(_10930_),
    .B(_11589_),
    .Y(_11590_));
 sg13g2_nor2_1 _20553_ (.A(_10930_),
    .B(_11035_),
    .Y(_11591_));
 sg13g2_nand2_1 _20554_ (.Y(_11592_),
    .A(net8314),
    .B(_11021_));
 sg13g2_nor4_1 _20555_ (.A(_11047_),
    .B(_11073_),
    .C(_11500_),
    .D(_11538_),
    .Y(_11593_));
 sg13g2_nor4_1 _20556_ (.A(_11047_),
    .B(_11073_),
    .C(_11082_),
    .D(_11503_),
    .Y(_11594_));
 sg13g2_or2_1 _20557_ (.X(_11595_),
    .B(_11072_),
    .A(_11046_));
 sg13g2_a221oi_1 _20558_ (.B2(_11045_),
    .C1(_11594_),
    .B1(_11595_),
    .A1(_11488_),
    .Y(_11596_),
    .A2(_11593_));
 sg13g2_nand2_1 _20559_ (.Y(_11597_),
    .A(net8314),
    .B(_11022_));
 sg13g2_nand2_1 _20560_ (.Y(_11598_),
    .A(_10993_),
    .B(_11021_));
 sg13g2_inv_1 _20561_ (.Y(_11599_),
    .A(_11598_));
 sg13g2_and2_1 _20562_ (.A(_11597_),
    .B(_11598_),
    .X(_11600_));
 sg13g2_o21ai_1 _20563_ (.B1(_11592_),
    .Y(_11601_),
    .A1(_11596_),
    .A2(_11600_));
 sg13g2_inv_1 _20564_ (.Y(_11602_),
    .A(_11601_));
 sg13g2_nor2_1 _20565_ (.A(_10966_),
    .B(_11031_),
    .Y(_11603_));
 sg13g2_mux2_1 _20566_ (.A0(_11603_),
    .A1(_11032_),
    .S(_11596_),
    .X(_11604_));
 sg13g2_mux2_1 _20567_ (.A0(_11604_),
    .A1(_11601_),
    .S(_11591_),
    .X(_11605_));
 sg13g2_a21oi_1 _20568_ (.A1(_11590_),
    .A2(_11601_),
    .Y(_11606_),
    .B1(_10967_));
 sg13g2_o21ai_1 _20569_ (.B1(_11606_),
    .Y(_11607_),
    .A1(_11590_),
    .A2(_11605_));
 sg13g2_nor2b_1 _20570_ (.A(_11588_),
    .B_N(_11607_),
    .Y(_11608_));
 sg13g2_and2_1 _20571_ (.A(_10930_),
    .B(_11027_),
    .X(_11609_));
 sg13g2_a221oi_1 _20572_ (.B2(_11587_),
    .C1(_11609_),
    .B1(_11608_),
    .A1(_11586_),
    .Y(_11610_),
    .A2(_11588_));
 sg13g2_nor2_1 _20573_ (.A(_11031_),
    .B(_11035_),
    .Y(_11611_));
 sg13g2_nand2_1 _20574_ (.Y(_11612_),
    .A(_10929_),
    .B(_11028_));
 sg13g2_nor2_1 _20575_ (.A(_10964_),
    .B(_11612_),
    .Y(_11613_));
 sg13g2_inv_1 _20576_ (.Y(_11614_),
    .A(_11613_));
 sg13g2_nand2_1 _20577_ (.Y(_11615_),
    .A(_11596_),
    .B(_11613_));
 sg13g2_nor2_1 _20578_ (.A(net8529),
    .B(_11612_),
    .Y(_11616_));
 sg13g2_inv_1 _20579_ (.Y(_11617_),
    .A(_11616_));
 sg13g2_o21ai_1 _20580_ (.B1(_11615_),
    .Y(_11618_),
    .A1(_11596_),
    .A2(_11617_));
 sg13g2_nor2_1 _20581_ (.A(_11030_),
    .B(_11589_),
    .Y(_11619_));
 sg13g2_nor2_1 _20582_ (.A(_11031_),
    .B(_11589_),
    .Y(_11620_));
 sg13g2_nand2_1 _20583_ (.Y(_11621_),
    .A(_11028_),
    .B(_11619_));
 sg13g2_nor3_1 _20584_ (.A(_10947_),
    .B(_10964_),
    .C(_11031_),
    .Y(_11622_));
 sg13g2_mux2_1 _20585_ (.A0(_11611_),
    .A1(_11620_),
    .S(_11601_),
    .X(_11623_));
 sg13g2_or2_1 _20586_ (.X(_11624_),
    .B(net7677),
    .A(net7679));
 sg13g2_nand2b_1 _20587_ (.Y(_11625_),
    .B(_11620_),
    .A_N(_11601_));
 sg13g2_mux2_1 _20588_ (.A0(_11614_),
    .A1(_11617_),
    .S(_11596_),
    .X(_11626_));
 sg13g2_mux2_1 _20589_ (.A0(_11613_),
    .A1(_11616_),
    .S(_11596_),
    .X(_11627_));
 sg13g2_a21oi_1 _20590_ (.A1(_11601_),
    .A2(_11611_),
    .Y(_11628_),
    .B1(_11627_));
 sg13g2_o21ai_1 _20591_ (.B1(_11626_),
    .Y(_11629_),
    .A1(_11601_),
    .A2(_11621_));
 sg13g2_and2_1 _20592_ (.A(_11601_),
    .B(_11622_),
    .X(_11630_));
 sg13g2_nand2_1 _20593_ (.Y(_11631_),
    .A(_11625_),
    .B(_11628_));
 sg13g2_inv_1 _20594_ (.Y(_11632_),
    .A(net7669));
 sg13g2_nand3_1 _20595_ (.B(_11036_),
    .C(_11596_),
    .A(_11034_),
    .Y(_11633_));
 sg13g2_nor4_1 _20596_ (.A(_10929_),
    .B(_10948_),
    .C(_11028_),
    .D(_11041_),
    .Y(_11634_));
 sg13g2_inv_1 _20597_ (.Y(_11635_),
    .A(net8266));
 sg13g2_nor3_1 _20598_ (.A(_10947_),
    .B(_11028_),
    .C(_11030_),
    .Y(_11636_));
 sg13g2_nand4_1 _20599_ (.B(_11026_),
    .C(_11027_),
    .A(_10948_),
    .Y(_11637_),
    .D(_11029_));
 sg13g2_nor2_2 _20600_ (.A(net8529),
    .B(net8260),
    .Y(_11638_));
 sg13g2_nand2_1 _20601_ (.Y(_11639_),
    .A(_10964_),
    .B(net8263));
 sg13g2_nand2_1 _20602_ (.Y(_11640_),
    .A(net8004),
    .B(net8003));
 sg13g2_nand2_2 _20603_ (.Y(_11641_),
    .A(net8529),
    .B(net8263));
 sg13g2_o21ai_1 _20604_ (.B1(_11182_),
    .Y(_11642_),
    .A1(net8298),
    .A2(_11641_));
 sg13g2_a21oi_1 _20605_ (.A1(net8529),
    .A2(net8263),
    .Y(_11643_),
    .B1(_10880_));
 sg13g2_nand4_1 _20606_ (.B(_10929_),
    .C(_11026_),
    .A(_10890_),
    .Y(_11644_),
    .D(_11027_));
 sg13g2_nor2_2 _20607_ (.A(_11024_),
    .B(_11644_),
    .Y(_11645_));
 sg13g2_or2_1 _20608_ (.X(_11646_),
    .B(_11644_),
    .A(_11024_));
 sg13g2_o21ai_1 _20609_ (.B1(net7999),
    .Y(_11647_),
    .A1(net8298),
    .A2(net8256));
 sg13g2_a22oi_1 _20610_ (.Y(_11648_),
    .B1(_11642_),
    .B2(_11647_),
    .A2(_11640_),
    .A1(_11572_));
 sg13g2_a21oi_2 _20611_ (.B1(net8519),
    .Y(_11649_),
    .A2(_11166_),
    .A1(_11165_));
 sg13g2_a21o_2 _20612_ (.A2(_11166_),
    .A1(_11165_),
    .B1(net8519),
    .X(_11650_));
 sg13g2_nor2_2 _20613_ (.A(net8425),
    .B(_11650_),
    .Y(_11651_));
 sg13g2_nand2_1 _20614_ (.Y(_11652_),
    .A(net8390),
    .B(_11571_));
 sg13g2_nor2_2 _20615_ (.A(net8410),
    .B(_11652_),
    .Y(_11653_));
 sg13g2_nor2_2 _20616_ (.A(_10966_),
    .B(_11644_),
    .Y(_11654_));
 sg13g2_or2_2 _20617_ (.X(_11655_),
    .B(_11644_),
    .A(_10966_));
 sg13g2_nor2_2 _20618_ (.A(net8439),
    .B(_11655_),
    .Y(_11656_));
 sg13g2_nand2_1 _20619_ (.Y(_11657_),
    .A(net8432),
    .B(_11654_));
 sg13g2_nand2_1 _20620_ (.Y(_11658_),
    .A(_11653_),
    .B(_11656_));
 sg13g2_nand3_1 _20621_ (.B(_11653_),
    .C(_11656_),
    .A(net8444),
    .Y(_11659_));
 sg13g2_nor2_2 _20622_ (.A(net8450),
    .B(_11655_),
    .Y(_11660_));
 sg13g2_nand2_1 _20623_ (.Y(_11661_),
    .A(net8445),
    .B(_11654_));
 sg13g2_nor2_1 _20624_ (.A(net8387),
    .B(net8277),
    .Y(_11662_));
 sg13g2_a21oi_1 _20625_ (.A1(net8387),
    .A2(net8283),
    .Y(_11663_),
    .B1(_11662_));
 sg13g2_nand2_1 _20626_ (.Y(_11664_),
    .A(net8387),
    .B(net8282));
 sg13g2_o21ai_1 _20627_ (.B1(_11664_),
    .Y(_11665_),
    .A1(net8387),
    .A2(net8280));
 sg13g2_nor2_1 _20628_ (.A(net8396),
    .B(_11665_),
    .Y(_11666_));
 sg13g2_a21oi_2 _20629_ (.B1(_11666_),
    .Y(_11667_),
    .A2(_11663_),
    .A1(net8397));
 sg13g2_nand2_1 _20630_ (.Y(_11668_),
    .A(net8386),
    .B(_11349_));
 sg13g2_nor2_1 _20631_ (.A(net8386),
    .B(net8285),
    .Y(_11669_));
 sg13g2_a21oi_1 _20632_ (.A1(net8386),
    .A2(_11349_),
    .Y(_11670_),
    .B1(_11669_));
 sg13g2_nor2_1 _20633_ (.A(net8386),
    .B(_11335_),
    .Y(_11671_));
 sg13g2_a21oi_2 _20634_ (.B1(_11671_),
    .Y(_11672_),
    .A2(net8289),
    .A1(net8386));
 sg13g2_mux2_1 _20635_ (.A0(_11670_),
    .A1(_11672_),
    .S(net8407),
    .X(_11673_));
 sg13g2_nor2_1 _20636_ (.A(net8422),
    .B(_11667_),
    .Y(_11674_));
 sg13g2_a21oi_2 _20637_ (.B1(_11674_),
    .Y(_11675_),
    .A2(_11673_),
    .A1(net8422));
 sg13g2_nand2_1 _20638_ (.Y(_11676_),
    .A(net8514),
    .B(net8270));
 sg13g2_o21ai_1 _20639_ (.B1(_11676_),
    .Y(_11677_),
    .A1(net8514),
    .A2(_11463_));
 sg13g2_nor2_1 _20640_ (.A(net8385),
    .B(net8274),
    .Y(_11678_));
 sg13g2_a21oi_1 _20641_ (.A1(net8385),
    .A2(net8275),
    .Y(_11679_),
    .B1(_11678_));
 sg13g2_nand2_1 _20642_ (.Y(_11680_),
    .A(net8404),
    .B(_11679_));
 sg13g2_o21ai_1 _20643_ (.B1(_11680_),
    .Y(_11681_),
    .A1(net8404),
    .A2(_11677_));
 sg13g2_nand2_1 _20644_ (.Y(_11682_),
    .A(net8308),
    .B(net8514));
 sg13g2_o21ai_1 _20645_ (.B1(_11682_),
    .Y(_11683_),
    .A1(net8514),
    .A2(_11492_));
 sg13g2_nand2_1 _20646_ (.Y(_11684_),
    .A(_11052_),
    .B(net8384));
 sg13g2_o21ai_1 _20647_ (.B1(_11684_),
    .Y(_11685_),
    .A1(_10993_),
    .A2(net8384));
 sg13g2_mux2_1 _20648_ (.A0(_11683_),
    .A1(_11685_),
    .S(net8408),
    .X(_11686_));
 sg13g2_nand2_1 _20649_ (.Y(_11687_),
    .A(net8417),
    .B(_11686_));
 sg13g2_o21ai_1 _20650_ (.B1(_11687_),
    .Y(_11688_),
    .A1(net8419),
    .A2(_11681_));
 sg13g2_mux2_1 _20651_ (.A0(_11675_),
    .A1(_11688_),
    .S(net8439),
    .X(_11689_));
 sg13g2_nor2_1 _20652_ (.A(_11143_),
    .B(net8509),
    .Y(_11690_));
 sg13g2_nand2_1 _20653_ (.Y(_11691_),
    .A(net8302),
    .B(net8509));
 sg13g2_nor2b_1 _20654_ (.A(_11690_),
    .B_N(_11691_),
    .Y(_11692_));
 sg13g2_nand2_1 _20655_ (.Y(_11693_),
    .A(net8300),
    .B(net8509));
 sg13g2_nand2_1 _20656_ (.Y(_11694_),
    .A(net8305),
    .B(net8511));
 sg13g2_o21ai_1 _20657_ (.B1(_11694_),
    .Y(_11695_),
    .A1(net8303),
    .A2(net8511));
 sg13g2_nand2_1 _20658_ (.Y(_11696_),
    .A(_11087_),
    .B(net8511));
 sg13g2_o21ai_1 _20659_ (.B1(_11696_),
    .Y(_11697_),
    .A1(_11096_),
    .A2(net8511));
 sg13g2_nor2_1 _20660_ (.A(net8391),
    .B(_11697_),
    .Y(_11698_));
 sg13g2_a21oi_1 _20661_ (.A1(net8391),
    .A2(_11695_),
    .Y(_11699_),
    .B1(_11698_));
 sg13g2_nor2_1 _20662_ (.A(net8451),
    .B(net8441),
    .Y(_11700_));
 sg13g2_nand2_2 _20663_ (.Y(_11701_),
    .A(net8446),
    .B(net8431));
 sg13g2_nor2_1 _20664_ (.A(net8400),
    .B(_11571_),
    .Y(_11702_));
 sg13g2_a221oi_1 _20665_ (.B2(_11702_),
    .C1(net8409),
    .B1(_11693_),
    .A1(net8401),
    .Y(_11703_),
    .A2(_11692_));
 sg13g2_o21ai_1 _20666_ (.B1(net8253),
    .Y(_11704_),
    .A1(net8427),
    .A2(_11699_));
 sg13g2_nor2_2 _20667_ (.A(_10947_),
    .B(_11644_),
    .Y(_11705_));
 sg13g2_nand2b_2 _20668_ (.Y(_11706_),
    .B(_10948_),
    .A_N(_11644_));
 sg13g2_nor2_1 _20669_ (.A(net8451),
    .B(net8436),
    .Y(_11707_));
 sg13g2_nand2_2 _20670_ (.Y(_11708_),
    .A(net8444),
    .B(net8439));
 sg13g2_nand2_1 _20671_ (.Y(_11709_),
    .A(net8388),
    .B(_11207_));
 sg13g2_nand2_1 _20672_ (.Y(_11710_),
    .A(net8511),
    .B(_11246_));
 sg13g2_and3_1 _20673_ (.X(_11711_),
    .A(net8391),
    .B(_11709_),
    .C(_11710_));
 sg13g2_nor2_1 _20674_ (.A(net8383),
    .B(net8297),
    .Y(_11712_));
 sg13g2_a21oi_1 _20675_ (.A1(net8388),
    .A2(_11221_),
    .Y(_11713_),
    .B1(_11712_));
 sg13g2_a21oi_1 _20676_ (.A1(net8403),
    .A2(_11713_),
    .Y(_11714_),
    .B1(_11711_));
 sg13g2_nand2_1 _20677_ (.Y(_11715_),
    .A(net8513),
    .B(_11303_));
 sg13g2_o21ai_1 _20678_ (.B1(_11715_),
    .Y(_11716_),
    .A1(net8513),
    .A2(_11291_));
 sg13g2_nor2_1 _20679_ (.A(net8387),
    .B(net8294),
    .Y(_11717_));
 sg13g2_a21oi_1 _20680_ (.A1(net8387),
    .A2(net8295),
    .Y(_11718_),
    .B1(_11717_));
 sg13g2_nand2_1 _20681_ (.Y(_11719_),
    .A(net8406),
    .B(_11718_));
 sg13g2_o21ai_1 _20682_ (.B1(_11719_),
    .Y(_11720_),
    .A1(net8403),
    .A2(_11716_));
 sg13g2_nor2_1 _20683_ (.A(net8420),
    .B(_11714_),
    .Y(_11721_));
 sg13g2_a21oi_2 _20684_ (.B1(_11721_),
    .Y(_11722_),
    .A2(_11720_),
    .A1(net8420));
 sg13g2_o21ai_1 _20685_ (.B1(_11705_),
    .Y(_11723_),
    .A1(_11703_),
    .A2(_11704_));
 sg13g2_a221oi_1 _20686_ (.B2(_11722_),
    .C1(_11723_),
    .B1(net8247),
    .A1(net8447),
    .Y(_11724_),
    .A2(_11689_));
 sg13g2_inv_1 _20687_ (.Y(_11725_),
    .A(_11724_));
 sg13g2_nand4_1 _20688_ (.B(_11648_),
    .C(_11659_),
    .A(_11633_),
    .Y(_11726_),
    .D(_11725_));
 sg13g2_a221oi_1 _20689_ (.B2(net8519),
    .C1(_11726_),
    .B1(net7673),
    .A1(_11037_),
    .Y(_11727_),
    .A2(_11602_));
 sg13g2_o21ai_1 _20690_ (.B1(_11727_),
    .Y(_11728_),
    .A1(net8298),
    .A2(_11632_));
 sg13g2_nor2_2 _20691_ (.A(_11610_),
    .B(_11728_),
    .Y(_11729_));
 sg13g2_o21ai_1 _20692_ (.B1(_10869_),
    .Y(_11730_),
    .A1(_11610_),
    .A2(_11728_));
 sg13g2_nand2_2 _20693_ (.Y(_11731_),
    .A(_10832_),
    .B(net8975));
 sg13g2_nor2_1 _20694_ (.A(net9203),
    .B(_11731_),
    .Y(_11732_));
 sg13g2_nor2_2 _20695_ (.A(_10984_),
    .B(_11732_),
    .Y(_11733_));
 sg13g2_o21ai_1 _20696_ (.B1(_10985_),
    .Y(_11734_),
    .A1(net9204),
    .A2(_11731_));
 sg13g2_nor2_1 _20697_ (.A(net8977),
    .B(_10979_),
    .Y(_11735_));
 sg13g2_nand3_1 _20698_ (.B(_10838_),
    .C(net8974),
    .A(net8980),
    .Y(_11736_));
 sg13g2_nand2_1 _20699_ (.Y(_11737_),
    .A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[0] ),
    .B(net8836));
 sg13g2_or2_1 _20700_ (.X(_11738_),
    .B(_10847_),
    .A(_10841_));
 sg13g2_nor2_1 _20701_ (.A(_10836_),
    .B(_11738_),
    .Y(_11739_));
 sg13g2_or2_1 _20702_ (.X(_11740_),
    .B(_11738_),
    .A(_10836_));
 sg13g2_a21oi_1 _20703_ (.A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[0] ),
    .A2(net8701),
    .Y(_11741_),
    .B1(net8696));
 sg13g2_o21ai_1 _20704_ (.B1(net8662),
    .Y(_11742_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[0] ),
    .A2(net8690));
 sg13g2_a21oi_1 _20705_ (.A1(_11737_),
    .A2(_11741_),
    .Y(_11743_),
    .B1(_11742_));
 sg13g2_nor2_1 _20706_ (.A(net8708),
    .B(_11743_),
    .Y(_11744_));
 sg13g2_nand3_1 _20707_ (.B(net8634),
    .C(_11740_),
    .A(net8664),
    .Y(_11745_));
 sg13g2_nor4_2 _20708_ (.A(net8743),
    .B(_10851_),
    .C(net8702),
    .Y(_11746_),
    .D(_11745_));
 sg13g2_a21oi_1 _20709_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[0] ),
    .A2(net8730),
    .Y(_11747_),
    .B1(net8627));
 sg13g2_nor2_1 _20710_ (.A(net8500),
    .B(_11747_),
    .Y(_11748_));
 sg13g2_inv_1 _20711_ (.Y(_11749_),
    .A(_11748_));
 sg13g2_a21o_1 _20712_ (.A2(_11744_),
    .A1(_11730_),
    .B1(_11749_),
    .X(_11750_));
 sg13g2_nand3_1 _20713_ (.B(_10832_),
    .C(_10838_),
    .A(net9198),
    .Y(_11751_));
 sg13g2_nand2_1 _20714_ (.Y(_11752_),
    .A(\soc_I.kianv_I.datapath_unit_I.ALUOut[0] ),
    .B(_11751_));
 sg13g2_nand3_1 _20715_ (.B(net9197),
    .C(_10832_),
    .A(net9196),
    .Y(_11753_));
 sg13g2_o21ai_1 _20716_ (.B1(_11752_),
    .Y(_11754_),
    .A1(net8977),
    .A2(_11753_));
 sg13g2_nand2_1 _20717_ (.Y(_11755_),
    .A(net8504),
    .B(_11754_));
 sg13g2_and2_1 _20718_ (.A(_11750_),
    .B(_11755_),
    .X(_11756_));
 sg13g2_and2_2 _20719_ (.A(\soc_I.PC[0] ),
    .B(_10858_),
    .X(_11757_));
 sg13g2_a21oi_2 _20720_ (.B1(_10858_),
    .Y(_11758_),
    .A2(_11755_),
    .A1(_11750_));
 sg13g2_or2_2 _20721_ (.X(\soc_I.clint_I.addr[0] ),
    .B(_11758_),
    .A(_11757_));
 sg13g2_nor2_2 _20722_ (.A(\soc_I.PC[1] ),
    .B(net8576),
    .Y(_11759_));
 sg13g2_and2_2 _20723_ (.A(net8504),
    .B(_11751_),
    .X(_11760_));
 sg13g2_o21ai_1 _20724_ (.B1(net7997),
    .Y(_11761_),
    .A1(net8299),
    .A2(net8001));
 sg13g2_nor2_1 _20725_ (.A(net8517),
    .B(net8277),
    .Y(_11762_));
 sg13g2_nand2_1 _20726_ (.Y(_11763_),
    .A(net8515),
    .B(net8282));
 sg13g2_nor2b_1 _20727_ (.A(_11762_),
    .B_N(_11763_),
    .Y(_11764_));
 sg13g2_nand2_1 _20728_ (.Y(_11765_),
    .A(net8516),
    .B(net8286));
 sg13g2_o21ai_1 _20729_ (.B1(_11765_),
    .Y(_11766_),
    .A1(net8515),
    .A2(net8280));
 sg13g2_nor2_1 _20730_ (.A(net8395),
    .B(_11766_),
    .Y(_11767_));
 sg13g2_a21oi_2 _20731_ (.B1(_11767_),
    .Y(_11768_),
    .A2(_11764_),
    .A1(net8397));
 sg13g2_nor2_1 _20732_ (.A(net8515),
    .B(net8285),
    .Y(_11769_));
 sg13g2_a21oi_1 _20733_ (.A1(net8515),
    .A2(net8289),
    .Y(_11770_),
    .B1(_11769_));
 sg13g2_nand2_1 _20734_ (.Y(_11771_),
    .A(net8395),
    .B(_11770_));
 sg13g2_nor2_1 _20735_ (.A(net8515),
    .B(_11335_),
    .Y(_11772_));
 sg13g2_nand2_1 _20736_ (.Y(_11773_),
    .A(net8515),
    .B(net8271));
 sg13g2_nand2b_1 _20737_ (.Y(_11774_),
    .B(_11773_),
    .A_N(_11772_));
 sg13g2_o21ai_1 _20738_ (.B1(_11771_),
    .Y(_11775_),
    .A1(net8395),
    .A2(_11774_));
 sg13g2_nand2_1 _20739_ (.Y(_11776_),
    .A(net8415),
    .B(_11775_));
 sg13g2_o21ai_1 _20740_ (.B1(_11776_),
    .Y(_11777_),
    .A1(net8415),
    .A2(_11768_));
 sg13g2_nand2_1 _20741_ (.Y(_11778_),
    .A(net8434),
    .B(_11777_));
 sg13g2_nand2_1 _20742_ (.Y(_11779_),
    .A(net8384),
    .B(_11472_));
 sg13g2_o21ai_1 _20743_ (.B1(_11779_),
    .Y(_11780_),
    .A1(net8384),
    .A2(_11440_));
 sg13g2_nor2_1 _20744_ (.A(net8514),
    .B(net8274),
    .Y(_11781_));
 sg13g2_a21oi_1 _20745_ (.A1(net8514),
    .A2(net8269),
    .Y(_11782_),
    .B1(_11781_));
 sg13g2_nand2_1 _20746_ (.Y(_11783_),
    .A(net8404),
    .B(_11782_));
 sg13g2_o21ai_1 _20747_ (.B1(_11783_),
    .Y(_11784_),
    .A1(net8404),
    .A2(_11780_));
 sg13g2_nand2_1 _20748_ (.Y(_11785_),
    .A(net8308),
    .B(net8384));
 sg13g2_o21ai_1 _20749_ (.B1(_11785_),
    .Y(_11786_),
    .A1(_11053_),
    .A2(net8384));
 sg13g2_nand2_1 _20750_ (.Y(_11787_),
    .A(net8393),
    .B(_11786_));
 sg13g2_a21oi_2 _20751_ (.B1(net8315),
    .Y(_11788_),
    .A2(_11705_),
    .A1(_10964_));
 sg13g2_o21ai_1 _20752_ (.B1(_10993_),
    .Y(_11789_),
    .A1(_10965_),
    .A2(net8249));
 sg13g2_o21ai_1 _20753_ (.B1(_11789_),
    .Y(_11790_),
    .A1(net8314),
    .A2(net8514));
 sg13g2_o21ai_1 _20754_ (.B1(_11787_),
    .Y(_11791_),
    .A1(net8393),
    .A2(_11790_));
 sg13g2_nand2_1 _20755_ (.Y(_11792_),
    .A(net8416),
    .B(_11791_));
 sg13g2_o21ai_1 _20756_ (.B1(_11792_),
    .Y(_11793_),
    .A1(net8416),
    .A2(_11784_));
 sg13g2_o21ai_1 _20757_ (.B1(_11778_),
    .Y(_11794_),
    .A1(net8432),
    .A2(_11793_));
 sg13g2_nor2_1 _20758_ (.A(net8302),
    .B(net8508),
    .Y(_11795_));
 sg13g2_nand2_1 _20759_ (.Y(_11796_),
    .A(net8303),
    .B(net8508));
 sg13g2_nand2b_1 _20760_ (.Y(_11797_),
    .B(_11796_),
    .A_N(_11795_));
 sg13g2_nor2_1 _20761_ (.A(net8299),
    .B(net8511),
    .Y(_11798_));
 sg13g2_a21oi_1 _20762_ (.A1(_11143_),
    .A2(net8511),
    .Y(_11799_),
    .B1(_11798_));
 sg13g2_a21oi_1 _20763_ (.A1(net8401),
    .A2(_11797_),
    .Y(_11800_),
    .B1(net8411));
 sg13g2_o21ai_1 _20764_ (.B1(_11800_),
    .Y(_11801_),
    .A1(net8401),
    .A2(_11799_));
 sg13g2_nand2_1 _20765_ (.Y(_11802_),
    .A(_11097_),
    .B(net8508));
 sg13g2_o21ai_1 _20766_ (.B1(_11802_),
    .Y(_11803_),
    .A1(net8304),
    .A2(net8508));
 sg13g2_nor2_1 _20767_ (.A(_11086_),
    .B(net8508),
    .Y(_11804_));
 sg13g2_a21oi_1 _20768_ (.A1(net8511),
    .A2(_11207_),
    .Y(_11805_),
    .B1(_11804_));
 sg13g2_nand2_1 _20769_ (.Y(_11806_),
    .A(net8402),
    .B(_11805_));
 sg13g2_o21ai_1 _20770_ (.B1(_11806_),
    .Y(_11807_),
    .A1(net8401),
    .A2(_11803_));
 sg13g2_a21oi_1 _20771_ (.A1(net8412),
    .A2(_11807_),
    .Y(_11808_),
    .B1(net8251));
 sg13g2_nand2_1 _20772_ (.Y(_11809_),
    .A(net8383),
    .B(_11246_));
 sg13g2_o21ai_1 _20773_ (.B1(_11809_),
    .Y(_11810_),
    .A1(net8383),
    .A2(_11222_));
 sg13g2_nor2_1 _20774_ (.A(net8512),
    .B(net8297),
    .Y(_11811_));
 sg13g2_a21oi_1 _20775_ (.A1(net8513),
    .A2(_11292_),
    .Y(_11812_),
    .B1(_11811_));
 sg13g2_nand2_1 _20776_ (.Y(_11813_),
    .A(net8402),
    .B(_11812_));
 sg13g2_o21ai_1 _20777_ (.B1(_11813_),
    .Y(_11814_),
    .A1(net8402),
    .A2(_11810_));
 sg13g2_or2_1 _20778_ (.X(_11815_),
    .B(_11814_),
    .A(net8411));
 sg13g2_nand2_1 _20779_ (.Y(_11816_),
    .A(net8383),
    .B(net8291));
 sg13g2_nand2_1 _20780_ (.Y(_11817_),
    .A(net8513),
    .B(net8295));
 sg13g2_nand2_1 _20781_ (.Y(_11818_),
    .A(_11816_),
    .B(_11817_));
 sg13g2_nor2_1 _20782_ (.A(net8517),
    .B(net8294),
    .Y(_11819_));
 sg13g2_a21oi_1 _20783_ (.A1(net8517),
    .A2(net8283),
    .Y(_11820_),
    .B1(_11819_));
 sg13g2_nand2_1 _20784_ (.Y(_11821_),
    .A(net8406),
    .B(_11820_));
 sg13g2_o21ai_1 _20785_ (.B1(_11821_),
    .Y(_11822_),
    .A1(net8402),
    .A2(_11818_));
 sg13g2_o21ai_1 _20786_ (.B1(_11815_),
    .Y(_11823_),
    .A1(net8427),
    .A2(_11822_));
 sg13g2_inv_1 _20787_ (.Y(_11824_),
    .A(_11823_));
 sg13g2_a221oi_1 _20788_ (.B2(net8245),
    .C1(net8250),
    .B1(_11823_),
    .A1(_11801_),
    .Y(_11825_),
    .A2(_11808_));
 sg13g2_o21ai_1 _20789_ (.B1(_11825_),
    .Y(_11826_),
    .A1(net8446),
    .A2(_11794_));
 sg13g2_o21ai_1 _20790_ (.B1(_11187_),
    .Y(_11827_),
    .A1(net8299),
    .A2(net8510));
 sg13g2_nand2b_1 _20791_ (.Y(_11828_),
    .B(net8390),
    .A_N(_11827_));
 sg13g2_nor2_1 _20792_ (.A(net8414),
    .B(_11828_),
    .Y(_11829_));
 sg13g2_nand2_2 _20793_ (.Y(_11830_),
    .A(_11656_),
    .B(_11829_));
 sg13g2_nor2_1 _20794_ (.A(net8400),
    .B(net8262),
    .Y(_11831_));
 sg13g2_a21oi_1 _20795_ (.A1(net8400),
    .A2(net8256),
    .Y(_11832_),
    .B1(_11831_));
 sg13g2_nand2_1 _20796_ (.Y(_11833_),
    .A(net8400),
    .B(_11761_));
 sg13g2_o21ai_1 _20797_ (.B1(_11833_),
    .Y(_11834_),
    .A1(net8449),
    .A2(_11830_));
 sg13g2_a221oi_1 _20798_ (.B2(net8299),
    .C1(_11834_),
    .B1(_11832_),
    .A1(_11573_),
    .Y(_11835_),
    .A2(net8265));
 sg13g2_nand2_1 _20799_ (.Y(_11836_),
    .A(_11826_),
    .B(_11835_));
 sg13g2_a221oi_1 _20800_ (.B2(net8300),
    .C1(_11836_),
    .B1(net7669),
    .A1(net8400),
    .Y(_11837_),
    .A2(net7672));
 sg13g2_o21ai_1 _20801_ (.B1(net8659),
    .Y(_11838_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[1] ),
    .A2(net8691));
 sg13g2_nand2_2 _20802_ (.Y(_11839_),
    .A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[1] ),
    .B(net8839));
 sg13g2_a21oi_2 _20803_ (.B1(net8697),
    .Y(_11840_),
    .A2(net8702),
    .A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[1] ));
 sg13g2_a21oi_1 _20804_ (.A1(_11839_),
    .A2(_11840_),
    .Y(_11841_),
    .B1(_11838_));
 sg13g2_nor2_1 _20805_ (.A(net8706),
    .B(_11841_),
    .Y(_11842_));
 sg13g2_o21ai_1 _20806_ (.B1(_11842_),
    .Y(_11843_),
    .A1(net8659),
    .A2(_11837_));
 sg13g2_a21oi_1 _20807_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[1] ),
    .A2(net8735),
    .Y(_11844_),
    .B1(net8634));
 sg13g2_nor2_1 _20808_ (.A(net8503),
    .B(_11844_),
    .Y(_11845_));
 sg13g2_a22oi_1 _20809_ (.Y(_11846_),
    .B1(_11843_),
    .B2(_11845_),
    .A2(net8377),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[1] ));
 sg13g2_a21oi_2 _20810_ (.B1(_11759_),
    .Y(\soc_I.clint_I.addr[1] ),
    .A2(net7668),
    .A1(net8577));
 sg13g2_nor2_2 _20811_ (.A(\soc_I.qqspi_I.xfer_cycles[1] ),
    .B(\soc_I.qqspi_I.xfer_cycles[0] ),
    .Y(_11847_));
 sg13g2_nor3_1 _20812_ (.A(\soc_I.qqspi_I.xfer_cycles[4] ),
    .B(\soc_I.qqspi_I.xfer_cycles[3] ),
    .C(\soc_I.qqspi_I.xfer_cycles[2] ),
    .Y(_11848_));
 sg13g2_nand2_1 _20813_ (.Y(_11849_),
    .A(_11847_),
    .B(_11848_));
 sg13g2_nor2_1 _20814_ (.A(\soc_I.qqspi_I.xfer_cycles[5] ),
    .B(_11849_),
    .Y(_11850_));
 sg13g2_or2_1 _20815_ (.X(_11851_),
    .B(_11849_),
    .A(\soc_I.qqspi_I.xfer_cycles[5] ));
 sg13g2_o21ai_1 _20816_ (.B1(net7996),
    .Y(_11852_),
    .A1(_11096_),
    .A2(net8000));
 sg13g2_a21oi_1 _20817_ (.A1(net8521),
    .A2(net8255),
    .Y(_11853_),
    .B1(_11097_));
 sg13g2_nand2b_1 _20818_ (.Y(_11854_),
    .B(net8261),
    .A_N(net8521));
 sg13g2_a21o_1 _20819_ (.A2(_11852_),
    .A1(net8521),
    .B1(_11853_),
    .X(_11855_));
 sg13g2_o21ai_1 _20820_ (.B1(_11694_),
    .Y(_11856_),
    .A1(_11097_),
    .A2(net8508));
 sg13g2_o21ai_1 _20821_ (.B1(_11691_),
    .Y(_11857_),
    .A1(net8303),
    .A2(net8508));
 sg13g2_mux2_1 _20822_ (.A0(_11856_),
    .A1(_11857_),
    .S(net8401),
    .X(_11858_));
 sg13g2_nor2_1 _20823_ (.A(net8411),
    .B(_11858_),
    .Y(_11859_));
 sg13g2_nor2b_1 _20824_ (.A(_11690_),
    .B_N(_11693_),
    .Y(_11860_));
 sg13g2_nand2_1 _20825_ (.Y(_11861_),
    .A(net8389),
    .B(_11860_));
 sg13g2_o21ai_1 _20826_ (.B1(_11861_),
    .Y(_11862_),
    .A1(net8390),
    .A2(_11571_));
 sg13g2_a21oi_2 _20827_ (.B1(_11859_),
    .Y(_11863_),
    .A2(_11862_),
    .A1(net8409));
 sg13g2_nor2_2 _20828_ (.A(net8439),
    .B(net7994),
    .Y(_11864_));
 sg13g2_inv_1 _20829_ (.Y(_11865_),
    .A(_11864_));
 sg13g2_nor2_1 _20830_ (.A(net8395),
    .B(_11677_),
    .Y(_11866_));
 sg13g2_a21oi_2 _20831_ (.B1(_11866_),
    .Y(_11867_),
    .A2(_11672_),
    .A1(net8396));
 sg13g2_nand2_1 _20832_ (.Y(_11868_),
    .A(net8394),
    .B(_11679_));
 sg13g2_o21ai_1 _20833_ (.B1(_11868_),
    .Y(_11869_),
    .A1(net8394),
    .A2(_11683_));
 sg13g2_nand2_1 _20834_ (.Y(_11870_),
    .A(net8417),
    .B(_11869_));
 sg13g2_o21ai_1 _20835_ (.B1(_11870_),
    .Y(_11871_),
    .A1(net8416),
    .A2(_11867_));
 sg13g2_nand2_1 _20836_ (.Y(_11872_),
    .A(net8434),
    .B(_11871_));
 sg13g2_nor2_1 _20837_ (.A(net8428),
    .B(_11788_),
    .Y(_11873_));
 sg13g2_nand2_1 _20838_ (.Y(_11874_),
    .A(net8393),
    .B(_11685_));
 sg13g2_o21ai_1 _20839_ (.B1(_11874_),
    .Y(_11875_),
    .A1(net8393),
    .A2(_11788_));
 sg13g2_a21o_1 _20840_ (.A2(_11875_),
    .A1(net8428),
    .B1(_11873_),
    .X(_11876_));
 sg13g2_o21ai_1 _20841_ (.B1(_11872_),
    .Y(_11877_),
    .A1(net8435),
    .A2(_11876_));
 sg13g2_mux2_1 _20842_ (.A0(_11663_),
    .A1(_11718_),
    .S(net8397),
    .X(_11878_));
 sg13g2_nor2_1 _20843_ (.A(net8422),
    .B(_11878_),
    .Y(_11879_));
 sg13g2_nor2_1 _20844_ (.A(net8406),
    .B(_11665_),
    .Y(_11880_));
 sg13g2_a21oi_2 _20845_ (.B1(_11880_),
    .Y(_11881_),
    .A2(_11670_),
    .A1(net8407));
 sg13g2_a21oi_2 _20846_ (.B1(_11879_),
    .Y(_11882_),
    .A2(_11881_),
    .A1(net8422));
 sg13g2_nand3_1 _20847_ (.B(_11709_),
    .C(_11710_),
    .A(net8403),
    .Y(_11883_));
 sg13g2_o21ai_1 _20848_ (.B1(_11883_),
    .Y(_11884_),
    .A1(net8403),
    .A2(_11697_));
 sg13g2_nor2_1 _20849_ (.A(net8392),
    .B(_11716_),
    .Y(_11885_));
 sg13g2_a21oi_2 _20850_ (.B1(_11885_),
    .Y(_11886_),
    .A2(_11713_),
    .A1(net8392));
 sg13g2_o21ai_1 _20851_ (.B1(net8253),
    .Y(_11887_),
    .A1(net8421),
    .A2(_11884_));
 sg13g2_a21oi_1 _20852_ (.A1(net8420),
    .A2(_11886_),
    .Y(_11888_),
    .B1(_11887_));
 sg13g2_a221oi_1 _20853_ (.B2(net8245),
    .C1(_11888_),
    .B1(_11882_),
    .A1(_11124_),
    .Y(_11889_),
    .A2(_11877_));
 sg13g2_nor2_1 _20854_ (.A(net8249),
    .B(_11889_),
    .Y(_11890_));
 sg13g2_a221oi_1 _20855_ (.B2(_11864_),
    .C1(_11890_),
    .B1(_11863_),
    .A1(_11854_),
    .Y(_11891_),
    .A2(_11855_));
 sg13g2_o21ai_1 _20856_ (.B1(_11891_),
    .Y(_11892_),
    .A1(_11563_),
    .A2(net8004));
 sg13g2_a221oi_1 _20857_ (.B2(_11096_),
    .C1(_11892_),
    .B1(net7669),
    .A1(net8521),
    .Y(_11893_),
    .A2(net7672));
 sg13g2_o21ai_1 _20858_ (.B1(_11208_),
    .Y(_11894_),
    .A1(net7676),
    .A2(net7675));
 sg13g2_nor2_1 _20859_ (.A(net8433),
    .B(_11788_),
    .Y(_11895_));
 sg13g2_a21oi_1 _20860_ (.A1(net8435),
    .A2(_11688_),
    .Y(_11896_),
    .B1(net7938));
 sg13g2_mux4_1 _20861_ (.S0(net8432),
    .A0(_11675_),
    .A1(_11722_),
    .A2(_11789_),
    .A3(_11688_),
    .S1(net8448),
    .X(_11897_));
 sg13g2_nor2_1 _20862_ (.A(net8431),
    .B(_11653_),
    .Y(_11898_));
 sg13g2_nand2_1 _20863_ (.Y(_11899_),
    .A(net8389),
    .B(_11857_));
 sg13g2_o21ai_1 _20864_ (.B1(_11899_),
    .Y(_11900_),
    .A1(net8389),
    .A2(_11860_));
 sg13g2_and2_1 _20865_ (.A(net8411),
    .B(_11900_),
    .X(_11901_));
 sg13g2_nand2_1 _20866_ (.Y(_11902_),
    .A(_11696_),
    .B(_11709_));
 sg13g2_nand2_1 _20867_ (.Y(_11903_),
    .A(net8402),
    .B(_11856_));
 sg13g2_o21ai_1 _20868_ (.B1(_11903_),
    .Y(_11904_),
    .A1(net8402),
    .A2(_11902_));
 sg13g2_a21oi_2 _20869_ (.B1(_11901_),
    .Y(_11905_),
    .A2(_11904_),
    .A1(net8429));
 sg13g2_a21oi_2 _20870_ (.B1(_11898_),
    .Y(_11906_),
    .A2(_11905_),
    .A1(net8431));
 sg13g2_o21ai_1 _20871_ (.B1(net7996),
    .Y(_11907_),
    .A1(_11208_),
    .A2(net8000));
 sg13g2_nor2_1 _20872_ (.A(net8507),
    .B(net8262),
    .Y(_11908_));
 sg13g2_a21oi_1 _20873_ (.A1(net8507),
    .A2(net8255),
    .Y(_11909_),
    .B1(_11908_));
 sg13g2_a22oi_1 _20874_ (.Y(_11910_),
    .B1(_11909_),
    .B2(_11208_),
    .A2(_11907_),
    .A1(net8507));
 sg13g2_o21ai_1 _20875_ (.B1(_11910_),
    .Y(_11911_),
    .A1(net8249),
    .A2(_11897_));
 sg13g2_a221oi_1 _20876_ (.B2(_11906_),
    .C1(_11911_),
    .B1(net7995),
    .A1(_11558_),
    .Y(_11912_),
    .A2(net8267));
 sg13g2_o21ai_1 _20877_ (.B1(net8507),
    .Y(_11913_),
    .A1(net7679),
    .A2(net7677));
 sg13g2_nand3_1 _20878_ (.B(_11912_),
    .C(_11913_),
    .A(_11894_),
    .Y(_11914_));
 sg13g2_o21ai_1 _20879_ (.B1(net7996),
    .Y(_11915_),
    .A1(_11144_),
    .A2(net8000));
 sg13g2_nand2_1 _20880_ (.Y(_11916_),
    .A(_11570_),
    .B(net8265));
 sg13g2_and2_1 _20881_ (.A(net8428),
    .B(_11881_),
    .X(_11917_));
 sg13g2_a21oi_2 _20882_ (.B1(_11917_),
    .Y(_11918_),
    .A2(_11867_),
    .A1(net8415));
 sg13g2_nand2_1 _20883_ (.Y(_11919_),
    .A(net8419),
    .B(_11875_));
 sg13g2_o21ai_1 _20884_ (.B1(_11919_),
    .Y(_11920_),
    .A1(net8417),
    .A2(_11869_));
 sg13g2_nor2_1 _20885_ (.A(net8434),
    .B(_11920_),
    .Y(_11921_));
 sg13g2_a21oi_2 _20886_ (.B1(_11921_),
    .Y(_11922_),
    .A2(_11918_),
    .A1(net8434));
 sg13g2_o21ai_1 _20887_ (.B1(net8429),
    .Y(_11923_),
    .A1(net8391),
    .A2(_11695_));
 sg13g2_a21oi_1 _20888_ (.A1(net8391),
    .A2(_11692_),
    .Y(_11924_),
    .B1(_11923_));
 sg13g2_a21o_1 _20889_ (.A2(_11884_),
    .A1(net8411),
    .B1(_11924_),
    .X(_11925_));
 sg13g2_nor2_1 _20890_ (.A(net8430),
    .B(_11878_),
    .Y(_11926_));
 sg13g2_a21oi_2 _20891_ (.B1(_11926_),
    .Y(_11927_),
    .A2(_11886_),
    .A1(net8430));
 sg13g2_a22oi_1 _20892_ (.Y(_11928_),
    .B1(_11927_),
    .B2(net8245),
    .A2(_11925_),
    .A1(net8253));
 sg13g2_o21ai_1 _20893_ (.B1(_11928_),
    .Y(_11929_),
    .A1(net8446),
    .A2(_11922_));
 sg13g2_nor3_1 _20894_ (.A(net8438),
    .B(net8409),
    .C(_11862_),
    .Y(_11930_));
 sg13g2_o21ai_1 _20895_ (.B1(_11144_),
    .Y(_11931_),
    .A1(net8427),
    .A2(_11645_));
 sg13g2_a21oi_1 _20896_ (.A1(net8427),
    .A2(net8261),
    .Y(_11932_),
    .B1(_11931_));
 sg13g2_a221oi_1 _20897_ (.B2(net7995),
    .C1(_11932_),
    .B1(_11930_),
    .A1(_11705_),
    .Y(_11933_),
    .A2(_11929_));
 sg13g2_nand2_1 _20898_ (.Y(_11934_),
    .A(net8414),
    .B(_11915_));
 sg13g2_nand3_1 _20899_ (.B(_11933_),
    .C(_11934_),
    .A(_11916_),
    .Y(_11935_));
 sg13g2_a221oi_1 _20900_ (.B2(_11144_),
    .C1(_11935_),
    .B1(net7669),
    .A1(net8414),
    .Y(_11936_),
    .A2(net7672));
 sg13g2_o21ai_1 _20901_ (.B1(_11053_),
    .Y(_11937_),
    .A1(_11629_),
    .A2(_11630_));
 sg13g2_o21ai_1 _20902_ (.B1(net8008),
    .Y(_11938_),
    .A1(net7680),
    .A2(net7678));
 sg13g2_a21oi_1 _20903_ (.A1(net8447),
    .A2(_11789_),
    .Y(_11939_),
    .B1(net8249));
 sg13g2_o21ai_1 _20904_ (.B1(_11705_),
    .Y(_11940_),
    .A1(net8442),
    .A2(_11788_));
 sg13g2_a21o_1 _20905_ (.A2(_11876_),
    .A1(net8433),
    .B1(_11895_),
    .X(_11941_));
 sg13g2_nand2_1 _20906_ (.Y(_11942_),
    .A(net8443),
    .B(_11941_));
 sg13g2_nor2_1 _20907_ (.A(net8431),
    .B(_11863_),
    .Y(_11943_));
 sg13g2_o21ai_1 _20908_ (.B1(_11715_),
    .Y(_11944_),
    .A1(net8513),
    .A2(_11268_));
 sg13g2_a21oi_1 _20909_ (.A1(net8383),
    .A2(_11292_),
    .Y(_11945_),
    .B1(_11712_));
 sg13g2_nand2_1 _20910_ (.Y(_11946_),
    .A(net8403),
    .B(_11945_));
 sg13g2_o21ai_1 _20911_ (.B1(_11946_),
    .Y(_11947_),
    .A1(net8406),
    .A2(_11944_));
 sg13g2_o21ai_1 _20912_ (.B1(_11710_),
    .Y(_11948_),
    .A1(net8512),
    .A2(_11222_));
 sg13g2_mux2_1 _20913_ (.A0(_11902_),
    .A1(_11948_),
    .S(net8391),
    .X(_11949_));
 sg13g2_nand2_1 _20914_ (.Y(_11950_),
    .A(net8421),
    .B(_11949_));
 sg13g2_o21ai_1 _20915_ (.B1(_11950_),
    .Y(_11951_),
    .A1(net8420),
    .A2(_11947_));
 sg13g2_a21oi_1 _20916_ (.A1(net8433),
    .A2(_11951_),
    .Y(_11952_),
    .B1(_11943_));
 sg13g2_nand2_1 _20917_ (.Y(_11953_),
    .A(net8447),
    .B(_11952_));
 sg13g2_a21oi_1 _20918_ (.A1(net8386),
    .A2(net8289),
    .Y(_11954_),
    .B1(_11669_));
 sg13g2_o21ai_1 _20919_ (.B1(_11668_),
    .Y(_11955_),
    .A1(net8386),
    .A2(net8279));
 sg13g2_nor2_1 _20920_ (.A(net8396),
    .B(_11955_),
    .Y(_11956_));
 sg13g2_a21oi_1 _20921_ (.A1(net8396),
    .A2(_11954_),
    .Y(_11957_),
    .B1(_11956_));
 sg13g2_nor2b_1 _20922_ (.A(_11662_),
    .B_N(_11664_),
    .Y(_11958_));
 sg13g2_a21oi_1 _20923_ (.A1(net8387),
    .A2(net8283),
    .Y(_11959_),
    .B1(_11717_));
 sg13g2_mux2_1 _20924_ (.A0(_11958_),
    .A1(_11959_),
    .S(net8406),
    .X(_11960_));
 sg13g2_nor2_1 _20925_ (.A(net8423),
    .B(_11957_),
    .Y(_11961_));
 sg13g2_a21oi_2 _20926_ (.B1(_11961_),
    .Y(_11962_),
    .A2(_11960_),
    .A1(net8422));
 sg13g2_o21ai_1 _20927_ (.B1(_11953_),
    .Y(_11963_),
    .A1(_11708_),
    .A2(_11962_));
 sg13g2_nor2_1 _20928_ (.A(_11070_),
    .B(net8264),
    .Y(_11964_));
 sg13g2_o21ai_1 _20929_ (.B1(net7999),
    .Y(_11965_),
    .A1(_11053_),
    .A2(net8002));
 sg13g2_a21oi_1 _20930_ (.A1(net8008),
    .A2(net8257),
    .Y(_11966_),
    .B1(_11964_));
 sg13g2_a22oi_1 _20931_ (.Y(_11967_),
    .B1(_11966_),
    .B2(_11053_),
    .A2(_11965_),
    .A1(net8008));
 sg13g2_o21ai_1 _20932_ (.B1(_11676_),
    .Y(_11968_),
    .A1(net8518),
    .A2(_11440_));
 sg13g2_nor2_1 _20933_ (.A(net8405),
    .B(_11968_),
    .Y(_11969_));
 sg13g2_a21oi_1 _20934_ (.A1(net8386),
    .A2(net8271),
    .Y(_11970_),
    .B1(_11671_));
 sg13g2_a21oi_1 _20935_ (.A1(net8405),
    .A2(_11970_),
    .Y(_11971_),
    .B1(_11969_));
 sg13g2_inv_1 _20936_ (.Y(_11972_),
    .A(_11971_));
 sg13g2_a21oi_1 _20937_ (.A1(net8385),
    .A2(net8269),
    .Y(_11973_),
    .B1(_11678_));
 sg13g2_nand3_1 _20938_ (.B(_11682_),
    .C(_11684_),
    .A(net8394),
    .Y(_11974_));
 sg13g2_a21oi_1 _20939_ (.A1(net8404),
    .A2(_11973_),
    .Y(_11975_),
    .B1(net8418));
 sg13g2_a22oi_1 _20940_ (.Y(_11976_),
    .B1(_11974_),
    .B2(_11975_),
    .A2(_11971_),
    .A1(net8419));
 sg13g2_nand2_1 _20941_ (.Y(_11977_),
    .A(_11864_),
    .B(_11976_));
 sg13g2_nand2_1 _20942_ (.Y(_11978_),
    .A(_11967_),
    .B(_11977_));
 sg13g2_nor2_2 _20943_ (.A(net8445),
    .B(_11655_),
    .Y(_11979_));
 sg13g2_a221oi_1 _20944_ (.B2(_11654_),
    .C1(_11978_),
    .B1(_11963_),
    .A1(net7936),
    .Y(_11980_),
    .A2(_11942_));
 sg13g2_nand2b_1 _20945_ (.Y(_11981_),
    .B(net8266),
    .A_N(_11508_));
 sg13g2_nand4_1 _20946_ (.B(_11938_),
    .C(_11980_),
    .A(_11937_),
    .Y(_11982_),
    .D(_11981_));
 sg13g2_o21ai_1 _20947_ (.B1(net8382),
    .Y(_11983_),
    .A1(net7679),
    .A2(net7677));
 sg13g2_a21oi_1 _20948_ (.A1(_10993_),
    .A2(_11649_),
    .Y(_11984_),
    .B1(_11788_));
 sg13g2_nand2_1 _20949_ (.Y(_11985_),
    .A(net8416),
    .B(_11984_));
 sg13g2_nand2_1 _20950_ (.Y(_11986_),
    .A(net8393),
    .B(_11782_));
 sg13g2_o21ai_1 _20951_ (.B1(_11986_),
    .Y(_11987_),
    .A1(net8393),
    .A2(_11786_));
 sg13g2_o21ai_1 _20952_ (.B1(_11985_),
    .Y(_11988_),
    .A1(net8416),
    .A2(_11987_));
 sg13g2_a21oi_2 _20953_ (.B1(net7938),
    .Y(_11989_),
    .A2(_11988_),
    .A1(net8432));
 sg13g2_nor2_1 _20954_ (.A(net8404),
    .B(_11766_),
    .Y(_11990_));
 sg13g2_a21oi_2 _20955_ (.B1(_11990_),
    .Y(_11991_),
    .A2(_11770_),
    .A1(net8404));
 sg13g2_nand2b_1 _20956_ (.Y(_11992_),
    .B(net8395),
    .A_N(_11774_));
 sg13g2_o21ai_1 _20957_ (.B1(_11992_),
    .Y(_11993_),
    .A1(net8394),
    .A2(_11780_));
 sg13g2_nor2_1 _20958_ (.A(net8429),
    .B(_11993_),
    .Y(_11994_));
 sg13g2_a21oi_1 _20959_ (.A1(net8428),
    .A2(_11991_),
    .Y(_11995_),
    .B1(_11994_));
 sg13g2_nor2_1 _20960_ (.A(net8392),
    .B(_11818_),
    .Y(_11996_));
 sg13g2_a21oi_1 _20961_ (.A1(net8392),
    .A2(_11812_),
    .Y(_11997_),
    .B1(_11996_));
 sg13g2_mux2_1 _20962_ (.A0(_11764_),
    .A1(_11820_),
    .S(net8397),
    .X(_11998_));
 sg13g2_nor2_1 _20963_ (.A(net8413),
    .B(_11997_),
    .Y(_11999_));
 sg13g2_a21oi_1 _20964_ (.A1(net8413),
    .A2(_11998_),
    .Y(_12000_),
    .B1(_11999_));
 sg13g2_nor2_1 _20965_ (.A(net8251),
    .B(_12000_),
    .Y(_12001_));
 sg13g2_a221oi_1 _20966_ (.B2(net8246),
    .C1(_12001_),
    .B1(_11995_),
    .A1(net8451),
    .Y(_12002_),
    .A2(_11989_));
 sg13g2_a21oi_1 _20967_ (.A1(_11143_),
    .A2(net8509),
    .Y(_12003_),
    .B1(_11795_));
 sg13g2_nor2_1 _20968_ (.A(net8390),
    .B(_11827_),
    .Y(_12004_));
 sg13g2_a21oi_2 _20969_ (.B1(_12004_),
    .Y(_12005_),
    .A2(_12003_),
    .A1(net8390));
 sg13g2_nand2b_2 _20970_ (.Y(_12006_),
    .B(net8427),
    .A_N(_12005_));
 sg13g2_a21oi_1 _20971_ (.A1(_11097_),
    .A2(net8508),
    .Y(_12007_),
    .B1(_11804_));
 sg13g2_nand2_1 _20972_ (.Y(_12008_),
    .A(net8389),
    .B(_12007_));
 sg13g2_o21ai_1 _20973_ (.B1(_11796_),
    .Y(_12009_),
    .A1(net8304),
    .A2(net8509));
 sg13g2_o21ai_1 _20974_ (.B1(_12008_),
    .Y(_12010_),
    .A1(net8389),
    .A2(_12009_));
 sg13g2_nand2_1 _20975_ (.Y(_12011_),
    .A(net8410),
    .B(_12010_));
 sg13g2_a21oi_2 _20976_ (.B1(_11811_),
    .Y(_12012_),
    .A2(_11221_),
    .A1(net8512));
 sg13g2_o21ai_1 _20977_ (.B1(_11809_),
    .Y(_12013_),
    .A1(net8383),
    .A2(_11208_));
 sg13g2_nor2_1 _20978_ (.A(net8389),
    .B(_12013_),
    .Y(_12014_));
 sg13g2_a21oi_2 _20979_ (.B1(_12014_),
    .Y(_12015_),
    .A2(_12012_),
    .A1(net8390));
 sg13g2_o21ai_1 _20980_ (.B1(_12011_),
    .Y(_12016_),
    .A1(net8414),
    .A2(_12015_));
 sg13g2_nor2_1 _20981_ (.A(net8440),
    .B(_12016_),
    .Y(_12017_));
 sg13g2_a21oi_2 _20982_ (.B1(_12017_),
    .Y(_12018_),
    .A2(_12006_),
    .A1(net8438));
 sg13g2_nor2_1 _20983_ (.A(net8382),
    .B(net8262),
    .Y(_12019_));
 sg13g2_a21oi_1 _20984_ (.A1(net8382),
    .A2(net8256),
    .Y(_12020_),
    .B1(_12019_));
 sg13g2_o21ai_1 _20985_ (.B1(net7999),
    .Y(_12021_),
    .A1(net8296),
    .A2(net8003));
 sg13g2_a22oi_1 _20986_ (.Y(_12022_),
    .B1(_12020_),
    .B2(net8296),
    .A2(_12018_),
    .A1(net7995));
 sg13g2_o21ai_1 _20987_ (.B1(_12022_),
    .Y(_12023_),
    .A1(net8249),
    .A2(_12002_));
 sg13g2_a221oi_1 _20988_ (.B2(net8382),
    .C1(_12023_),
    .B1(_12021_),
    .A1(_11551_),
    .Y(_12024_),
    .A2(net8265));
 sg13g2_o21ai_1 _20989_ (.B1(net8296),
    .Y(_12025_),
    .A1(net7676),
    .A2(net7675));
 sg13g2_nand3_1 _20990_ (.B(_12024_),
    .C(_12025_),
    .A(_11983_),
    .Y(_12026_));
 sg13g2_o21ai_1 _20991_ (.B1(net8522),
    .Y(_12027_),
    .A1(net7679),
    .A2(net7677));
 sg13g2_o21ai_1 _20992_ (.B1(net7996),
    .Y(_12028_),
    .A1(_11086_),
    .A2(net8000));
 sg13g2_a21oi_1 _20993_ (.A1(net8522),
    .A2(net8255),
    .Y(_12029_),
    .B1(_11087_));
 sg13g2_nand2b_1 _20994_ (.Y(_12030_),
    .B(net8261),
    .A_N(net8522));
 sg13g2_a21o_1 _20995_ (.A2(_12028_),
    .A1(net8522),
    .B1(_12029_),
    .X(_12031_));
 sg13g2_nor2_1 _20996_ (.A(net8410),
    .B(_12010_),
    .Y(_12032_));
 sg13g2_a21oi_2 _20997_ (.B1(_12032_),
    .Y(_12033_),
    .A2(_12005_),
    .A1(net8409));
 sg13g2_and2_1 _20998_ (.A(net8419),
    .B(_11987_),
    .X(_12034_));
 sg13g2_a21oi_1 _20999_ (.A1(net8428),
    .A2(_11993_),
    .Y(_12035_),
    .B1(_12034_));
 sg13g2_nor2_1 _21000_ (.A(net8439),
    .B(_12035_),
    .Y(_12036_));
 sg13g2_nor2_1 _21001_ (.A(_11873_),
    .B(_11984_),
    .Y(_12037_));
 sg13g2_a21oi_1 _21002_ (.A1(net8439),
    .A2(_12037_),
    .Y(_12038_),
    .B1(_12036_));
 sg13g2_nor2_1 _21003_ (.A(net8413),
    .B(_11998_),
    .Y(_12039_));
 sg13g2_a21oi_1 _21004_ (.A1(net8415),
    .A2(_11991_),
    .Y(_12040_),
    .B1(_12039_));
 sg13g2_nand2_1 _21005_ (.Y(_12041_),
    .A(net8391),
    .B(_11805_));
 sg13g2_o21ai_1 _21006_ (.B1(_12041_),
    .Y(_12042_),
    .A1(net8389),
    .A2(_11810_));
 sg13g2_nor2_1 _21007_ (.A(net8411),
    .B(_12042_),
    .Y(_12043_));
 sg13g2_a21oi_1 _21008_ (.A1(net8413),
    .A2(_11997_),
    .Y(_12044_),
    .B1(_12043_));
 sg13g2_a22oi_1 _21009_ (.Y(_12045_),
    .B1(_12044_),
    .B2(net8253),
    .A2(_12040_),
    .A1(net8246));
 sg13g2_o21ai_1 _21010_ (.B1(_12045_),
    .Y(_12046_),
    .A1(net8444),
    .A2(_12038_));
 sg13g2_nand2_1 _21011_ (.Y(_12047_),
    .A(_11705_),
    .B(_12046_));
 sg13g2_o21ai_1 _21012_ (.B1(_12047_),
    .Y(_12048_),
    .A1(_11562_),
    .A2(net8004));
 sg13g2_a221oi_1 _21013_ (.B2(_11864_),
    .C1(_12048_),
    .B1(_12033_),
    .A1(_12030_),
    .Y(_12049_),
    .A2(_12031_));
 sg13g2_o21ai_1 _21014_ (.B1(_11086_),
    .Y(_12050_),
    .A1(net7676),
    .A2(net7675));
 sg13g2_and3_2 _21015_ (.X(_12051_),
    .A(_12027_),
    .B(_12049_),
    .C(_12050_));
 sg13g2_nand3_1 _21016_ (.B(_12049_),
    .C(_12050_),
    .A(_12027_),
    .Y(_12052_));
 sg13g2_nand2_1 _21017_ (.Y(_12053_),
    .A(net8427),
    .B(_11949_));
 sg13g2_o21ai_1 _21018_ (.B1(_12053_),
    .Y(_12054_),
    .A1(net8429),
    .A2(_11858_));
 sg13g2_or3_1 _21019_ (.A(net8431),
    .B(net8409),
    .C(_11862_),
    .X(_12055_));
 sg13g2_o21ai_1 _21020_ (.B1(_12055_),
    .Y(_12056_),
    .A1(net8438),
    .A2(_12054_));
 sg13g2_o21ai_1 _21021_ (.B1(net7996),
    .Y(_12057_),
    .A1(_11222_),
    .A2(net8000));
 sg13g2_o21ai_1 _21022_ (.B1(_11222_),
    .Y(_12058_),
    .A1(net8506),
    .A2(net8264));
 sg13g2_a21oi_1 _21023_ (.A1(net8506),
    .A2(net8255),
    .Y(_12059_),
    .B1(_12058_));
 sg13g2_a221oi_1 _21024_ (.B2(net8506),
    .C1(_12059_),
    .B1(_12057_),
    .A1(net7995),
    .Y(_12060_),
    .A2(_12056_));
 sg13g2_a21oi_1 _21025_ (.A1(net8434),
    .A2(_11920_),
    .Y(_12061_),
    .B1(net7938));
 sg13g2_nand2_1 _21026_ (.Y(_12062_),
    .A(net8451),
    .B(_12061_));
 sg13g2_a22oi_1 _21027_ (.Y(_12063_),
    .B1(_11927_),
    .B2(net8253),
    .A2(_11918_),
    .A1(net8245));
 sg13g2_a21oi_1 _21028_ (.A1(_12062_),
    .A2(_12063_),
    .Y(_12064_),
    .B1(net8250));
 sg13g2_nor2b_1 _21029_ (.A(_12064_),
    .B_N(_12060_),
    .Y(_12065_));
 sg13g2_o21ai_1 _21030_ (.B1(_12065_),
    .Y(_12066_),
    .A1(_11554_),
    .A2(net8004));
 sg13g2_a21oi_1 _21031_ (.A1(net8506),
    .A2(net7672),
    .Y(_12067_),
    .B1(_12066_));
 sg13g2_a221oi_1 _21032_ (.B2(_11222_),
    .C1(_12066_),
    .B1(net7669),
    .A1(net8506),
    .Y(_12068_),
    .A2(net7672));
 sg13g2_o21ai_1 _21033_ (.B1(_12067_),
    .Y(_12069_),
    .A1(_11221_),
    .A2(_11632_));
 sg13g2_o21ai_1 _21034_ (.B1(_11465_),
    .Y(_12070_),
    .A1(net7679),
    .A2(net7678));
 sg13g2_nand2_1 _21035_ (.Y(_12071_),
    .A(_11581_),
    .B(net8266));
 sg13g2_o21ai_1 _21036_ (.B1(net7936),
    .Y(_12072_),
    .A1(net8447),
    .A2(_11896_));
 sg13g2_a21oi_2 _21037_ (.B1(net8258),
    .Y(_12073_),
    .A2(net8263),
    .A1(_10965_));
 sg13g2_nand2_1 _21038_ (.Y(_12074_),
    .A(_11641_),
    .B(net8257));
 sg13g2_o21ai_1 _21039_ (.B1(_10881_),
    .Y(_12075_),
    .A1(net8271),
    .A2(_12073_));
 sg13g2_a22oi_1 _21040_ (.Y(_12076_),
    .B1(_12075_),
    .B2(_11465_),
    .A2(_11979_),
    .A1(_11906_));
 sg13g2_xnor2_1 _21041_ (.Y(_12077_),
    .A(_11463_),
    .B(_11465_));
 sg13g2_o21ai_1 _21042_ (.B1(_12076_),
    .Y(_12078_),
    .A1(net8260),
    .A2(_12077_));
 sg13g2_nor2_1 _21043_ (.A(net8391),
    .B(_11948_),
    .Y(_12079_));
 sg13g2_a21oi_2 _21044_ (.B1(_12079_),
    .Y(_12080_),
    .A2(_11945_),
    .A1(net8392));
 sg13g2_nand2_1 _21045_ (.Y(_12081_),
    .A(net8397),
    .B(_11959_));
 sg13g2_o21ai_1 _21046_ (.B1(_12081_),
    .Y(_12082_),
    .A1(net8397),
    .A2(_11944_));
 sg13g2_nor2_1 _21047_ (.A(net8422),
    .B(_12082_),
    .Y(_12083_));
 sg13g2_a21oi_2 _21048_ (.B1(_12083_),
    .Y(_12084_),
    .A2(_12080_),
    .A1(net8421));
 sg13g2_mux2_1 _21049_ (.A0(_11954_),
    .A1(_11970_),
    .S(net8396),
    .X(_12085_));
 sg13g2_inv_1 _21050_ (.Y(_12086_),
    .A(_12085_));
 sg13g2_nor2_1 _21051_ (.A(net8406),
    .B(_11955_),
    .Y(_12087_));
 sg13g2_a21oi_2 _21052_ (.B1(_12087_),
    .Y(_12088_),
    .A2(_11958_),
    .A1(net8406));
 sg13g2_o21ai_1 _21053_ (.B1(net8437),
    .Y(_12089_),
    .A1(net8423),
    .A2(_12085_));
 sg13g2_a21oi_1 _21054_ (.A1(net8423),
    .A2(_12088_),
    .Y(_12090_),
    .B1(_12089_));
 sg13g2_a21oi_1 _21055_ (.A1(net8441),
    .A2(_12084_),
    .Y(_12091_),
    .B1(_12090_));
 sg13g2_o21ai_1 _21056_ (.B1(_12072_),
    .Y(_12092_),
    .A1(net7994),
    .A2(_12091_));
 sg13g2_nor2_1 _21057_ (.A(_12078_),
    .B(_12092_),
    .Y(_12093_));
 sg13g2_o21ai_1 _21058_ (.B1(_11463_),
    .Y(_12094_),
    .A1(net7676),
    .A2(net7675));
 sg13g2_nand4_1 _21059_ (.B(_12071_),
    .C(_12093_),
    .A(_12070_),
    .Y(_12095_),
    .D(_12094_));
 sg13g2_o21ai_1 _21060_ (.B1(_11476_),
    .Y(_12096_),
    .A1(net7680),
    .A2(net7678));
 sg13g2_nand2b_1 _21061_ (.Y(_12097_),
    .B(net8266),
    .A_N(_11543_));
 sg13g2_a21o_1 _21062_ (.A2(_11793_),
    .A1(net8433),
    .B1(net7938),
    .X(_12098_));
 sg13g2_nand2_1 _21063_ (.Y(_12099_),
    .A(net8442),
    .B(_12098_));
 sg13g2_o21ai_1 _21064_ (.B1(_11816_),
    .Y(_12100_),
    .A1(net8383),
    .A2(net8292));
 sg13g2_nor2_1 _21065_ (.A(net8402),
    .B(_12100_),
    .Y(_12101_));
 sg13g2_a21oi_1 _21066_ (.A1(net8403),
    .A2(_12012_),
    .Y(_12102_),
    .B1(_12101_));
 sg13g2_nor2_1 _21067_ (.A(net8429),
    .B(_12102_),
    .Y(_12103_));
 sg13g2_a21oi_1 _21068_ (.A1(net8517),
    .A2(net8283),
    .Y(_12104_),
    .B1(_11762_));
 sg13g2_nand2_1 _21069_ (.Y(_12105_),
    .A(net8397),
    .B(_12104_));
 sg13g2_o21ai_1 _21070_ (.B1(_11817_),
    .Y(_12106_),
    .A1(net8513),
    .A2(net8294));
 sg13g2_o21ai_1 _21071_ (.B1(_12105_),
    .Y(_12107_),
    .A1(net8397),
    .A2(_12106_));
 sg13g2_a21oi_2 _21072_ (.B1(_12103_),
    .Y(_12108_),
    .A2(_12107_),
    .A1(net8428));
 sg13g2_nand2_1 _21073_ (.Y(_12109_),
    .A(_11773_),
    .B(_11779_));
 sg13g2_nor2_1 _21074_ (.A(net8404),
    .B(_12109_),
    .Y(_12110_));
 sg13g2_a21oi_1 _21075_ (.A1(net8515),
    .A2(net8288),
    .Y(_12111_),
    .B1(_11772_));
 sg13g2_a21oi_1 _21076_ (.A1(net8405),
    .A2(_12111_),
    .Y(_12112_),
    .B1(_12110_));
 sg13g2_inv_1 _21077_ (.Y(_12113_),
    .A(_12112_));
 sg13g2_a21oi_1 _21078_ (.A1(net8516),
    .A2(net8286),
    .Y(_12114_),
    .B1(_11769_));
 sg13g2_o21ai_1 _21079_ (.B1(_11763_),
    .Y(_12115_),
    .A1(net8515),
    .A2(net8279));
 sg13g2_nor2_1 _21080_ (.A(net8395),
    .B(_12115_),
    .Y(_12116_));
 sg13g2_a21oi_1 _21081_ (.A1(net8395),
    .A2(_12114_),
    .Y(_12117_),
    .B1(_12116_));
 sg13g2_a21oi_1 _21082_ (.A1(net8418),
    .A2(_12117_),
    .Y(_12118_),
    .B1(net8439));
 sg13g2_o21ai_1 _21083_ (.B1(_12118_),
    .Y(_12119_),
    .A1(net8417),
    .A2(_12113_));
 sg13g2_o21ai_1 _21084_ (.B1(_12119_),
    .Y(_12120_),
    .A1(net8434),
    .A2(_12108_));
 sg13g2_nand2_1 _21085_ (.Y(_12121_),
    .A(net8400),
    .B(_12003_));
 sg13g2_o21ai_1 _21086_ (.B1(_12121_),
    .Y(_12122_),
    .A1(net8400),
    .A2(_12009_));
 sg13g2_nor2_1 _21087_ (.A(net8401),
    .B(_12013_),
    .Y(_12123_));
 sg13g2_a21oi_2 _21088_ (.B1(_12123_),
    .Y(_12124_),
    .A2(_12007_),
    .A1(net8401));
 sg13g2_nor2_1 _21089_ (.A(net8410),
    .B(_12124_),
    .Y(_12125_));
 sg13g2_a21oi_2 _21090_ (.B1(_12125_),
    .Y(_12126_),
    .A2(_12122_),
    .A1(net8410));
 sg13g2_nand2_1 _21091_ (.Y(_12127_),
    .A(net8431),
    .B(_12126_));
 sg13g2_o21ai_1 _21092_ (.B1(_12127_),
    .Y(_12128_),
    .A1(net8431),
    .A2(_11829_));
 sg13g2_inv_1 _21093_ (.Y(_12129_),
    .A(_12128_));
 sg13g2_xnor2_1 _21094_ (.Y(_12130_),
    .A(_11473_),
    .B(_11476_));
 sg13g2_o21ai_1 _21095_ (.B1(_10881_),
    .Y(_12131_),
    .A1(_11472_),
    .A2(_12073_));
 sg13g2_a22oi_1 _21096_ (.Y(_12132_),
    .B1(_12131_),
    .B2(_11476_),
    .A2(_12129_),
    .A1(_11979_));
 sg13g2_o21ai_1 _21097_ (.B1(_12132_),
    .Y(_12133_),
    .A1(net8260),
    .A2(_12130_));
 sg13g2_a221oi_1 _21098_ (.B2(net7995),
    .C1(_12133_),
    .B1(_12120_),
    .A1(net7936),
    .Y(_12134_),
    .A2(_12099_));
 sg13g2_o21ai_1 _21099_ (.B1(_11473_),
    .Y(_12135_),
    .A1(_11629_),
    .A2(_11630_));
 sg13g2_nand4_1 _21100_ (.B(_12097_),
    .C(_12134_),
    .A(_12096_),
    .Y(_12136_),
    .D(_12135_));
 sg13g2_o21ai_1 _21101_ (.B1(net7998),
    .Y(_12137_),
    .A1(_11492_),
    .A2(net8002));
 sg13g2_o21ai_1 _21102_ (.B1(_11492_),
    .Y(_12138_),
    .A1(_11629_),
    .A2(_11630_));
 sg13g2_nand2b_1 _21103_ (.Y(_12139_),
    .B(net8266),
    .A_N(_11544_));
 sg13g2_nand2_1 _21104_ (.Y(_12140_),
    .A(net8410),
    .B(_11652_));
 sg13g2_o21ai_1 _21105_ (.B1(_12140_),
    .Y(_12141_),
    .A1(net8409),
    .A2(_11900_));
 sg13g2_nand2_1 _21106_ (.Y(_12142_),
    .A(net8440),
    .B(_12141_));
 sg13g2_nand2_1 _21107_ (.Y(_12143_),
    .A(net8421),
    .B(_11904_));
 sg13g2_o21ai_1 _21108_ (.B1(_12143_),
    .Y(_12144_),
    .A1(net8420),
    .A2(_12080_));
 sg13g2_o21ai_1 _21109_ (.B1(_12142_),
    .Y(_12145_),
    .A1(net8440),
    .A2(_12144_));
 sg13g2_nor2_1 _21110_ (.A(net8430),
    .B(_12082_),
    .Y(_12146_));
 sg13g2_a21oi_2 _21111_ (.B1(_12146_),
    .Y(_12147_),
    .A2(_12088_),
    .A1(net8430));
 sg13g2_a21oi_1 _21112_ (.A1(net8394),
    .A2(_11973_),
    .Y(_12148_),
    .B1(net8418));
 sg13g2_o21ai_1 _21113_ (.B1(_12148_),
    .Y(_12149_),
    .A1(net8394),
    .A2(_11968_));
 sg13g2_a21oi_1 _21114_ (.A1(net8417),
    .A2(_12086_),
    .Y(_12150_),
    .B1(net8251));
 sg13g2_a22oi_1 _21115_ (.Y(_12151_),
    .B1(_12149_),
    .B2(_12150_),
    .A2(_12147_),
    .A1(net8248));
 sg13g2_o21ai_1 _21116_ (.B1(_12151_),
    .Y(_12152_),
    .A1(net8442),
    .A2(_12145_));
 sg13g2_a21oi_1 _21117_ (.A1(_11495_),
    .A2(net8259),
    .Y(_12153_),
    .B1(net8268));
 sg13g2_o21ai_1 _21118_ (.B1(_12153_),
    .Y(_12154_),
    .A1(_11495_),
    .A2(net8258));
 sg13g2_a21o_1 _21119_ (.A2(_11686_),
    .A1(net8428),
    .B1(_11873_),
    .X(_12155_));
 sg13g2_a21oi_2 _21120_ (.B1(net7938),
    .Y(_12156_),
    .A2(_12155_),
    .A1(net8433));
 sg13g2_o21ai_1 _21121_ (.B1(net7937),
    .Y(_12157_),
    .A1(net8450),
    .A2(_12156_));
 sg13g2_nand2_1 _21122_ (.Y(_12158_),
    .A(_11496_),
    .B(_12137_));
 sg13g2_nand3_1 _21123_ (.B(_12157_),
    .C(_12158_),
    .A(_12154_),
    .Y(_12159_));
 sg13g2_a21oi_1 _21124_ (.A1(_11654_),
    .A2(_12152_),
    .Y(_12160_),
    .B1(_12159_));
 sg13g2_o21ai_1 _21125_ (.B1(_11496_),
    .Y(_12161_),
    .A1(net7680),
    .A2(net7678));
 sg13g2_nand4_1 _21126_ (.B(_12139_),
    .C(_12160_),
    .A(_12138_),
    .Y(_12162_),
    .D(_12161_));
 sg13g2_o21ai_1 _21127_ (.B1(_11350_),
    .Y(_12163_),
    .A1(net7676),
    .A2(net7675));
 sg13g2_mux2_2 _21128_ (.A0(_11673_),
    .A1(_11681_),
    .S(net8415),
    .X(_12164_));
 sg13g2_nor2_1 _21129_ (.A(net8435),
    .B(_12155_),
    .Y(_12165_));
 sg13g2_a21oi_2 _21130_ (.B1(_12165_),
    .Y(_12166_),
    .A2(_12164_),
    .A1(net8433));
 sg13g2_nand2_1 _21131_ (.Y(_12167_),
    .A(net8443),
    .B(_12166_));
 sg13g2_o21ai_1 _21132_ (.B1(net7994),
    .Y(_12168_),
    .A1(_11657_),
    .A2(_12141_));
 sg13g2_nor2_1 _21133_ (.A(_11708_),
    .B(_12144_),
    .Y(_12169_));
 sg13g2_nor2_1 _21134_ (.A(_11701_),
    .B(_12147_),
    .Y(_12170_));
 sg13g2_nor2_1 _21135_ (.A(_12169_),
    .B(_12170_),
    .Y(_12171_));
 sg13g2_a21oi_1 _21136_ (.A1(_11353_),
    .A2(net8257),
    .Y(_12172_),
    .B1(net8286));
 sg13g2_o21ai_1 _21137_ (.B1(_12172_),
    .Y(_12173_),
    .A1(_11353_),
    .A2(net8263));
 sg13g2_o21ai_1 _21138_ (.B1(net7999),
    .Y(_12174_),
    .A1(_11350_),
    .A2(net8003));
 sg13g2_a22oi_1 _21139_ (.Y(_12175_),
    .B1(_12174_),
    .B2(_11353_),
    .A2(_12167_),
    .A1(net7936));
 sg13g2_nand2_1 _21140_ (.Y(_12176_),
    .A(_12173_),
    .B(_12175_));
 sg13g2_a221oi_1 _21141_ (.B2(_12171_),
    .C1(_12176_),
    .B1(_12168_),
    .A1(_11521_),
    .Y(_12177_),
    .A2(net8267));
 sg13g2_o21ai_1 _21142_ (.B1(_11353_),
    .Y(_12178_),
    .A1(net7679),
    .A2(net7677));
 sg13g2_and3_2 _21143_ (.X(_12179_),
    .A(_12163_),
    .B(_12177_),
    .C(_12178_));
 sg13g2_nand3_1 _21144_ (.B(_12177_),
    .C(_12178_),
    .A(_12163_),
    .Y(_12180_));
 sg13g2_nor2_1 _21145_ (.A(net8439),
    .B(_12037_),
    .Y(_12181_));
 sg13g2_o21ai_1 _21146_ (.B1(net8442),
    .Y(_12182_),
    .A1(net7938),
    .A2(_12181_));
 sg13g2_o21ai_1 _21147_ (.B1(_11599_),
    .Y(_12183_),
    .A1(_11611_),
    .A2(net8258));
 sg13g2_a22oi_1 _21148_ (.Y(_12184_),
    .B1(_11598_),
    .B2(_11619_),
    .A2(_11021_),
    .A1(_10880_));
 sg13g2_nand4_1 _21149_ (.B(_11641_),
    .C(_12183_),
    .A(_11621_),
    .Y(_12185_),
    .D(_12184_));
 sg13g2_a22oi_1 _21150_ (.Y(_12186_),
    .B1(_12185_),
    .B2(_11597_),
    .A2(_12182_),
    .A1(net7937));
 sg13g2_nor2_1 _21151_ (.A(net8432),
    .B(_12033_),
    .Y(_12187_));
 sg13g2_mux2_1 _21152_ (.A0(_12100_),
    .A1(_12106_),
    .S(net8392),
    .X(_12188_));
 sg13g2_mux2_1 _21153_ (.A0(_12015_),
    .A1(_12188_),
    .S(net8429),
    .X(_12189_));
 sg13g2_a21oi_2 _21154_ (.B1(_12187_),
    .Y(_12190_),
    .A2(_12189_),
    .A1(net8432));
 sg13g2_a21oi_1 _21155_ (.A1(net8514),
    .A2(net8275),
    .Y(_12191_),
    .B1(_11781_));
 sg13g2_nand2_1 _21156_ (.Y(_12192_),
    .A(net8394),
    .B(_12191_));
 sg13g2_o21ai_1 _21157_ (.B1(_12192_),
    .Y(_12193_),
    .A1(net8394),
    .A2(_12109_));
 sg13g2_nand2_1 _21158_ (.Y(_12194_),
    .A(net8419),
    .B(_12193_));
 sg13g2_a21oi_1 _21159_ (.A1(net8315),
    .A2(_11649_),
    .Y(_12195_),
    .B1(net8419));
 sg13g2_o21ai_1 _21160_ (.B1(_11785_),
    .Y(_12196_),
    .A1(net8384),
    .A2(_11492_));
 sg13g2_nor3_1 _21161_ (.A(_11053_),
    .B(net8408),
    .C(net8384),
    .Y(_12197_));
 sg13g2_a21oi_1 _21162_ (.A1(net8408),
    .A2(_12196_),
    .Y(_12198_),
    .B1(_12197_));
 sg13g2_a21oi_1 _21163_ (.A1(_12195_),
    .A2(_12198_),
    .Y(_12199_),
    .B1(_11701_));
 sg13g2_nand2_1 _21164_ (.Y(_12200_),
    .A(net8406),
    .B(_12104_));
 sg13g2_o21ai_1 _21165_ (.B1(_12200_),
    .Y(_12201_),
    .A1(net8405),
    .A2(_12115_));
 sg13g2_and2_1 _21166_ (.A(net8395),
    .B(_12111_),
    .X(_12202_));
 sg13g2_a21oi_1 _21167_ (.A1(net8405),
    .A2(_12114_),
    .Y(_12203_),
    .B1(_12202_));
 sg13g2_nor2_1 _21168_ (.A(net8418),
    .B(_12203_),
    .Y(_12204_));
 sg13g2_a21oi_1 _21169_ (.A1(net8418),
    .A2(_12201_),
    .Y(_12205_),
    .B1(_12204_));
 sg13g2_a221oi_1 _21170_ (.B2(net8248),
    .C1(_11655_),
    .B1(_12205_),
    .A1(_12194_),
    .Y(_12206_),
    .A2(_12199_));
 sg13g2_o21ai_1 _21171_ (.B1(_12206_),
    .Y(_12207_),
    .A1(net8445),
    .A2(_12190_));
 sg13g2_nand2_1 _21172_ (.Y(_12208_),
    .A(_12186_),
    .B(_12207_));
 sg13g2_a221oi_1 _21173_ (.B2(_10993_),
    .C1(_12208_),
    .B1(_11627_),
    .A1(_11021_),
    .Y(_12209_),
    .A2(net7680));
 sg13g2_o21ai_1 _21174_ (.B1(_12209_),
    .Y(_12210_),
    .A1(_11507_),
    .A2(net8005));
 sg13g2_o21ai_1 _21175_ (.B1(_11454_),
    .Y(_12211_),
    .A1(net7680),
    .A2(net7677));
 sg13g2_or2_1 _21176_ (.X(_12212_),
    .B(_11989_),
    .A(net8450));
 sg13g2_o21ai_1 _21177_ (.B1(net8273),
    .Y(_12213_),
    .A1(_11453_),
    .A2(_12074_));
 sg13g2_a21oi_1 _21178_ (.A1(_11453_),
    .A2(net8259),
    .Y(_12214_),
    .B1(_12213_));
 sg13g2_o21ai_1 _21179_ (.B1(_10881_),
    .Y(_12215_),
    .A1(net8273),
    .A2(net8259));
 sg13g2_a221oi_1 _21180_ (.B2(_11454_),
    .C1(_12214_),
    .B1(_12215_),
    .A1(_11979_),
    .Y(_12216_),
    .A2(_12018_));
 sg13g2_o21ai_1 _21181_ (.B1(net8435),
    .Y(_12217_),
    .A1(net8417),
    .A2(_12193_));
 sg13g2_a21oi_1 _21182_ (.A1(net8417),
    .A2(_12203_),
    .Y(_12218_),
    .B1(_12217_));
 sg13g2_nor2_1 _21183_ (.A(net8415),
    .B(_12201_),
    .Y(_12219_));
 sg13g2_a21oi_2 _21184_ (.B1(_12219_),
    .Y(_12220_),
    .A2(_12188_),
    .A1(net8415));
 sg13g2_a21oi_1 _21185_ (.A1(net8440),
    .A2(_12220_),
    .Y(_12221_),
    .B1(_12218_));
 sg13g2_o21ai_1 _21186_ (.B1(_12216_),
    .Y(_12222_),
    .A1(net7994),
    .A2(_12221_));
 sg13g2_a221oi_1 _21187_ (.B2(_12212_),
    .C1(_12222_),
    .B1(net7937),
    .A1(_11513_),
    .Y(_12223_),
    .A2(net8266));
 sg13g2_o21ai_1 _21188_ (.B1(net8273),
    .Y(_12224_),
    .A1(net7676),
    .A2(net7675));
 sg13g2_nand3_1 _21189_ (.B(_12223_),
    .C(_12224_),
    .A(_12211_),
    .Y(_12225_));
 sg13g2_or2_1 _21190_ (.X(_12226_),
    .B(_12061_),
    .A(net8451));
 sg13g2_o21ai_1 _21191_ (.B1(_10881_),
    .Y(_12227_),
    .A1(_11440_),
    .A2(net8260));
 sg13g2_nand2_1 _21192_ (.Y(_12228_),
    .A(net8006),
    .B(_12073_));
 sg13g2_o21ai_1 _21193_ (.B1(_12228_),
    .Y(_12229_),
    .A1(net8006),
    .A2(net8263));
 sg13g2_nor2_1 _21194_ (.A(_11439_),
    .B(_12229_),
    .Y(_12230_));
 sg13g2_a221oi_1 _21195_ (.B2(net8006),
    .C1(_12230_),
    .B1(_12227_),
    .A1(_11979_),
    .Y(_12231_),
    .A2(_12056_));
 sg13g2_a21oi_1 _21196_ (.A1(net8422),
    .A2(_11957_),
    .Y(_12232_),
    .B1(net8441));
 sg13g2_o21ai_1 _21197_ (.B1(_12232_),
    .Y(_12233_),
    .A1(net8423),
    .A2(_11972_));
 sg13g2_or2_1 _21198_ (.X(_12234_),
    .B(_11960_),
    .A(net8422));
 sg13g2_o21ai_1 _21199_ (.B1(_12234_),
    .Y(_12235_),
    .A1(_11152_),
    .A2(_11947_));
 sg13g2_o21ai_1 _21200_ (.B1(_12233_),
    .Y(_12236_),
    .A1(net8437),
    .A2(_12235_));
 sg13g2_a22oi_1 _21201_ (.Y(_12237_),
    .B1(_12236_),
    .B2(_11660_),
    .A2(_12226_),
    .A1(net7936));
 sg13g2_a21oi_1 _21202_ (.A1(_11514_),
    .A2(_11515_),
    .Y(_12238_),
    .B1(net8005));
 sg13g2_nand3b_1 _21203_ (.B(_12237_),
    .C(_12231_),
    .Y(_12239_),
    .A_N(_12238_));
 sg13g2_a221oi_1 _21204_ (.B2(_11440_),
    .C1(_12239_),
    .B1(net7670),
    .A1(net8006),
    .Y(_12240_),
    .A2(net7673));
 sg13g2_o21ai_1 _21205_ (.B1(net7998),
    .Y(_12241_),
    .A1(net8293),
    .A2(net8002));
 sg13g2_nor2_1 _21206_ (.A(net8381),
    .B(net8263),
    .Y(_12242_));
 sg13g2_a21oi_1 _21207_ (.A1(net8381),
    .A2(net8257),
    .Y(_12243_),
    .B1(_12242_));
 sg13g2_a22oi_1 _21208_ (.Y(_12244_),
    .B1(_12243_),
    .B2(net8293),
    .A2(_12241_),
    .A1(net8381));
 sg13g2_nand2_1 _21209_ (.Y(_12245_),
    .A(net7995),
    .B(_12190_));
 sg13g2_nor3_1 _21210_ (.A(net8442),
    .B(net7938),
    .C(_12181_),
    .Y(_12246_));
 sg13g2_nand2_1 _21211_ (.Y(_12247_),
    .A(net8252),
    .B(_12040_));
 sg13g2_o21ai_1 _21212_ (.B1(_12247_),
    .Y(_12248_),
    .A1(_11708_),
    .A2(_12035_));
 sg13g2_o21ai_1 _21213_ (.B1(_11705_),
    .Y(_12249_),
    .A1(_12246_),
    .A2(_12248_));
 sg13g2_o21ai_1 _21214_ (.B1(_12249_),
    .Y(_12250_),
    .A1(_11519_),
    .A2(net8004));
 sg13g2_nand3b_1 _21215_ (.B(_12245_),
    .C(_12244_),
    .Y(_12251_),
    .A_N(_12250_));
 sg13g2_a221oi_1 _21216_ (.B2(net8293),
    .C1(_12251_),
    .B1(net7670),
    .A1(net8381),
    .Y(_12252_),
    .A2(net7673));
 sg13g2_nand2_1 _21217_ (.Y(_12253_),
    .A(_11541_),
    .B(net8267));
 sg13g2_o21ai_1 _21218_ (.B1(net7936),
    .Y(_12254_),
    .A1(net8448),
    .A2(_11877_));
 sg13g2_a21oi_1 _21219_ (.A1(_11656_),
    .A2(_11863_),
    .Y(_12255_),
    .B1(_11660_));
 sg13g2_a221oi_1 _21220_ (.B2(net8252),
    .C1(_12255_),
    .B1(_11962_),
    .A1(net8248),
    .Y(_12256_),
    .A2(_11951_));
 sg13g2_o21ai_1 _21221_ (.B1(_11326_),
    .Y(_12257_),
    .A1(net8288),
    .A2(net8259));
 sg13g2_nor3_1 _21222_ (.A(net8288),
    .B(_11326_),
    .C(net8258),
    .Y(_12258_));
 sg13g2_nor2_1 _21223_ (.A(_11323_),
    .B(_11638_),
    .Y(_12259_));
 sg13g2_o21ai_1 _21224_ (.B1(net7999),
    .Y(_12260_),
    .A1(_12258_),
    .A2(_12259_));
 sg13g2_a21oi_1 _21225_ (.A1(_12257_),
    .A2(_12260_),
    .Y(_12261_),
    .B1(_12256_));
 sg13g2_nand3_1 _21226_ (.B(_12254_),
    .C(_12261_),
    .A(_12253_),
    .Y(_12262_));
 sg13g2_a221oi_1 _21227_ (.B2(_11323_),
    .C1(_12262_),
    .B1(net7670),
    .A1(_11327_),
    .Y(_12263_),
    .A2(net7674));
 sg13g2_o21ai_1 _21228_ (.B1(net7998),
    .Y(_12264_),
    .A1(_11268_),
    .A2(net8002));
 sg13g2_nand2_1 _21229_ (.Y(_12265_),
    .A(_11546_),
    .B(net8265));
 sg13g2_a22oi_1 _21230_ (.Y(_12266_),
    .B1(_11882_),
    .B2(net8252),
    .A2(_11871_),
    .A1(net8248));
 sg13g2_o21ai_1 _21231_ (.B1(_12266_),
    .Y(_12267_),
    .A1(net8443),
    .A2(_11941_));
 sg13g2_nand2_1 _21232_ (.Y(_12268_),
    .A(_11705_),
    .B(_12267_));
 sg13g2_a21oi_1 _21233_ (.A1(_11272_),
    .A2(net8257),
    .Y(_12269_),
    .B1(net8295));
 sg13g2_o21ai_1 _21234_ (.B1(_12269_),
    .Y(_12270_),
    .A1(_11272_),
    .A2(net8262));
 sg13g2_a22oi_1 _21235_ (.Y(_12271_),
    .B1(_12264_),
    .B2(_11272_),
    .A2(_11952_),
    .A1(net7995));
 sg13g2_nand4_1 _21236_ (.B(_12268_),
    .C(_12270_),
    .A(_12265_),
    .Y(_12272_),
    .D(_12271_));
 sg13g2_a221oi_1 _21237_ (.B2(_11268_),
    .C1(_12272_),
    .B1(net7670),
    .A1(_11272_),
    .Y(_12273_),
    .A2(net7673));
 sg13g2_nand2_1 _21238_ (.Y(_12274_),
    .A(net8443),
    .B(_11922_));
 sg13g2_nor2_1 _21239_ (.A(net8253),
    .B(_11930_),
    .Y(_12275_));
 sg13g2_o21ai_1 _21240_ (.B1(_12275_),
    .Y(_12276_),
    .A1(net8449),
    .A2(_12054_));
 sg13g2_a21oi_1 _21241_ (.A1(net8252),
    .A2(_12235_),
    .Y(_12277_),
    .B1(_11655_));
 sg13g2_o21ai_1 _21242_ (.B1(_10881_),
    .Y(_12278_),
    .A1(_11392_),
    .A2(net8260));
 sg13g2_nand2_1 _21243_ (.Y(_12279_),
    .A(net8379),
    .B(_12073_));
 sg13g2_o21ai_1 _21244_ (.B1(_12279_),
    .Y(_12280_),
    .A1(net8379),
    .A2(net8263));
 sg13g2_a22oi_1 _21245_ (.Y(_12281_),
    .B1(_12278_),
    .B2(net8379),
    .A2(_12274_),
    .A1(net7936));
 sg13g2_o21ai_1 _21246_ (.B1(_12281_),
    .Y(_12282_),
    .A1(net8281),
    .A2(_12280_));
 sg13g2_a221oi_1 _21247_ (.B2(_12277_),
    .C1(_12282_),
    .B1(_12276_),
    .A1(_11526_),
    .Y(_12283_),
    .A2(net8267));
 sg13g2_inv_1 _21248_ (.Y(_12284_),
    .A(_12283_));
 sg13g2_a221oi_1 _21249_ (.B2(_11392_),
    .C1(_12284_),
    .B1(net7671),
    .A1(net8379),
    .Y(_12285_),
    .A2(net7674));
 sg13g2_a21oi_1 _21250_ (.A1(_11625_),
    .A2(_11628_),
    .Y(_12286_),
    .B1(net8307));
 sg13g2_a21o_1 _21251_ (.A2(_11791_),
    .A1(net8428),
    .B1(_11873_),
    .X(_12287_));
 sg13g2_a21oi_2 _21252_ (.B1(net7938),
    .Y(_12288_),
    .A2(_12287_),
    .A1(net8432));
 sg13g2_o21ai_1 _21253_ (.B1(net7937),
    .Y(_12289_),
    .A1(net8450),
    .A2(_12288_));
 sg13g2_nor2b_1 _21254_ (.A(net8007),
    .B_N(net8307),
    .Y(_12290_));
 sg13g2_nor2b_1 _21255_ (.A(net8307),
    .B_N(net8007),
    .Y(_12291_));
 sg13g2_nor3_1 _21256_ (.A(net8259),
    .B(_12290_),
    .C(_12291_),
    .Y(_12292_));
 sg13g2_a221oi_1 _21257_ (.B2(_12291_),
    .C1(_12292_),
    .B1(_12074_),
    .A1(_10880_),
    .Y(_12293_),
    .A2(net8007));
 sg13g2_nor2_1 _21258_ (.A(net8409),
    .B(_12122_),
    .Y(_12294_));
 sg13g2_a21oi_2 _21259_ (.B1(_12294_),
    .Y(_12295_),
    .A2(_11828_),
    .A1(net8409));
 sg13g2_mux2_1 _21260_ (.A0(_12102_),
    .A1(_12124_),
    .S(net8413),
    .X(_12296_));
 sg13g2_nand2_1 _21261_ (.Y(_12297_),
    .A(net8436),
    .B(_12296_));
 sg13g2_o21ai_1 _21262_ (.B1(_12297_),
    .Y(_12298_),
    .A1(net8431),
    .A2(_12295_));
 sg13g2_nand2_1 _21263_ (.Y(_12299_),
    .A(net8447),
    .B(_12298_));
 sg13g2_a21oi_1 _21264_ (.A1(net8393),
    .A2(_12196_),
    .Y(_12300_),
    .B1(net8419));
 sg13g2_o21ai_1 _21265_ (.B1(_12300_),
    .Y(_12301_),
    .A1(net8393),
    .A2(_12191_));
 sg13g2_a21oi_1 _21266_ (.A1(net8417),
    .A2(_12113_),
    .Y(_12302_),
    .B1(net8251));
 sg13g2_nor2_1 _21267_ (.A(net8416),
    .B(_12117_),
    .Y(_12303_));
 sg13g2_a21oi_2 _21268_ (.B1(_12303_),
    .Y(_12304_),
    .A2(_12107_),
    .A1(net8415));
 sg13g2_a22oi_1 _21269_ (.Y(_12305_),
    .B1(_12304_),
    .B2(net8248),
    .A2(_12302_),
    .A1(_12301_));
 sg13g2_nand3_1 _21270_ (.B(_12299_),
    .C(_12305_),
    .A(_11654_),
    .Y(_12306_));
 sg13g2_nand3_1 _21271_ (.B(_12293_),
    .C(_12306_),
    .A(_12289_),
    .Y(_12307_));
 sg13g2_a21oi_1 _21272_ (.A1(_11540_),
    .A2(net8266),
    .Y(_12308_),
    .B1(_12307_));
 sg13g2_o21ai_1 _21273_ (.B1(net8007),
    .Y(_12309_),
    .A1(net7680),
    .A2(net7678));
 sg13g2_nand3b_1 _21274_ (.B(_12308_),
    .C(_12309_),
    .Y(_12310_),
    .A_N(_12286_));
 sg13g2_a21oi_1 _21275_ (.A1(net8442),
    .A2(_12038_),
    .Y(_12311_),
    .B1(_11940_));
 sg13g2_a21oi_1 _21276_ (.A1(_11656_),
    .A2(_12033_),
    .Y(_12312_),
    .B1(_11660_));
 sg13g2_a221oi_1 _21277_ (.B2(net8252),
    .C1(_12312_),
    .B1(_12205_),
    .A1(net8248),
    .Y(_12313_),
    .A2(_12189_));
 sg13g2_nand2_1 _21278_ (.Y(_12314_),
    .A(net8287),
    .B(net8264));
 sg13g2_nand3_1 _21279_ (.B(_11340_),
    .C(net8257),
    .A(net8287),
    .Y(_12315_));
 sg13g2_o21ai_1 _21280_ (.B1(_12315_),
    .Y(_12316_),
    .A1(net8287),
    .A2(_11638_));
 sg13g2_a22oi_1 _21281_ (.Y(_12317_),
    .B1(_12316_),
    .B2(net7998),
    .A2(_12314_),
    .A1(_11339_));
 sg13g2_nor3_1 _21282_ (.A(_12311_),
    .B(_12313_),
    .C(_12317_),
    .Y(_12318_));
 sg13g2_o21ai_1 _21283_ (.B1(_12318_),
    .Y(_12319_),
    .A1(_11537_),
    .A2(net8005));
 sg13g2_a221oi_1 _21284_ (.B2(net8287),
    .C1(_12319_),
    .B1(net7670),
    .A1(_11340_),
    .Y(_12320_),
    .A2(net7673));
 sg13g2_o21ai_1 _21285_ (.B1(net7996),
    .Y(_12321_),
    .A1(net8304),
    .A2(net8000));
 sg13g2_nor2_1 _21286_ (.A(net8520),
    .B(net8262),
    .Y(_12322_));
 sg13g2_a21oi_1 _21287_ (.A1(net8520),
    .A2(net8255),
    .Y(_12323_),
    .B1(_12322_));
 sg13g2_a22oi_1 _21288_ (.Y(_12324_),
    .B1(_12323_),
    .B2(net8304),
    .A2(_12321_),
    .A1(net8520));
 sg13g2_nand2_1 _21289_ (.Y(_12325_),
    .A(_11656_),
    .B(_12295_));
 sg13g2_nand2_1 _21290_ (.Y(_12326_),
    .A(_11864_),
    .B(_12295_));
 sg13g2_mux2_1 _21291_ (.A0(_11775_),
    .A1(_11784_),
    .S(net8416),
    .X(_12327_));
 sg13g2_nand2_1 _21292_ (.Y(_12328_),
    .A(net8434),
    .B(_12327_));
 sg13g2_o21ai_1 _21293_ (.B1(_12328_),
    .Y(_12329_),
    .A1(net8432),
    .A2(_12287_));
 sg13g2_nand2_1 _21294_ (.Y(_12330_),
    .A(net8447),
    .B(_12329_));
 sg13g2_nor2_1 _21295_ (.A(net8413),
    .B(_11822_),
    .Y(_12331_));
 sg13g2_a21oi_1 _21296_ (.A1(net8413),
    .A2(_11768_),
    .Y(_12332_),
    .B1(_12331_));
 sg13g2_mux2_1 _21297_ (.A0(_11807_),
    .A1(_11814_),
    .S(net8411),
    .X(_12333_));
 sg13g2_a22oi_1 _21298_ (.Y(_12334_),
    .B1(_12333_),
    .B2(net8253),
    .A2(_12332_),
    .A1(net8245));
 sg13g2_nand2_1 _21299_ (.Y(_12335_),
    .A(_12330_),
    .B(_12334_));
 sg13g2_a22oi_1 _21300_ (.Y(_12336_),
    .B1(_11705_),
    .B2(_12335_),
    .A2(net8265),
    .A1(_11565_));
 sg13g2_nand3_1 _21301_ (.B(_12326_),
    .C(_12336_),
    .A(_12324_),
    .Y(_12337_));
 sg13g2_a221oi_1 _21302_ (.B2(net8306),
    .C1(_12337_),
    .B1(net7671),
    .A1(net8520),
    .Y(_12338_),
    .A2(net7672));
 sg13g2_nand2_1 _21303_ (.Y(_12339_),
    .A(_11580_),
    .B(net8266));
 sg13g2_o21ai_1 _21304_ (.B1(net7937),
    .Y(_12340_),
    .A1(net8450),
    .A2(_11794_));
 sg13g2_o21ai_1 _21305_ (.B1(net7998),
    .Y(_12341_),
    .A1(net8276),
    .A2(net8002));
 sg13g2_o21ai_1 _21306_ (.B1(net8276),
    .Y(_12342_),
    .A1(_11416_),
    .A2(net8258));
 sg13g2_nand2_1 _21307_ (.Y(_12343_),
    .A(_11417_),
    .B(_12341_));
 sg13g2_a22oi_1 _21308_ (.Y(_12344_),
    .B1(_12342_),
    .B2(_12343_),
    .A2(net8259),
    .A1(_11416_));
 sg13g2_nand2_1 _21309_ (.Y(_12345_),
    .A(net7994),
    .B(_11830_));
 sg13g2_a22oi_1 _21310_ (.Y(_12346_),
    .B1(_12126_),
    .B2(net8247),
    .A2(_12108_),
    .A1(net8252));
 sg13g2_a21oi_1 _21311_ (.A1(_12345_),
    .A2(_12346_),
    .Y(_12347_),
    .B1(_12344_));
 sg13g2_nand3_1 _21312_ (.B(_12340_),
    .C(_12347_),
    .A(_12339_),
    .Y(_12348_));
 sg13g2_a221oi_1 _21313_ (.B2(net8276),
    .C1(_12348_),
    .B1(net7671),
    .A1(_11417_),
    .Y(_12349_),
    .A2(net7673));
 sg13g2_o21ai_1 _21314_ (.B1(net8505),
    .Y(_12350_),
    .A1(net7679),
    .A2(net7677));
 sg13g2_nor2_1 _21315_ (.A(net8444),
    .B(_12098_),
    .Y(_12351_));
 sg13g2_a221oi_1 _21316_ (.B2(net8253),
    .C1(_12351_),
    .B1(_11824_),
    .A1(net8246),
    .Y(_12352_),
    .A2(_11777_));
 sg13g2_a21oi_1 _21317_ (.A1(net8505),
    .A2(net8255),
    .Y(_12353_),
    .B1(_11246_));
 sg13g2_o21ai_1 _21318_ (.B1(net7996),
    .Y(_12354_),
    .A1(_11247_),
    .A2(net8000));
 sg13g2_a21o_1 _21319_ (.A2(_12354_),
    .A1(net8505),
    .B1(_12353_),
    .X(_12355_));
 sg13g2_o21ai_1 _21320_ (.B1(_12355_),
    .Y(_12356_),
    .A1(net8505),
    .A2(net8262));
 sg13g2_o21ai_1 _21321_ (.B1(_12356_),
    .Y(_12357_),
    .A1(net8249),
    .A2(_12352_));
 sg13g2_a221oi_1 _21322_ (.B2(_12129_),
    .C1(_12357_),
    .B1(net7995),
    .A1(_11557_),
    .Y(_12358_),
    .A2(net8265));
 sg13g2_o21ai_1 _21323_ (.B1(_11247_),
    .Y(_12359_),
    .A1(net7676),
    .A2(net7675));
 sg13g2_nand3_1 _21324_ (.B(_12358_),
    .C(_12359_),
    .A(_12350_),
    .Y(_12360_));
 sg13g2_o21ai_1 _21325_ (.B1(net7996),
    .Y(_12361_),
    .A1(net8301),
    .A2(net8001));
 sg13g2_nand2_1 _21326_ (.Y(_12362_),
    .A(_11569_),
    .B(net8265));
 sg13g2_nand2_1 _21327_ (.Y(_12363_),
    .A(net8434),
    .B(_11995_));
 sg13g2_o21ai_1 _21328_ (.B1(_12363_),
    .Y(_12364_),
    .A1(net8433),
    .A2(_11988_));
 sg13g2_nand2_1 _21329_ (.Y(_12365_),
    .A(net8412),
    .B(_12042_));
 sg13g2_nand2_1 _21330_ (.Y(_12366_),
    .A(net8401),
    .B(_11803_));
 sg13g2_a21oi_1 _21331_ (.A1(net8389),
    .A2(_11797_),
    .Y(_12367_),
    .B1(net8411));
 sg13g2_a21oi_1 _21332_ (.A1(_12366_),
    .A2(_12367_),
    .Y(_12368_),
    .B1(net8251));
 sg13g2_a221oi_1 _21333_ (.B2(_12368_),
    .C1(net8249),
    .B1(_12365_),
    .A1(net8245),
    .Y(_12369_),
    .A2(_12000_));
 sg13g2_o21ai_1 _21334_ (.B1(_12369_),
    .Y(_12370_),
    .A1(net8446),
    .A2(_12364_));
 sg13g2_nor3_1 _21335_ (.A(net8449),
    .B(_11657_),
    .C(_12006_),
    .Y(_12371_));
 sg13g2_nor2_1 _21336_ (.A(net8438),
    .B(net8262),
    .Y(_12372_));
 sg13g2_a21oi_1 _21337_ (.A1(net8438),
    .A2(net8255),
    .Y(_12373_),
    .B1(_12372_));
 sg13g2_a221oi_1 _21338_ (.B2(net8301),
    .C1(_12371_),
    .B1(_12373_),
    .A1(net8438),
    .Y(_12374_),
    .A2(_12361_));
 sg13g2_nand3_1 _21339_ (.B(_12370_),
    .C(_12374_),
    .A(_12362_),
    .Y(_12375_));
 sg13g2_a221oi_1 _21340_ (.B2(net8302),
    .C1(_12375_),
    .B1(net7669),
    .A1(net8438),
    .Y(_12376_),
    .A2(net7672));
 sg13g2_nand2b_2 _21341_ (.Y(_12377_),
    .B(_12376_),
    .A_N(_12360_));
 sg13g2_a21o_1 _21342_ (.A2(_11532_),
    .A1(_11531_),
    .B1(net8005),
    .X(_12378_));
 sg13g2_o21ai_1 _21343_ (.B1(net7937),
    .Y(_12379_),
    .A1(net8448),
    .A2(_12364_));
 sg13g2_o21ai_1 _21344_ (.B1(_11661_),
    .Y(_12380_),
    .A1(_11657_),
    .A2(_12006_));
 sg13g2_nor2_1 _21345_ (.A(_11708_),
    .B(_12016_),
    .Y(_12381_));
 sg13g2_a21o_1 _21346_ (.A2(net8264),
    .A1(net8279),
    .B1(_11404_),
    .X(_12382_));
 sg13g2_o21ai_1 _21347_ (.B1(net7998),
    .Y(_12383_),
    .A1(net8279),
    .A2(net8002));
 sg13g2_a21oi_1 _21348_ (.A1(_11404_),
    .A2(net8257),
    .Y(_12384_),
    .B1(_11402_));
 sg13g2_o21ai_1 _21349_ (.B1(_12382_),
    .Y(_12385_),
    .A1(_12383_),
    .A2(_12384_));
 sg13g2_o21ai_1 _21350_ (.B1(_12380_),
    .Y(_12386_),
    .A1(net8251),
    .A2(_12220_));
 sg13g2_o21ai_1 _21351_ (.B1(_12379_),
    .Y(_12387_),
    .A1(_12381_),
    .A2(_12386_));
 sg13g2_nand3b_1 _21352_ (.B(_12385_),
    .C(_12378_),
    .Y(_12388_),
    .A_N(_12387_));
 sg13g2_a221oi_1 _21353_ (.B2(net8280),
    .C1(_12388_),
    .B1(net7670),
    .A1(_11404_),
    .Y(_12389_),
    .A2(net7673));
 sg13g2_nand2b_1 _21354_ (.Y(_12390_),
    .B(net8442),
    .A_N(_12329_));
 sg13g2_nand2_1 _21355_ (.Y(_12391_),
    .A(net7994),
    .B(_12325_));
 sg13g2_a22oi_1 _21356_ (.Y(_12392_),
    .B1(_12304_),
    .B2(net8254),
    .A2(_12296_),
    .A1(net8248));
 sg13g2_o21ai_1 _21357_ (.B1(net7998),
    .Y(_12393_),
    .A1(net8284),
    .A2(net8002));
 sg13g2_nand2_1 _21358_ (.Y(_12394_),
    .A(_11365_),
    .B(_12393_));
 sg13g2_o21ai_1 _21359_ (.B1(net8284),
    .Y(_12395_),
    .A1(_11366_),
    .A2(net8258));
 sg13g2_a22oi_1 _21360_ (.Y(_12396_),
    .B1(_12394_),
    .B2(_12395_),
    .A2(net8259),
    .A1(_11366_));
 sg13g2_a221oi_1 _21361_ (.B2(_12392_),
    .C1(_12396_),
    .B1(_12391_),
    .A1(net7936),
    .Y(_12397_),
    .A2(_12390_));
 sg13g2_o21ai_1 _21362_ (.B1(_12397_),
    .Y(_12398_),
    .A1(_11530_),
    .A2(net8005));
 sg13g2_a221oi_1 _21363_ (.B2(net8284),
    .C1(_12398_),
    .B1(net7670),
    .A1(_11365_),
    .Y(_12399_),
    .A2(net7674));
 sg13g2_o21ai_1 _21364_ (.B1(net7997),
    .Y(_12400_),
    .A1(_11118_),
    .A2(net8000));
 sg13g2_o21ai_1 _21365_ (.B1(_11118_),
    .Y(_12401_),
    .A1(net7676),
    .A2(net7675));
 sg13g2_nor2_1 _21366_ (.A(_11567_),
    .B(net8004),
    .Y(_12402_));
 sg13g2_nand2b_1 _21367_ (.Y(_12403_),
    .B(net8448),
    .A_N(_12166_));
 sg13g2_nor2_1 _21368_ (.A(net8420),
    .B(_11720_),
    .Y(_12404_));
 sg13g2_a21oi_2 _21369_ (.B1(_12404_),
    .Y(_12405_),
    .A2(_11667_),
    .A1(net8420));
 sg13g2_nand2_1 _21370_ (.Y(_12406_),
    .A(net8420),
    .B(_11714_));
 sg13g2_a21oi_1 _21371_ (.A1(net8427),
    .A2(_11699_),
    .Y(_12407_),
    .B1(net8251));
 sg13g2_a22oi_1 _21372_ (.Y(_12408_),
    .B1(_12406_),
    .B2(_12407_),
    .A2(_12405_),
    .A1(net8245));
 sg13g2_a21oi_2 _21373_ (.B1(net8250),
    .Y(_12409_),
    .A2(_12408_),
    .A1(_12403_));
 sg13g2_a21oi_1 _21374_ (.A1(net8446),
    .A2(net8261),
    .Y(_12410_),
    .B1(net8303));
 sg13g2_o21ai_1 _21375_ (.B1(net8450),
    .Y(_12411_),
    .A1(net7679),
    .A2(net7677));
 sg13g2_nand2_1 _21376_ (.Y(_12412_),
    .A(net8449),
    .B(net8255));
 sg13g2_a22oi_1 _21377_ (.Y(_12413_),
    .B1(_12410_),
    .B2(_12412_),
    .A2(_12400_),
    .A1(net8449));
 sg13g2_o21ai_1 _21378_ (.B1(_12413_),
    .Y(_12414_),
    .A1(_11865_),
    .A2(_12141_));
 sg13g2_nor3_2 _21379_ (.A(_12402_),
    .B(_12409_),
    .C(_12414_),
    .Y(_12415_));
 sg13g2_and3_2 _21380_ (.X(_12416_),
    .A(_12401_),
    .B(_12411_),
    .C(_12415_));
 sg13g2_nand3_1 _21381_ (.B(_12411_),
    .C(_12415_),
    .A(_12401_),
    .Y(_12417_));
 sg13g2_nand2_1 _21382_ (.Y(_12418_),
    .A(_11547_),
    .B(net8265));
 sg13g2_a21oi_1 _21383_ (.A1(net8442),
    .A2(_11689_),
    .Y(_12419_),
    .B1(_11940_));
 sg13g2_o21ai_1 _21384_ (.B1(net7998),
    .Y(_12420_),
    .A1(_11379_),
    .A2(net8002));
 sg13g2_nor2_1 _21385_ (.A(_11383_),
    .B(net8258),
    .Y(_12421_));
 sg13g2_a21oi_1 _21386_ (.A1(_11383_),
    .A2(net8259),
    .Y(_12422_),
    .B1(_12421_));
 sg13g2_a221oi_1 _21387_ (.B2(_11379_),
    .C1(_12419_),
    .B1(_12422_),
    .A1(_11382_),
    .Y(_12423_),
    .A2(_12420_));
 sg13g2_a22oi_1 _21388_ (.Y(_12424_),
    .B1(net8247),
    .B2(_11905_),
    .A2(_11661_),
    .A1(_11658_));
 sg13g2_o21ai_1 _21389_ (.B1(_12424_),
    .Y(_12425_),
    .A1(net8251),
    .A2(_12084_));
 sg13g2_nand3_1 _21390_ (.B(_12423_),
    .C(_12425_),
    .A(_12418_),
    .Y(_12426_));
 sg13g2_a221oi_1 _21391_ (.B2(_11379_),
    .C1(_12426_),
    .B1(net7670),
    .A1(_11382_),
    .Y(_12427_),
    .A2(net7673));
 sg13g2_o21ai_1 _21392_ (.B1(net7997),
    .Y(_12428_),
    .A1(net8292),
    .A2(net8001));
 sg13g2_nor2_1 _21393_ (.A(net8380),
    .B(net8262),
    .Y(_12429_));
 sg13g2_a21oi_1 _21394_ (.A1(net8380),
    .A2(net8256),
    .Y(_12430_),
    .B1(_12429_));
 sg13g2_a22oi_1 _21395_ (.Y(_12431_),
    .B1(_12430_),
    .B2(net8292),
    .A2(_12428_),
    .A1(net8380));
 sg13g2_o21ai_1 _21396_ (.B1(_12431_),
    .Y(_12432_),
    .A1(net7994),
    .A2(_12145_));
 sg13g2_nand2_1 _21397_ (.Y(_12433_),
    .A(net8447),
    .B(_12156_));
 sg13g2_a22oi_1 _21398_ (.Y(_12434_),
    .B1(_12405_),
    .B2(net8252),
    .A2(_12164_),
    .A1(net8245));
 sg13g2_a21oi_1 _21399_ (.A1(_12433_),
    .A2(_12434_),
    .Y(_12435_),
    .B1(net8250));
 sg13g2_nor2_1 _21400_ (.A(_12432_),
    .B(_12435_),
    .Y(_12436_));
 sg13g2_o21ai_1 _21401_ (.B1(_12436_),
    .Y(_12437_),
    .A1(_11555_),
    .A2(net8004));
 sg13g2_a221oi_1 _21402_ (.B2(net8292),
    .C1(_12437_),
    .B1(net7669),
    .A1(net8380),
    .Y(_12438_),
    .A2(net7672));
 sg13g2_nand2_1 _21403_ (.Y(_12439_),
    .A(net8291),
    .B(_11638_));
 sg13g2_nand2_1 _21404_ (.Y(_12440_),
    .A(net8447),
    .B(_12288_));
 sg13g2_a22oi_1 _21405_ (.Y(_12441_),
    .B1(_12332_),
    .B2(net8252),
    .A2(_12327_),
    .A1(net8246));
 sg13g2_a21oi_1 _21406_ (.A1(_12440_),
    .A2(_12441_),
    .Y(_12442_),
    .B1(net8249));
 sg13g2_nor2_1 _21407_ (.A(net7994),
    .B(_12298_),
    .Y(_12443_));
 sg13g2_nand2_1 _21408_ (.Y(_12444_),
    .A(net8290),
    .B(net8261));
 sg13g2_o21ai_1 _21409_ (.B1(_12444_),
    .Y(_12445_),
    .A1(net8290),
    .A2(net8258));
 sg13g2_nor2_1 _21410_ (.A(net8291),
    .B(_12445_),
    .Y(_12446_));
 sg13g2_a21oi_1 _21411_ (.A1(net7997),
    .A2(_12439_),
    .Y(_12447_),
    .B1(net8290));
 sg13g2_nor4_1 _21412_ (.A(_12442_),
    .B(_12443_),
    .C(_12446_),
    .D(_12447_),
    .Y(_12448_));
 sg13g2_o21ai_1 _21413_ (.B1(_12448_),
    .Y(_12449_),
    .A1(_11553_),
    .A2(net8004));
 sg13g2_a221oi_1 _21414_ (.B2(_11304_),
    .C1(_12449_),
    .B1(net7669),
    .A1(_11308_),
    .Y(_12450_),
    .A2(net7674));
 sg13g2_inv_1 _21415_ (.Y(_12451_),
    .A(_12450_));
 sg13g2_nand4_1 _21416_ (.B(_12240_),
    .C(_12338_),
    .A(_11893_),
    .Y(_12452_),
    .D(_12416_));
 sg13g2_nand4_1 _21417_ (.B(_12252_),
    .C(_12273_),
    .A(_12051_),
    .Y(_12453_),
    .D(_12438_));
 sg13g2_nand2_1 _21418_ (.Y(_12454_),
    .A(_11936_),
    .B(_12179_));
 sg13g2_or4_1 _21419_ (.A(_11982_),
    .B(_12095_),
    .C(_12136_),
    .D(_12225_),
    .X(_12455_));
 sg13g2_or3_1 _21420_ (.A(_12162_),
    .B(_12210_),
    .C(_12310_),
    .X(_12456_));
 sg13g2_nor4_1 _21421_ (.A(_12452_),
    .B(_12453_),
    .C(_12455_),
    .D(_12456_),
    .Y(_12457_));
 sg13g2_nor4_2 _21422_ (.A(_11914_),
    .B(_12026_),
    .C(_12069_),
    .Y(_12458_),
    .D(_12451_));
 sg13g2_nand4_1 _21423_ (.B(_12285_),
    .C(_12349_),
    .A(_11837_),
    .Y(_12459_),
    .D(_12389_));
 sg13g2_nand4_1 _21424_ (.B(_12320_),
    .C(_12399_),
    .A(_12263_),
    .Y(_12460_),
    .D(_12427_));
 sg13g2_nor4_1 _21425_ (.A(_12377_),
    .B(_12454_),
    .C(_12459_),
    .D(_12460_),
    .Y(_12461_));
 sg13g2_nand4_1 _21426_ (.B(_12457_),
    .C(_12458_),
    .A(_11729_),
    .Y(_12462_),
    .D(_12461_));
 sg13g2_nand2_1 _21427_ (.Y(_12463_),
    .A(net8837),
    .B(_11751_));
 sg13g2_nor3_1 _21428_ (.A(_11732_),
    .B(net8697),
    .C(_12463_),
    .Y(_12464_));
 sg13g2_o21ai_1 _21429_ (.B1(_12464_),
    .Y(_12465_),
    .A1(_10836_),
    .A2(_11753_));
 sg13g2_nor3_1 _21430_ (.A(net8577),
    .B(_10867_),
    .C(_12465_),
    .Y(_12466_));
 sg13g2_o21ai_1 _21431_ (.B1(_12466_),
    .Y(_12467_),
    .A1(_10877_),
    .A2(_12462_));
 sg13g2_inv_2 _21432_ (.Y(_12468_),
    .A(net7480));
 sg13g2_nand2b_2 _21433_ (.Y(_12469_),
    .B(net7480),
    .A_N(net9271));
 sg13g2_a21o_1 _21434_ (.A2(net8704),
    .A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[27] ),
    .B1(net8699),
    .X(_12470_));
 sg13g2_a21oi_1 _21435_ (.A1(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[27] ),
    .A2(net8839),
    .Y(_12471_),
    .B1(_12470_));
 sg13g2_o21ai_1 _21436_ (.B1(net8660),
    .Y(_12472_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[27] ),
    .A2(net8692));
 sg13g2_o21ai_1 _21437_ (.B1(net8634),
    .Y(_12473_),
    .A1(_12471_),
    .A2(_12472_));
 sg13g2_a21o_1 _21438_ (.A2(_12225_),
    .A1(_10869_),
    .B1(_12473_),
    .X(_12474_));
 sg13g2_a21oi_1 _21439_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[27] ),
    .A2(net8738),
    .Y(_12475_),
    .B1(net8628));
 sg13g2_nor2_2 _21440_ (.A(net8500),
    .B(_12475_),
    .Y(_12476_));
 sg13g2_a22oi_1 _21441_ (.Y(_12477_),
    .B1(_12474_),
    .B2(_12476_),
    .A2(net8375),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[27] ));
 sg13g2_nand2_1 _21442_ (.Y(_12478_),
    .A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[26] ),
    .B(net8839));
 sg13g2_a21oi_1 _21443_ (.A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[26] ),
    .A2(net8705),
    .Y(_12479_),
    .B1(net8700));
 sg13g2_o21ai_1 _21444_ (.B1(net8662),
    .Y(_12480_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[26] ),
    .A2(net8690));
 sg13g2_a21oi_1 _21445_ (.A1(_12478_),
    .A2(_12479_),
    .Y(_12481_),
    .B1(_12480_));
 sg13g2_nor2_1 _21446_ (.A(net8707),
    .B(_12481_),
    .Y(_12482_));
 sg13g2_o21ai_1 _21447_ (.B1(_12482_),
    .Y(_12483_),
    .A1(net8662),
    .A2(_12240_));
 sg13g2_a21oi_1 _21448_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[26] ),
    .A2(net8736),
    .Y(_12484_),
    .B1(net8632));
 sg13g2_nor2_1 _21449_ (.A(net8503),
    .B(_12484_),
    .Y(_12485_));
 sg13g2_a22oi_1 _21450_ (.Y(_12486_),
    .B1(_12483_),
    .B2(_12485_),
    .A2(net8378),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[26] ));
 sg13g2_a221oi_1 _21451_ (.B2(_12476_),
    .C1(_10858_),
    .B1(_12474_),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[27] ),
    .Y(_12487_),
    .A2(net8375));
 sg13g2_nor2_1 _21452_ (.A(\soc_I.PC[27] ),
    .B(\soc_I.PC[26] ),
    .Y(_12488_));
 sg13g2_a22oi_1 _21453_ (.Y(_12489_),
    .B1(_12488_),
    .B2(_10858_),
    .A2(_12487_),
    .A1(_12486_));
 sg13g2_a21o_1 _21454_ (.A2(net8705),
    .A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[25] ),
    .B1(net8700),
    .X(_12490_));
 sg13g2_a21oi_1 _21455_ (.A1(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[25] ),
    .A2(net8840),
    .Y(_12491_),
    .B1(_12490_));
 sg13g2_o21ai_1 _21456_ (.B1(net8661),
    .Y(_12492_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[25] ),
    .A2(net8694));
 sg13g2_o21ai_1 _21457_ (.B1(net8632),
    .Y(_12493_),
    .A1(_12491_),
    .A2(_12492_));
 sg13g2_a21o_1 _21458_ (.A2(_12136_),
    .A1(net8655),
    .B1(_12493_),
    .X(_12494_));
 sg13g2_a21oi_1 _21459_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[25] ),
    .A2(net8736),
    .Y(_12495_),
    .B1(net8633));
 sg13g2_nor2_1 _21460_ (.A(net8503),
    .B(_12495_),
    .Y(_12496_));
 sg13g2_a22oi_1 _21461_ (.Y(_12497_),
    .B1(_12494_),
    .B2(_12496_),
    .A2(net8377),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[25] ));
 sg13g2_nor2_1 _21462_ (.A(\soc_I.PC[25] ),
    .B(net8577),
    .Y(_12498_));
 sg13g2_a21oi_2 _21463_ (.B1(_12498_),
    .Y(_12499_),
    .A2(_12497_),
    .A1(net8577));
 sg13g2_or2_2 _21464_ (.X(_12500_),
    .B(_12499_),
    .A(_12489_));
 sg13g2_nor2_2 _21465_ (.A(\soc_I.PC[24] ),
    .B(net8570),
    .Y(_12501_));
 sg13g2_a21o_1 _21466_ (.A2(net8704),
    .A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[24] ),
    .B1(net8699),
    .X(_12502_));
 sg13g2_a21oi_1 _21467_ (.A1(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[24] ),
    .A2(net8839),
    .Y(_12503_),
    .B1(_12502_));
 sg13g2_o21ai_1 _21468_ (.B1(net8661),
    .Y(_12504_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[24] ),
    .A2(net8693));
 sg13g2_o21ai_1 _21469_ (.B1(net8632),
    .Y(_12505_),
    .A1(_12503_),
    .A2(_12504_));
 sg13g2_a21o_1 _21470_ (.A2(_12095_),
    .A1(net8655),
    .B1(_12505_),
    .X(_12506_));
 sg13g2_a21oi_1 _21471_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[24] ),
    .A2(net8736),
    .Y(_12507_),
    .B1(net8632));
 sg13g2_nor2_1 _21472_ (.A(net8503),
    .B(_12507_),
    .Y(_12508_));
 sg13g2_a22oi_1 _21473_ (.Y(_12509_),
    .B1(_12506_),
    .B2(_12508_),
    .A2(net8377),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[24] ));
 sg13g2_a21oi_2 _21474_ (.B1(_12501_),
    .Y(_12510_),
    .A2(net7647),
    .A1(net8571));
 sg13g2_a21o_1 _21475_ (.A2(net7647),
    .A1(net8571),
    .B1(_12501_),
    .X(_12511_));
 sg13g2_a21o_1 _21476_ (.A2(net8704),
    .A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[28] ),
    .B1(net8699),
    .X(_12512_));
 sg13g2_a21oi_1 _21477_ (.A1(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[28] ),
    .A2(net8839),
    .Y(_12513_),
    .B1(_12512_));
 sg13g2_o21ai_1 _21478_ (.B1(net8660),
    .Y(_12514_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[28] ),
    .A2(net8692));
 sg13g2_o21ai_1 _21479_ (.B1(net8632),
    .Y(_12515_),
    .A1(_12513_),
    .A2(_12514_));
 sg13g2_a21o_1 _21480_ (.A2(_12162_),
    .A1(_10869_),
    .B1(_12515_),
    .X(_12516_));
 sg13g2_a21oi_1 _21481_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[28] ),
    .A2(net8736),
    .Y(_12517_),
    .B1(net8632));
 sg13g2_nor2_1 _21482_ (.A(net8504),
    .B(_12517_),
    .Y(_12518_));
 sg13g2_a22oi_1 _21483_ (.Y(_12519_),
    .B1(_12516_),
    .B2(_12518_),
    .A2(net8377),
    .A1(net2683));
 sg13g2_nor2_1 _21484_ (.A(\soc_I.PC[28] ),
    .B(net8575),
    .Y(_12520_));
 sg13g2_a21oi_2 _21485_ (.B1(_12520_),
    .Y(_12521_),
    .A2(net7641),
    .A1(net8575));
 sg13g2_or3_1 _21486_ (.A(_12500_),
    .B(_12510_),
    .C(_12521_),
    .X(_12522_));
 sg13g2_a21o_1 _21487_ (.A2(net8701),
    .A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[31] ),
    .B1(net8696),
    .X(_12523_));
 sg13g2_a21oi_1 _21488_ (.A1(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[31] ),
    .A2(net8836),
    .Y(_12524_),
    .B1(_12523_));
 sg13g2_o21ai_1 _21489_ (.B1(net8660),
    .Y(_12525_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[31] ),
    .A2(net8692));
 sg13g2_o21ai_1 _21490_ (.B1(net8628),
    .Y(_12526_),
    .A1(_12524_),
    .A2(_12525_));
 sg13g2_a21o_1 _21491_ (.A2(_12210_),
    .A1(net8655),
    .B1(_12526_),
    .X(_12527_));
 sg13g2_a21oi_1 _21492_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[31] ),
    .A2(net8730),
    .Y(_12528_),
    .B1(net8627));
 sg13g2_nor2_1 _21493_ (.A(net8499),
    .B(_12528_),
    .Y(_12529_));
 sg13g2_a22oi_1 _21494_ (.Y(_12530_),
    .B1(_12527_),
    .B2(_12529_),
    .A2(net8374),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[31] ));
 sg13g2_mux2_2 _21495_ (.A0(_10450_),
    .A1(_12530_),
    .S(net8570),
    .X(_12531_));
 sg13g2_o21ai_1 _21496_ (.B1(net8660),
    .Y(_12532_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[29] ),
    .A2(net8692));
 sg13g2_a21o_1 _21497_ (.A2(net8704),
    .A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[29] ),
    .B1(net8699),
    .X(_12533_));
 sg13g2_a21oi_1 _21498_ (.A1(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[29] ),
    .A2(net8839),
    .Y(_12534_),
    .B1(_12533_));
 sg13g2_o21ai_1 _21499_ (.B1(net8632),
    .Y(_12535_),
    .A1(_12532_),
    .A2(_12534_));
 sg13g2_a21o_1 _21500_ (.A2(_12310_),
    .A1(net8655),
    .B1(_12535_),
    .X(_12536_));
 sg13g2_a21oi_1 _21501_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[29] ),
    .A2(net8736),
    .Y(_12537_),
    .B1(net8632));
 sg13g2_nor2_1 _21502_ (.A(net8503),
    .B(_12537_),
    .Y(_12538_));
 sg13g2_a22oi_1 _21503_ (.Y(_12539_),
    .B1(_12536_),
    .B2(_12538_),
    .A2(net8377),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[29] ));
 sg13g2_mux2_2 _21504_ (.A0(_10452_),
    .A1(_12539_),
    .S(net8575),
    .X(_12540_));
 sg13g2_a21o_1 _21505_ (.A2(net8701),
    .A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[30] ),
    .B1(net8696),
    .X(_12541_));
 sg13g2_a21oi_1 _21506_ (.A1(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[30] ),
    .A2(net8837),
    .Y(_12542_),
    .B1(_12541_));
 sg13g2_o21ai_1 _21507_ (.B1(net8662),
    .Y(_12543_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[30] ),
    .A2(net8690));
 sg13g2_o21ai_1 _21508_ (.B1(net8628),
    .Y(_12544_),
    .A1(_12542_),
    .A2(_12543_));
 sg13g2_a21o_1 _21509_ (.A2(_11982_),
    .A1(net8655),
    .B1(_12544_),
    .X(_12545_));
 sg13g2_a21oi_1 _21510_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[30] ),
    .A2(net8730),
    .Y(_12546_),
    .B1(net8627));
 sg13g2_nor2_1 _21511_ (.A(net8499),
    .B(_12546_),
    .Y(_12547_));
 sg13g2_a22oi_1 _21512_ (.Y(_12548_),
    .B1(_12545_),
    .B2(_12547_),
    .A2(net8374),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[30] ));
 sg13g2_mux2_2 _21513_ (.A0(_10451_),
    .A1(net7624),
    .S(net8578),
    .X(_12549_));
 sg13g2_nand3b_1 _21514_ (.B(_12540_),
    .C(_12549_),
    .Y(_12550_),
    .A_N(_12522_));
 sg13g2_nand3_1 _21515_ (.B(_12531_),
    .C(_12549_),
    .A(_10856_),
    .Y(_12551_));
 sg13g2_or2_1 _21516_ (.X(_12552_),
    .B(_12551_),
    .A(_12540_));
 sg13g2_nor3_1 _21517_ (.A(_12469_),
    .B(_12522_),
    .C(_12552_),
    .Y(_12553_));
 sg13g2_nor3_2 _21518_ (.A(_12469_),
    .B(_12531_),
    .C(_12550_),
    .Y(_12554_));
 sg13g2_or3_1 _21519_ (.A(_12469_),
    .B(_12531_),
    .C(_12550_),
    .X(_12555_));
 sg13g2_nand2b_1 _21520_ (.Y(_12556_),
    .B(net7458),
    .A_N(_12553_));
 sg13g2_and2_1 _21521_ (.A(_00244_),
    .B(_12556_),
    .X(_12557_));
 sg13g2_inv_1 _21522_ (.Y(_12558_),
    .A(_12557_));
 sg13g2_nand2_1 _21523_ (.Y(_12559_),
    .A(net8683),
    .B(_12557_));
 sg13g2_nor2_2 _21524_ (.A(net9020),
    .B(net8677),
    .Y(_12560_));
 sg13g2_and2_1 _21525_ (.A(\soc_I.qqspi_I.state[3] ),
    .B(net8626),
    .X(_12561_));
 sg13g2_nand2_2 _21526_ (.Y(_12562_),
    .A(net4673),
    .B(net8626));
 sg13g2_a21oi_1 _21527_ (.A1(net5067),
    .A2(_12559_),
    .Y(_12563_),
    .B1(net9297));
 sg13g2_nand2_1 _21528_ (.Y(_00004_),
    .A(net8555),
    .B(_12563_));
 sg13g2_nor2_2 _21529_ (.A(net9297),
    .B(net8685),
    .Y(_12564_));
 sg13g2_nand2_1 _21530_ (.Y(_12565_),
    .A(net4977),
    .B(_12564_));
 sg13g2_nand3_1 _21531_ (.B(net9001),
    .C(net8683),
    .A(net4574),
    .Y(_12566_));
 sg13g2_o21ai_1 _21532_ (.B1(_12565_),
    .Y(_00005_),
    .A1(net8665),
    .A2(_12566_));
 sg13g2_a22oi_1 _21533_ (.Y(_12567_),
    .B1(_12564_),
    .B2(net4069),
    .A2(net8626),
    .A1(net3104));
 sg13g2_inv_1 _21534_ (.Y(_00006_),
    .A(net4070));
 sg13g2_a22oi_1 _21535_ (.Y(_12568_),
    .B1(_12564_),
    .B2(net4673),
    .A2(net8626),
    .A1(net9195));
 sg13g2_inv_1 _21536_ (.Y(_00007_),
    .A(net4674));
 sg13g2_nand2_1 _21537_ (.Y(_12569_),
    .A(net3104),
    .B(_12564_));
 sg13g2_nand2_1 _21538_ (.Y(_12570_),
    .A(\soc_I.qqspi_I.state[0] ),
    .B(net9001));
 sg13g2_o21ai_1 _21539_ (.B1(net3105),
    .Y(_00008_),
    .A1(_12559_),
    .A2(_12570_));
 sg13g2_a22oi_1 _21540_ (.Y(_12571_),
    .B1(_12564_),
    .B2(net9195),
    .A2(net8626),
    .A1(net4977));
 sg13g2_o21ai_1 _21541_ (.B1(net4978),
    .Y(_00009_),
    .A1(_10856_),
    .A2(_12566_));
 sg13g2_a22oi_1 _21542_ (.Y(_12572_),
    .B1(_12564_),
    .B2(net4574),
    .A2(net8626),
    .A1(net4069));
 sg13g2_inv_1 _21543_ (.Y(_00010_),
    .A(net4575));
 sg13g2_nand2_2 _21544_ (.Y(_12573_),
    .A(_11134_),
    .B(_11149_));
 sg13g2_a21o_1 _21545_ (.A2(net8711),
    .A1(\soc_I.kianv_I.Instr[25] ),
    .B1(_11122_),
    .X(_12574_));
 sg13g2_nand4_1 _21546_ (.B(_00213_),
    .C(_11210_),
    .A(net9427),
    .Y(_12575_),
    .D(_11236_));
 sg13g2_or4_2 _21547_ (.A(net9431),
    .B(_11098_),
    .C(_12574_),
    .D(_12575_),
    .X(_12576_));
 sg13g2_or2_2 _21548_ (.X(_12577_),
    .B(_12576_),
    .A(_12573_));
 sg13g2_nor2_1 _21549_ (.A(_11164_),
    .B(_12573_),
    .Y(_12578_));
 sg13g2_nand3_1 _21550_ (.B(_11149_),
    .C(_11163_),
    .A(_11134_),
    .Y(_12579_));
 sg13g2_nor3_2 _21551_ (.A(_00213_),
    .B(net8709),
    .C(_11236_),
    .Y(_12580_));
 sg13g2_nand2_1 _21552_ (.Y(_12581_),
    .A(_10898_),
    .B(_12580_));
 sg13g2_nor4_2 _21553_ (.A(\soc_I.kianv_I.Instr[26] ),
    .B(_11088_),
    .C(_12574_),
    .Y(_12582_),
    .D(_12581_));
 sg13g2_and2_1 _21554_ (.A(_12578_),
    .B(_12582_),
    .X(_12583_));
 sg13g2_nor3_1 _21555_ (.A(net9431),
    .B(\soc_I.kianv_I.Instr[26] ),
    .C(\soc_I.kianv_I.Instr[25] ),
    .Y(_12584_));
 sg13g2_nor2_1 _21556_ (.A(net8709),
    .B(_12584_),
    .Y(_12585_));
 sg13g2_nor2_1 _21557_ (.A(_11122_),
    .B(_12585_),
    .Y(_12586_));
 sg13g2_nand2b_2 _21558_ (.Y(_12587_),
    .B(_12586_),
    .A_N(_12575_));
 sg13g2_nor2_2 _21559_ (.A(_12579_),
    .B(_12587_),
    .Y(_12588_));
 sg13g2_nor3_1 _21560_ (.A(net8563),
    .B(_12579_),
    .C(_12587_),
    .Y(_12589_));
 sg13g2_nor2_1 _21561_ (.A(net7934),
    .B(net7928),
    .Y(_12590_));
 sg13g2_nor2b_1 _21562_ (.A(_12581_),
    .B_N(_12586_),
    .Y(_12591_));
 sg13g2_nor3_2 _21563_ (.A(_11163_),
    .B(net8562),
    .C(_12573_),
    .Y(_12592_));
 sg13g2_and2_1 _21564_ (.A(_12591_),
    .B(_12592_),
    .X(_12593_));
 sg13g2_nand3_1 _21565_ (.B(_11150_),
    .C(_11163_),
    .A(_11134_),
    .Y(_12594_));
 sg13g2_or2_1 _21566_ (.X(_12595_),
    .B(_12594_),
    .A(_12587_));
 sg13g2_nand2b_1 _21567_ (.Y(_12596_),
    .B(_12595_),
    .A_N(net7923));
 sg13g2_and2_2 _21568_ (.A(_12578_),
    .B(_12591_),
    .X(_12597_));
 sg13g2_and2_1 _21569_ (.A(_12582_),
    .B(_12592_),
    .X(_12598_));
 sg13g2_nand2_2 _21570_ (.Y(_12599_),
    .A(net8562),
    .B(_12588_));
 sg13g2_and3_1 _21571_ (.X(_12600_),
    .A(net9427),
    .B(_11210_),
    .C(_12584_));
 sg13g2_nand4_1 _21572_ (.B(_12580_),
    .C(_12592_),
    .A(_11122_),
    .Y(_12601_),
    .D(_12600_));
 sg13g2_inv_1 _21573_ (.Y(_12602_),
    .A(_12601_));
 sg13g2_or3_1 _21574_ (.A(net8562),
    .B(_12576_),
    .C(_12594_),
    .X(_12603_));
 sg13g2_nand3_1 _21575_ (.B(_12601_),
    .C(_12603_),
    .A(_12599_),
    .Y(_12604_));
 sg13g2_nor4_1 _21576_ (.A(_12596_),
    .B(net7918),
    .C(net7914),
    .D(_12604_),
    .Y(_12605_));
 sg13g2_nand3_1 _21577_ (.B(_12590_),
    .C(_12605_),
    .A(_12577_),
    .Y(_12606_));
 sg13g2_nor3_2 _21578_ (.A(net9709),
    .B(net9711),
    .C(\soc_I.kianv_I.Instr[9] ),
    .Y(_12607_));
 sg13g2_nor2_1 _21579_ (.A(\soc_I.kianv_I.Instr[8] ),
    .B(\soc_I.kianv_I.Instr[7] ),
    .Y(_12608_));
 sg13g2_nand2_2 _21580_ (.Y(_12609_),
    .A(_12607_),
    .B(_12608_));
 sg13g2_nand2_1 _21581_ (.Y(_12610_),
    .A(_10918_),
    .B(_12609_));
 sg13g2_a21oi_2 _21582_ (.B1(_10970_),
    .Y(_12611_),
    .A2(_12610_),
    .A1(_11002_));
 sg13g2_nand2_2 _21583_ (.Y(_12612_),
    .A(_12606_),
    .B(_12611_));
 sg13g2_nand2_1 _21584_ (.Y(_12613_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[32] ),
    .B(net7913));
 sg13g2_a22oi_1 _21585_ (.Y(_12614_),
    .B1(net7927),
    .B2(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[0] ),
    .A2(net7933),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[32] ));
 sg13g2_nand4_1 _21586_ (.B(_12601_),
    .C(_12613_),
    .A(_12599_),
    .Y(_12615_),
    .D(_12614_));
 sg13g2_nor3_2 _21587_ (.A(_11163_),
    .B(net8563),
    .C(_12577_),
    .Y(_12616_));
 sg13g2_nor3_2 _21588_ (.A(net8563),
    .B(_12576_),
    .C(_12579_),
    .Y(_12617_));
 sg13g2_a221oi_1 _21589_ (.B2(net5577),
    .C1(_12615_),
    .B1(net7904),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[0] ),
    .Y(_12618_),
    .A2(net7807));
 sg13g2_nor3_2 _21590_ (.A(_11164_),
    .B(_11174_),
    .C(_12577_),
    .Y(_12619_));
 sg13g2_nor3_1 _21591_ (.A(_11163_),
    .B(_11174_),
    .C(_12577_),
    .Y(_12620_));
 sg13g2_nor2_1 _21592_ (.A(net8563),
    .B(_12595_),
    .Y(_12621_));
 sg13g2_a22oi_1 _21593_ (.Y(_12622_),
    .B1(net7791),
    .B2(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[0] ),
    .A2(net7923),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[0] ));
 sg13g2_nor2_1 _21594_ (.A(_11174_),
    .B(_12595_),
    .Y(_12623_));
 sg13g2_a22oi_1 _21595_ (.Y(_12624_),
    .B1(net7785),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[0] ),
    .A2(net7918),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[0] ));
 sg13g2_nand2_1 _21596_ (.Y(_12625_),
    .A(_12622_),
    .B(_12624_));
 sg13g2_a221oi_1 _21597_ (.B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[0] ),
    .C1(_12625_),
    .B1(net7796),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[0] ),
    .Y(_12626_),
    .A2(net7802));
 sg13g2_a21oi_2 _21598_ (.B1(net7685),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[0] ),
    .A2(_12626_),
    .A1(_12618_));
 sg13g2_a21oi_1 _21599_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[1] ),
    .A2(net7923),
    .Y(_12627_),
    .B1(_12602_));
 sg13g2_a22oi_1 _21600_ (.Y(_12628_),
    .B1(net7785),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[1] ),
    .A2(net7791),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[1] ));
 sg13g2_a22oi_1 _21601_ (.Y(_12629_),
    .B1(net7904),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[1] ),
    .A2(net7807),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[1] ));
 sg13g2_a22oi_1 _21602_ (.Y(_12630_),
    .B1(net7910),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[33] ),
    .A2(net7934),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[33] ));
 sg13g2_a22oi_1 _21603_ (.Y(_12631_),
    .B1(net7918),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[1] ),
    .A2(net7928),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[1] ));
 sg13g2_nand2_1 _21604_ (.Y(_12632_),
    .A(_12630_),
    .B(_12631_));
 sg13g2_a221oi_1 _21605_ (.B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[1] ),
    .C1(_12632_),
    .B1(net7796),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[1] ),
    .Y(_12633_),
    .A2(net7802));
 sg13g2_nand4_1 _21606_ (.B(_12628_),
    .C(_12629_),
    .A(_12627_),
    .Y(_12634_),
    .D(_12633_));
 sg13g2_nor2b_2 _21607_ (.A(net7685),
    .B_N(_12634_),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[1] ));
 sg13g2_a22oi_1 _21608_ (.Y(_12635_),
    .B1(net7785),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[2] ),
    .A2(net7914),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[34] ));
 sg13g2_a22oi_1 _21609_ (.Y(_12636_),
    .B1(net7923),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[2] ),
    .A2(net7934),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[34] ));
 sg13g2_a22oi_1 _21610_ (.Y(_12637_),
    .B1(net7908),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[2] ),
    .A2(net7811),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[2] ));
 sg13g2_nand2_1 _21611_ (.Y(_12638_),
    .A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[2] ),
    .B(net7791));
 sg13g2_a22oi_1 _21612_ (.Y(_12639_),
    .B1(net7918),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[2] ),
    .A2(net7928),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[2] ));
 sg13g2_nand2_2 _21613_ (.Y(_12640_),
    .A(_12638_),
    .B(_12639_));
 sg13g2_a221oi_1 _21614_ (.B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[2] ),
    .C1(_12640_),
    .B1(net7796),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[2] ),
    .Y(_12641_),
    .A2(net7806));
 sg13g2_nand4_1 _21615_ (.B(_12636_),
    .C(_12637_),
    .A(_12635_),
    .Y(_12642_),
    .D(_12641_));
 sg13g2_nor2b_2 _21616_ (.A(net7689),
    .B_N(_12642_),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[2] ));
 sg13g2_nor4_1 _21617_ (.A(_10645_),
    .B(net8562),
    .C(_12576_),
    .D(_12594_),
    .Y(_12643_));
 sg13g2_a221oi_1 _21618_ (.B2(net4567),
    .C1(_12643_),
    .B1(net7904),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[3] ),
    .Y(_12644_),
    .A2(net7807));
 sg13g2_a22oi_1 _21619_ (.Y(_12645_),
    .B1(net7791),
    .B2(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[3] ),
    .A2(net7934),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[35] ));
 sg13g2_a22oi_1 _21620_ (.Y(_12646_),
    .B1(net7784),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[3] ),
    .A2(net7927),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[3] ));
 sg13g2_a21oi_1 _21621_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[3] ),
    .A2(net7918),
    .Y(_12647_),
    .B1(_12602_));
 sg13g2_a22oi_1 _21622_ (.Y(_12648_),
    .B1(net7913),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[35] ),
    .A2(net7922),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[3] ));
 sg13g2_nand4_1 _21623_ (.B(_12646_),
    .C(_12647_),
    .A(_12645_),
    .Y(_12649_),
    .D(_12648_));
 sg13g2_a221oi_1 _21624_ (.B2(net4660),
    .C1(_12649_),
    .B1(net7796),
    .A1(net4891),
    .Y(_12650_),
    .A2(net7802));
 sg13g2_a21oi_2 _21625_ (.B1(net7685),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[3] ),
    .A2(_12650_),
    .A1(_12644_));
 sg13g2_a22oi_1 _21626_ (.Y(_12651_),
    .B1(net7918),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[4] ),
    .A2(net7928),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[4] ));
 sg13g2_a22oi_1 _21627_ (.Y(_12652_),
    .B1(net7785),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[4] ),
    .A2(net7934),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[36] ));
 sg13g2_a22oi_1 _21628_ (.Y(_12653_),
    .B1(net7908),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[4] ),
    .A2(net7811),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[4] ));
 sg13g2_nand2_1 _21629_ (.Y(_12654_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[4] ),
    .B(net7923));
 sg13g2_a22oi_1 _21630_ (.Y(_12655_),
    .B1(net7791),
    .B2(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[4] ),
    .A2(net7914),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[36] ));
 sg13g2_nand2_1 _21631_ (.Y(_12656_),
    .A(_12654_),
    .B(_12655_));
 sg13g2_a221oi_1 _21632_ (.B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[4] ),
    .C1(_12656_),
    .B1(net7796),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[4] ),
    .Y(_12657_),
    .A2(net7802));
 sg13g2_nand4_1 _21633_ (.B(_12652_),
    .C(_12653_),
    .A(_12651_),
    .Y(_12658_),
    .D(_12657_));
 sg13g2_nor2b_1 _21634_ (.A(net7689),
    .B_N(_12658_),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[4] ));
 sg13g2_a21oi_2 _21635_ (.B1(_12602_),
    .Y(_12659_),
    .A2(net7910),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[37] ));
 sg13g2_a22oi_1 _21636_ (.Y(_12660_),
    .B1(net7791),
    .B2(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[5] ),
    .A2(net7934),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[37] ));
 sg13g2_a22oi_1 _21637_ (.Y(_12661_),
    .B1(net7908),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[5] ),
    .A2(net7811),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[5] ));
 sg13g2_a22oi_1 _21638_ (.Y(_12662_),
    .B1(net7785),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[5] ),
    .A2(net7918),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[5] ));
 sg13g2_a22oi_1 _21639_ (.Y(_12663_),
    .B1(net7923),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[5] ),
    .A2(net7928),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[5] ));
 sg13g2_nand2_1 _21640_ (.Y(_12664_),
    .A(_12662_),
    .B(_12663_));
 sg13g2_a221oi_1 _21641_ (.B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[5] ),
    .C1(_12664_),
    .B1(net7796),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[5] ),
    .Y(_12665_),
    .A2(net7802));
 sg13g2_nand4_1 _21642_ (.B(_12660_),
    .C(_12661_),
    .A(_12659_),
    .Y(_12666_),
    .D(_12665_));
 sg13g2_nor2b_2 _21643_ (.A(net7689),
    .B_N(_12666_),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[5] ));
 sg13g2_a22oi_1 _21644_ (.Y(_12667_),
    .B1(net7785),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[6] ),
    .A2(net7914),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[38] ));
 sg13g2_a22oi_1 _21645_ (.Y(_12668_),
    .B1(net7917),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[6] ),
    .A2(net7934),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[38] ));
 sg13g2_nand2_1 _21646_ (.Y(_12669_),
    .A(_12667_),
    .B(_12668_));
 sg13g2_a221oi_1 _21647_ (.B2(net4554),
    .C1(_12669_),
    .B1(net7908),
    .A1(net2805),
    .Y(_12670_),
    .A2(net7811));
 sg13g2_nand2_1 _21648_ (.Y(_12671_),
    .A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[6] ),
    .B(net7791));
 sg13g2_a22oi_1 _21649_ (.Y(_12672_),
    .B1(net7923),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[6] ),
    .A2(net7928),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[6] ));
 sg13g2_nand2_1 _21650_ (.Y(_12673_),
    .A(_12671_),
    .B(_12672_));
 sg13g2_a221oi_1 _21651_ (.B2(net5124),
    .C1(_12673_),
    .B1(net7796),
    .A1(net4732),
    .Y(_12674_),
    .A2(net7802));
 sg13g2_a21oi_2 _21652_ (.B1(net7689),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[6] ),
    .A2(_12674_),
    .A1(_12670_));
 sg13g2_nor4_1 _21653_ (.A(_10644_),
    .B(net8562),
    .C(_12576_),
    .D(_12594_),
    .Y(_12675_));
 sg13g2_a221oi_1 _21654_ (.B2(net4529),
    .C1(_12675_),
    .B1(net7904),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[7] ),
    .Y(_12676_),
    .A2(net7807));
 sg13g2_nand2_1 _21655_ (.Y(_12677_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[39] ),
    .B(net7910));
 sg13g2_a22oi_1 _21656_ (.Y(_12678_),
    .B1(net7917),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[7] ),
    .A2(net7927),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[7] ));
 sg13g2_a22oi_1 _21657_ (.Y(_12679_),
    .B1(net7784),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[7] ),
    .A2(net7789),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[7] ));
 sg13g2_a22oi_1 _21658_ (.Y(_12680_),
    .B1(net7922),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[7] ),
    .A2(net7933),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[39] ));
 sg13g2_nand4_1 _21659_ (.B(_12678_),
    .C(_12679_),
    .A(_12677_),
    .Y(_12681_),
    .D(_12680_));
 sg13g2_a221oi_1 _21660_ (.B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[7] ),
    .C1(_12681_),
    .B1(net7794),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[7] ),
    .Y(_12682_),
    .A2(net7798));
 sg13g2_a21oi_2 _21661_ (.B1(net7685),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[7] ),
    .A2(_12682_),
    .A1(_12676_));
 sg13g2_nand2_1 _21662_ (.Y(_12683_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[8] ),
    .B(net7917));
 sg13g2_o21ai_1 _21663_ (.B1(_12588_),
    .Y(_12684_),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[8] ),
    .A2(net8562));
 sg13g2_a22oi_1 _21664_ (.Y(_12685_),
    .B1(net7784),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[8] ),
    .A2(net7933),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[40] ));
 sg13g2_nand3_1 _21665_ (.B(_12684_),
    .C(_12685_),
    .A(_12683_),
    .Y(_12686_));
 sg13g2_a221oi_1 _21666_ (.B2(net4464),
    .C1(_12686_),
    .B1(net7907),
    .A1(net2802),
    .Y(_12687_),
    .A2(net7810));
 sg13g2_nand2_1 _21667_ (.Y(_12688_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[8] ),
    .B(net7922));
 sg13g2_a22oi_1 _21668_ (.Y(_12689_),
    .B1(net7789),
    .B2(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[8] ),
    .A2(net7910),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[40] ));
 sg13g2_nand2_1 _21669_ (.Y(_12690_),
    .A(_12688_),
    .B(_12689_));
 sg13g2_a221oi_1 _21670_ (.B2(net4396),
    .C1(_12690_),
    .B1(net7794),
    .A1(net4670),
    .Y(_12691_),
    .A2(net7798));
 sg13g2_a21oi_2 _21671_ (.B1(net7685),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[8] ),
    .A2(_12691_),
    .A1(_12687_));
 sg13g2_a22oi_1 _21672_ (.Y(_12692_),
    .B1(net7784),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[9] ),
    .A2(net7922),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[9] ));
 sg13g2_a22oi_1 _21673_ (.Y(_12693_),
    .B1(net7910),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[41] ),
    .A2(net7917),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[9] ));
 sg13g2_a22oi_1 _21674_ (.Y(_12694_),
    .B1(net7904),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[9] ),
    .A2(net7807),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[9] ));
 sg13g2_nand2_1 _21675_ (.Y(_12695_),
    .A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[9] ),
    .B(net7789));
 sg13g2_a22oi_1 _21676_ (.Y(_12696_),
    .B1(net7927),
    .B2(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[9] ),
    .A2(net7933),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[41] ));
 sg13g2_nand2_1 _21677_ (.Y(_12697_),
    .A(_12695_),
    .B(_12696_));
 sg13g2_a221oi_1 _21678_ (.B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[9] ),
    .C1(_12697_),
    .B1(net7794),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[9] ),
    .Y(_12698_),
    .A2(net7798));
 sg13g2_nand4_1 _21679_ (.B(_12693_),
    .C(_12694_),
    .A(_12692_),
    .Y(_12699_),
    .D(_12698_));
 sg13g2_nor2b_2 _21680_ (.A(net7685),
    .B_N(_12699_),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[9] ));
 sg13g2_a22oi_1 _21681_ (.Y(_12700_),
    .B1(net7784),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[10] ),
    .A2(net7922),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[10] ));
 sg13g2_a22oi_1 _21682_ (.Y(_12701_),
    .B1(net7789),
    .B2(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[10] ),
    .A2(net7933),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[42] ));
 sg13g2_a22oi_1 _21683_ (.Y(_12702_),
    .B1(net7904),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[10] ),
    .A2(net7807),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[10] ));
 sg13g2_nand2_1 _21684_ (.Y(_12703_),
    .A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[10] ),
    .B(net7927));
 sg13g2_a22oi_1 _21685_ (.Y(_12704_),
    .B1(net7910),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[42] ),
    .A2(net7917),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[10] ));
 sg13g2_nand2_1 _21686_ (.Y(_12705_),
    .A(_12703_),
    .B(_12704_));
 sg13g2_a221oi_1 _21687_ (.B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[10] ),
    .C1(_12705_),
    .B1(net7794),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[10] ),
    .Y(_12706_),
    .A2(net7798));
 sg13g2_nand4_1 _21688_ (.B(_12701_),
    .C(_12702_),
    .A(_12700_),
    .Y(_12707_),
    .D(_12706_));
 sg13g2_nor2b_2 _21689_ (.A(net7687),
    .B_N(_12707_),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[10] ));
 sg13g2_a22oi_1 _21690_ (.Y(_12708_),
    .B1(net7789),
    .B2(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[11] ),
    .A2(net7927),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[11] ));
 sg13g2_a22oi_1 _21691_ (.Y(_12709_),
    .B1(net7784),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[11] ),
    .A2(net7910),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[43] ));
 sg13g2_nand2_1 _21692_ (.Y(_12710_),
    .A(_12708_),
    .B(_12709_));
 sg13g2_a221oi_1 _21693_ (.B2(net4539),
    .C1(_12710_),
    .B1(net7904),
    .A1(net2656),
    .Y(_12711_),
    .A2(net7807));
 sg13g2_nand2_1 _21694_ (.Y(_12712_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[43] ),
    .B(net7933));
 sg13g2_a22oi_1 _21695_ (.Y(_12713_),
    .B1(net7917),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[11] ),
    .A2(net7922),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[11] ));
 sg13g2_nand2_1 _21696_ (.Y(_12714_),
    .A(_12712_),
    .B(_12713_));
 sg13g2_a221oi_1 _21697_ (.B2(net4757),
    .C1(_12714_),
    .B1(net7794),
    .A1(net4598),
    .Y(_12715_),
    .A2(net7798));
 sg13g2_a21oi_2 _21698_ (.B1(net7685),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[11] ),
    .A2(_12715_),
    .A1(_12711_));
 sg13g2_nand2_1 _21699_ (.Y(_12716_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[12] ),
    .B(net7917));
 sg13g2_o21ai_1 _21700_ (.B1(_12588_),
    .Y(_12717_),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[12] ),
    .A2(net8562));
 sg13g2_a22oi_1 _21701_ (.Y(_12718_),
    .B1(net7910),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[44] ),
    .A2(net7920),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[12] ));
 sg13g2_nand3_1 _21702_ (.B(_12717_),
    .C(_12718_),
    .A(_12716_),
    .Y(_12719_));
 sg13g2_a221oi_1 _21703_ (.B2(net4665),
    .C1(_12719_),
    .B1(net7904),
    .A1(net2696),
    .Y(_12720_),
    .A2(net7807));
 sg13g2_nand2_1 _21704_ (.Y(_12721_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[12] ),
    .B(net7784));
 sg13g2_a22oi_1 _21705_ (.Y(_12722_),
    .B1(net7789),
    .B2(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[12] ),
    .A2(net7933),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[44] ));
 sg13g2_nand2_1 _21706_ (.Y(_12723_),
    .A(_12721_),
    .B(_12722_));
 sg13g2_a221oi_1 _21707_ (.B2(net4744),
    .C1(_12723_),
    .B1(net7794),
    .A1(net4295),
    .Y(_12724_),
    .A2(net7801));
 sg13g2_a21oi_2 _21708_ (.B1(net7685),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[12] ),
    .A2(_12724_),
    .A1(_12720_));
 sg13g2_a22oi_1 _21709_ (.Y(_12725_),
    .B1(net7782),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[13] ),
    .A2(net7931),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[45] ));
 sg13g2_a22oi_1 _21710_ (.Y(_12726_),
    .B1(net7788),
    .B2(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[13] ),
    .A2(net7920),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[13] ));
 sg13g2_a22oi_1 _21711_ (.Y(_12727_),
    .B1(net7905),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[13] ),
    .A2(net7808),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[13] ));
 sg13g2_nand2_1 _21712_ (.Y(_12728_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[45] ),
    .B(net7911));
 sg13g2_a22oi_1 _21713_ (.Y(_12729_),
    .B1(net7915),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[13] ),
    .A2(net7925),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[13] ));
 sg13g2_nand2_1 _21714_ (.Y(_12730_),
    .A(_12728_),
    .B(_12729_));
 sg13g2_a221oi_1 _21715_ (.B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[13] ),
    .C1(_12730_),
    .B1(net7793),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[13] ),
    .Y(_12731_),
    .A2(net7799));
 sg13g2_nand4_1 _21716_ (.B(_12726_),
    .C(_12727_),
    .A(_12725_),
    .Y(_12732_),
    .D(_12731_));
 sg13g2_nor2b_1 _21717_ (.A(net7686),
    .B_N(_12732_),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[13] ));
 sg13g2_a22oi_1 _21718_ (.Y(_12733_),
    .B1(net7788),
    .B2(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[14] ),
    .A2(net7931),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[46] ));
 sg13g2_a22oi_1 _21719_ (.Y(_12734_),
    .B1(net7782),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[14] ),
    .A2(net7911),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[46] ));
 sg13g2_a22oi_1 _21720_ (.Y(_12735_),
    .B1(net7905),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[14] ),
    .A2(net7808),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[14] ));
 sg13g2_nand2_1 _21721_ (.Y(_12736_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[14] ),
    .B(net7915));
 sg13g2_a22oi_1 _21722_ (.Y(_12737_),
    .B1(net7920),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[14] ),
    .A2(net7925),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[14] ));
 sg13g2_nand2_1 _21723_ (.Y(_12738_),
    .A(_12736_),
    .B(_12737_));
 sg13g2_a221oi_1 _21724_ (.B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[14] ),
    .C1(_12738_),
    .B1(net7793),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[14] ),
    .Y(_12739_),
    .A2(net7799));
 sg13g2_nand4_1 _21725_ (.B(_12734_),
    .C(_12735_),
    .A(_12733_),
    .Y(_12740_),
    .D(_12739_));
 sg13g2_nor2b_1 _21726_ (.A(net7687),
    .B_N(_12740_),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[14] ));
 sg13g2_a22oi_1 _21727_ (.Y(_12741_),
    .B1(net7788),
    .B2(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[15] ),
    .A2(net7911),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[47] ));
 sg13g2_a22oi_1 _21728_ (.Y(_12742_),
    .B1(net7782),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[15] ),
    .A2(net7925),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[15] ));
 sg13g2_nand2_1 _21729_ (.Y(_12743_),
    .A(_12741_),
    .B(_12742_));
 sg13g2_a221oi_1 _21730_ (.B2(net4453),
    .C1(_12743_),
    .B1(net7905),
    .A1(net2803),
    .Y(_12744_),
    .A2(net7808));
 sg13g2_nand2_1 _21731_ (.Y(_12745_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[47] ),
    .B(net7931));
 sg13g2_a22oi_1 _21732_ (.Y(_12746_),
    .B1(net7915),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[15] ),
    .A2(net7920),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[15] ));
 sg13g2_nand2_2 _21733_ (.Y(_12747_),
    .A(_12745_),
    .B(_12746_));
 sg13g2_a221oi_1 _21734_ (.B2(net4349),
    .C1(_12747_),
    .B1(net7793),
    .A1(net4910),
    .Y(_12748_),
    .A2(net7799));
 sg13g2_a21oi_2 _21735_ (.B1(net7686),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[15] ),
    .A2(_12748_),
    .A1(_12744_));
 sg13g2_a22oi_1 _21736_ (.Y(_12749_),
    .B1(net7920),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[16] ),
    .A2(net7925),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[16] ));
 sg13g2_a22oi_1 _21737_ (.Y(_12750_),
    .B1(net7782),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[16] ),
    .A2(net7788),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[16] ));
 sg13g2_a22oi_1 _21738_ (.Y(_12751_),
    .B1(net7905),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[16] ),
    .A2(net7808),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[16] ));
 sg13g2_nand2_1 _21739_ (.Y(_12752_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[48] ),
    .B(net7931));
 sg13g2_a22oi_1 _21740_ (.Y(_12753_),
    .B1(net7911),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[48] ),
    .A2(net7915),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[16] ));
 sg13g2_nand2_1 _21741_ (.Y(_12754_),
    .A(_12752_),
    .B(_12753_));
 sg13g2_a221oi_1 _21742_ (.B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[16] ),
    .C1(_12754_),
    .B1(net7793),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[16] ),
    .Y(_12755_),
    .A2(net7799));
 sg13g2_nand4_1 _21743_ (.B(_12750_),
    .C(_12751_),
    .A(_12749_),
    .Y(_12756_),
    .D(_12755_));
 sg13g2_nor2b_1 _21744_ (.A(net7686),
    .B_N(_12756_),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[16] ));
 sg13g2_a22oi_1 _21745_ (.Y(_12757_),
    .B1(net7915),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[17] ),
    .A2(net7932),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[49] ));
 sg13g2_a22oi_1 _21746_ (.Y(_12758_),
    .B1(net7788),
    .B2(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[17] ),
    .A2(net7920),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[17] ));
 sg13g2_nand2_1 _21747_ (.Y(_12759_),
    .A(_12757_),
    .B(_12758_));
 sg13g2_a221oi_1 _21748_ (.B2(net4445),
    .C1(_12759_),
    .B1(net7905),
    .A1(net2777),
    .Y(_12760_),
    .A2(net7808));
 sg13g2_nand2_1 _21749_ (.Y(_12761_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[17] ),
    .B(net7782));
 sg13g2_a22oi_1 _21750_ (.Y(_12762_),
    .B1(net7912),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[49] ),
    .A2(net7925),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[17] ));
 sg13g2_nand2_1 _21751_ (.Y(_12763_),
    .A(_12761_),
    .B(_12762_));
 sg13g2_a221oi_1 _21752_ (.B2(net4357),
    .C1(_12763_),
    .B1(net7793),
    .A1(net4883),
    .Y(_12764_),
    .A2(net7799));
 sg13g2_a21oi_2 _21753_ (.B1(net7686),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[17] ),
    .A2(_12764_),
    .A1(_12760_));
 sg13g2_a22oi_1 _21754_ (.Y(_12765_),
    .B1(net7916),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[18] ),
    .A2(net7925),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[18] ));
 sg13g2_a22oi_1 _21755_ (.Y(_12766_),
    .B1(net7782),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[18] ),
    .A2(net7921),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[18] ));
 sg13g2_a22oi_1 _21756_ (.Y(_12767_),
    .B1(net7905),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[18] ),
    .A2(net7808),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[18] ));
 sg13g2_nand2_1 _21757_ (.Y(_12768_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[50] ),
    .B(net7931));
 sg13g2_a22oi_1 _21758_ (.Y(_12769_),
    .B1(net7788),
    .B2(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[18] ),
    .A2(net7911),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[50] ));
 sg13g2_nand2_1 _21759_ (.Y(_12770_),
    .A(_12768_),
    .B(_12769_));
 sg13g2_a221oi_1 _21760_ (.B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[18] ),
    .C1(_12770_),
    .B1(net7793),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[18] ),
    .Y(_12771_),
    .A2(net7799));
 sg13g2_nand4_1 _21761_ (.B(_12766_),
    .C(_12767_),
    .A(_12765_),
    .Y(_12772_),
    .D(_12771_));
 sg13g2_nor2b_2 _21762_ (.A(net7686),
    .B_N(_12772_),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[18] ));
 sg13g2_a22oi_1 _21763_ (.Y(_12773_),
    .B1(net7911),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[51] ),
    .A2(net7931),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[51] ));
 sg13g2_a22oi_1 _21764_ (.Y(_12774_),
    .B1(net7782),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[19] ),
    .A2(net7925),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[19] ));
 sg13g2_a22oi_1 _21765_ (.Y(_12775_),
    .B1(net7905),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[19] ),
    .A2(net7808),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[19] ));
 sg13g2_nand2_1 _21766_ (.Y(_12776_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[19] ),
    .B(net7921));
 sg13g2_a22oi_1 _21767_ (.Y(_12777_),
    .B1(net7788),
    .B2(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[19] ),
    .A2(net7915),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[19] ));
 sg13g2_nand2_1 _21768_ (.Y(_12778_),
    .A(_12776_),
    .B(_12777_));
 sg13g2_a221oi_1 _21769_ (.B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[19] ),
    .C1(_12778_),
    .B1(net7793),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[19] ),
    .Y(_12779_),
    .A2(net7799));
 sg13g2_nand4_1 _21770_ (.B(_12774_),
    .C(_12775_),
    .A(_12773_),
    .Y(_12780_),
    .D(_12779_));
 sg13g2_nor2b_2 _21771_ (.A(net7686),
    .B_N(_12780_),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[19] ));
 sg13g2_nand2_1 _21772_ (.Y(_12781_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[20] ),
    .B(net7785));
 sg13g2_a22oi_1 _21773_ (.Y(_12782_),
    .B1(net7916),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[20] ),
    .A2(net7926),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[20] ));
 sg13g2_nand3_1 _21774_ (.B(_12781_),
    .C(_12782_),
    .A(_12599_),
    .Y(_12783_));
 sg13g2_a221oi_1 _21775_ (.B2(net4538),
    .C1(_12783_),
    .B1(net7908),
    .A1(net2638),
    .Y(_12784_),
    .A2(net7811));
 sg13g2_a22oi_1 _21776_ (.Y(_12785_),
    .B1(net7788),
    .B2(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[20] ),
    .A2(net7911),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[52] ));
 sg13g2_a22oi_1 _21777_ (.Y(_12786_),
    .B1(net7921),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[20] ),
    .A2(net7931),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[52] ));
 sg13g2_nand2_2 _21778_ (.Y(_12787_),
    .A(_12785_),
    .B(_12786_));
 sg13g2_a221oi_1 _21779_ (.B2(net4678),
    .C1(_12787_),
    .B1(net7795),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[20] ),
    .Y(_12788_),
    .A2(net7805));
 sg13g2_a21oi_2 _21780_ (.B1(net7688),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[20] ),
    .A2(_12788_),
    .A1(_12784_));
 sg13g2_a22oi_1 _21781_ (.Y(_12789_),
    .B1(net7790),
    .B2(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[21] ),
    .A2(net7914),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[53] ));
 sg13g2_a22oi_1 _21782_ (.Y(_12790_),
    .B1(net7786),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[21] ),
    .A2(net7929),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[21] ));
 sg13g2_nand2_1 _21783_ (.Y(_12791_),
    .A(_12789_),
    .B(_12790_));
 sg13g2_a221oi_1 _21784_ (.B2(net4373),
    .C1(_12791_),
    .B1(net7909),
    .A1(net2667),
    .Y(_12792_),
    .A2(net7812));
 sg13g2_nand2_1 _21785_ (.Y(_12793_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[21] ),
    .B(net7915));
 sg13g2_a22oi_1 _21786_ (.Y(_12794_),
    .B1(net7920),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[21] ),
    .A2(net7931),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[53] ));
 sg13g2_nand2_2 _21787_ (.Y(_12795_),
    .A(_12793_),
    .B(_12794_));
 sg13g2_a221oi_1 _21788_ (.B2(net4727),
    .C1(_12795_),
    .B1(net7797),
    .A1(net5522),
    .Y(_12796_),
    .A2(net7803));
 sg13g2_a21oi_2 _21789_ (.B1(net7688),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[21] ),
    .A2(_12796_),
    .A1(_12792_));
 sg13g2_a22oi_1 _21790_ (.Y(_12797_),
    .B1(net7929),
    .B2(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[22] ),
    .A2(net7935),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[54] ));
 sg13g2_a22oi_1 _21791_ (.Y(_12798_),
    .B1(net7786),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[22] ),
    .A2(net7792),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[22] ));
 sg13g2_nand2_1 _21792_ (.Y(_12799_),
    .A(_12797_),
    .B(_12798_));
 sg13g2_a221oi_1 _21793_ (.B2(net4385),
    .C1(_12799_),
    .B1(net7909),
    .A1(net2668),
    .Y(_12800_),
    .A2(net7812));
 sg13g2_nand2_1 _21794_ (.Y(_12801_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[54] ),
    .B(net7911));
 sg13g2_a22oi_1 _21795_ (.Y(_12802_),
    .B1(net7915),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[22] ),
    .A2(net7920),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[22] ));
 sg13g2_nand2_2 _21796_ (.Y(_12803_),
    .A(_12801_),
    .B(_12802_));
 sg13g2_a221oi_1 _21797_ (.B2(net4741),
    .C1(_12803_),
    .B1(net7795),
    .A1(net4840),
    .Y(_12804_),
    .A2(net7804));
 sg13g2_a21oi_2 _21798_ (.B1(net7689),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[22] ),
    .A2(_12804_),
    .A1(_12800_));
 sg13g2_a22oi_1 _21799_ (.Y(_12805_),
    .B1(net7790),
    .B2(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[23] ),
    .A2(net7924),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[23] ));
 sg13g2_a22oi_1 _21800_ (.Y(_12806_),
    .B1(net7913),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[55] ),
    .A2(net7935),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[55] ));
 sg13g2_a22oi_1 _21801_ (.Y(_12807_),
    .B1(net7909),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[23] ),
    .A2(net7812),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[23] ));
 sg13g2_nand2_1 _21802_ (.Y(_12808_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[23] ),
    .B(net7786));
 sg13g2_a22oi_1 _21803_ (.Y(_12809_),
    .B1(net7919),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[23] ),
    .A2(net7929),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[23] ));
 sg13g2_nand2_1 _21804_ (.Y(_12810_),
    .A(_12808_),
    .B(_12809_));
 sg13g2_a221oi_1 _21805_ (.B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[23] ),
    .C1(_12810_),
    .B1(net7795),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[23] ),
    .Y(_12811_),
    .A2(net7805));
 sg13g2_nand4_1 _21806_ (.B(_12806_),
    .C(_12807_),
    .A(_12805_),
    .Y(_12812_),
    .D(_12811_));
 sg13g2_nor2b_2 _21807_ (.A(net7688),
    .B_N(_12812_),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[23] ));
 sg13g2_a22oi_1 _21808_ (.Y(_12813_),
    .B1(net7790),
    .B2(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[24] ),
    .A2(net7924),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[24] ));
 sg13g2_a22oi_1 _21809_ (.Y(_12814_),
    .B1(net7919),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[24] ),
    .A2(net7928),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[24] ));
 sg13g2_nand2_1 _21810_ (.Y(_12815_),
    .A(_12813_),
    .B(_12814_));
 sg13g2_a221oi_1 _21811_ (.B2(net4471),
    .C1(_12815_),
    .B1(net7908),
    .A1(net2772),
    .Y(_12816_),
    .A2(net7811));
 sg13g2_nand2_1 _21812_ (.Y(_12817_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[56] ),
    .B(net7932));
 sg13g2_a22oi_1 _21813_ (.Y(_12818_),
    .B1(net7782),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[24] ),
    .A2(net7912),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[56] ));
 sg13g2_nand2_2 _21814_ (.Y(_12819_),
    .A(_12817_),
    .B(_12818_));
 sg13g2_a221oi_1 _21815_ (.B2(net4577),
    .C1(_12819_),
    .B1(net7795),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[24] ),
    .Y(_12820_),
    .A2(net7803));
 sg13g2_a21oi_2 _21816_ (.B1(net7688),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[24] ),
    .A2(_12820_),
    .A1(_12816_));
 sg13g2_a22oi_1 _21817_ (.Y(_12821_),
    .B1(net7914),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[57] ),
    .A2(net7919),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[25] ));
 sg13g2_a22oi_1 _21818_ (.Y(_12822_),
    .B1(net7786),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[25] ),
    .A2(net7792),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[25] ));
 sg13g2_a22oi_1 _21819_ (.Y(_12823_),
    .B1(net7908),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[25] ),
    .A2(net7811),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[25] ));
 sg13g2_nand2_1 _21820_ (.Y(_12824_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[25] ),
    .B(net7922));
 sg13g2_a22oi_1 _21821_ (.Y(_12825_),
    .B1(net7925),
    .B2(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[25] ),
    .A2(net7935),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[57] ));
 sg13g2_nand2_2 _21822_ (.Y(_12826_),
    .A(_12824_),
    .B(_12825_));
 sg13g2_a221oi_1 _21823_ (.B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[25] ),
    .C1(_12826_),
    .B1(net7795),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[25] ),
    .Y(_12827_),
    .A2(net7803));
 sg13g2_nand4_1 _21824_ (.B(_12822_),
    .C(_12823_),
    .A(_12821_),
    .Y(_12828_),
    .D(_12827_));
 sg13g2_nor2b_2 _21825_ (.A(net7688),
    .B_N(_12828_),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[25] ));
 sg13g2_a22oi_1 _21826_ (.Y(_12829_),
    .B1(net7924),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[26] ),
    .A2(net7928),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[26] ));
 sg13g2_a22oi_1 _21827_ (.Y(_12830_),
    .B1(net7786),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[26] ),
    .A2(net7790),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[26] ));
 sg13g2_a22oi_1 _21828_ (.Y(_12831_),
    .B1(net7908),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[26] ),
    .A2(net7811),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[26] ));
 sg13g2_nand2_1 _21829_ (.Y(_12832_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[26] ),
    .B(net7918));
 sg13g2_a22oi_1 _21830_ (.Y(_12833_),
    .B1(net7912),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[58] ),
    .A2(net7932),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[58] ));
 sg13g2_nand2_2 _21831_ (.Y(_12834_),
    .A(_12832_),
    .B(_12833_));
 sg13g2_a221oi_1 _21832_ (.B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[26] ),
    .C1(_12834_),
    .B1(net7795),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[26] ),
    .Y(_12835_),
    .A2(net7803));
 sg13g2_nand4_1 _21833_ (.B(_12830_),
    .C(_12831_),
    .A(_12829_),
    .Y(_12836_),
    .D(_12835_));
 sg13g2_nor2b_2 _21834_ (.A(net7688),
    .B_N(_12836_),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[26] ));
 sg13g2_a22oi_1 _21835_ (.Y(_12837_),
    .B1(net7785),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[27] ),
    .A2(net7914),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[59] ));
 sg13g2_a22oi_1 _21836_ (.Y(_12838_),
    .B1(net7790),
    .B2(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[27] ),
    .A2(net7934),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[59] ));
 sg13g2_a22oi_1 _21837_ (.Y(_12839_),
    .B1(net7909),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[27] ),
    .A2(net7812),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[27] ));
 sg13g2_nand2_1 _21838_ (.Y(_12840_),
    .A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[27] ),
    .B(net7929));
 sg13g2_a22oi_1 _21839_ (.Y(_12841_),
    .B1(net7919),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[27] ),
    .A2(net7923),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[27] ));
 sg13g2_nand2_1 _21840_ (.Y(_12842_),
    .A(_12840_),
    .B(_12841_));
 sg13g2_a221oi_1 _21841_ (.B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[27] ),
    .C1(_12842_),
    .B1(net7795),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[27] ),
    .Y(_12843_),
    .A2(net7805));
 sg13g2_nand4_1 _21842_ (.B(_12838_),
    .C(_12839_),
    .A(_12837_),
    .Y(_12844_),
    .D(_12843_));
 sg13g2_nor2b_1 _21843_ (.A(net7688),
    .B_N(_12844_),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[27] ));
 sg13g2_a22oi_1 _21844_ (.Y(_12845_),
    .B1(net7790),
    .B2(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[28] ),
    .A2(net7919),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[28] ));
 sg13g2_a22oi_1 _21845_ (.Y(_12846_),
    .B1(net7912),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[60] ),
    .A2(net7926),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[28] ));
 sg13g2_a22oi_1 _21846_ (.Y(_12847_),
    .B1(net7906),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[28] ),
    .A2(net7809),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[28] ));
 sg13g2_nand2_1 _21847_ (.Y(_12848_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[28] ),
    .B(net7783));
 sg13g2_a22oi_1 _21848_ (.Y(_12849_),
    .B1(net7921),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[28] ),
    .A2(net7932),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[60] ));
 sg13g2_nand2_1 _21849_ (.Y(_12850_),
    .A(_12848_),
    .B(_12849_));
 sg13g2_a221oi_1 _21850_ (.B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[28] ),
    .C1(_12850_),
    .B1(net7794),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[28] ),
    .Y(_12851_),
    .A2(net7800));
 sg13g2_nand4_1 _21851_ (.B(_12846_),
    .C(_12847_),
    .A(_12845_),
    .Y(_12852_),
    .D(_12851_));
 sg13g2_nor2b_2 _21852_ (.A(net7688),
    .B_N(_12852_),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[28] ));
 sg13g2_a22oi_1 _21853_ (.Y(_12853_),
    .B1(net7921),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[29] ),
    .A2(net7932),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[61] ));
 sg13g2_a22oi_1 _21854_ (.Y(_12854_),
    .B1(net7783),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[29] ),
    .A2(net7912),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[61] ));
 sg13g2_a22oi_1 _21855_ (.Y(_12855_),
    .B1(net7905),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[29] ),
    .A2(net7808),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[29] ));
 sg13g2_nand2_1 _21856_ (.Y(_12856_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[29] ),
    .B(net7919));
 sg13g2_a22oi_1 _21857_ (.Y(_12857_),
    .B1(net7790),
    .B2(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[29] ),
    .A2(net7929),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[29] ));
 sg13g2_nand2_1 _21858_ (.Y(_12858_),
    .A(_12856_),
    .B(_12857_));
 sg13g2_a221oi_1 _21859_ (.B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[29] ),
    .C1(_12858_),
    .B1(net7795),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[29] ),
    .Y(_12859_),
    .A2(net7805));
 sg13g2_nand4_1 _21860_ (.B(_12854_),
    .C(_12855_),
    .A(_12853_),
    .Y(_12860_),
    .D(_12859_));
 sg13g2_nor2b_2 _21861_ (.A(net7686),
    .B_N(_12860_),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[29] ));
 sg13g2_nand2_1 _21862_ (.Y(_12861_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[30] ),
    .B(net7783));
 sg13g2_a22oi_1 _21863_ (.Y(_12862_),
    .B1(net7926),
    .B2(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[30] ),
    .A2(net7932),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[62] ));
 sg13g2_nand3_1 _21864_ (.B(_12861_),
    .C(_12862_),
    .A(_12599_),
    .Y(_12863_));
 sg13g2_a221oi_1 _21865_ (.B2(net4579),
    .C1(_12863_),
    .B1(net7906),
    .A1(net2739),
    .Y(_12864_),
    .A2(net7809));
 sg13g2_a22oi_1 _21866_ (.Y(_12865_),
    .B1(net7916),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[30] ),
    .A2(net7921),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[30] ));
 sg13g2_a22oi_1 _21867_ (.Y(_12866_),
    .B1(net7792),
    .B2(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[30] ),
    .A2(net7912),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[62] ));
 sg13g2_nand2_1 _21868_ (.Y(_12867_),
    .A(_12865_),
    .B(_12866_));
 sg13g2_a221oi_1 _21869_ (.B2(net4505),
    .C1(_12867_),
    .B1(net7797),
    .A1(net4711),
    .Y(_12868_),
    .A2(net7800));
 sg13g2_a21oi_2 _21870_ (.B1(net7687),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[30] ),
    .A2(_12868_),
    .A1(_12864_));
 sg13g2_a22oi_1 _21871_ (.Y(_12869_),
    .B1(net7912),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[63] ),
    .A2(net7926),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[31] ));
 sg13g2_a22oi_1 _21872_ (.Y(_12870_),
    .B1(net7789),
    .B2(net4481),
    .A2(net7916),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[31] ));
 sg13g2_a22oi_1 _21873_ (.Y(_12871_),
    .B1(net7906),
    .B2(net5562),
    .A2(net7809),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[31] ));
 sg13g2_nand2_1 _21874_ (.Y(_12872_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[31] ),
    .B(net7783));
 sg13g2_a22oi_1 _21875_ (.Y(_12873_),
    .B1(net7921),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[31] ),
    .A2(net7932),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[63] ));
 sg13g2_nand2_1 _21876_ (.Y(_12874_),
    .A(_12872_),
    .B(_12873_));
 sg13g2_a221oi_1 _21877_ (.B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[31] ),
    .C1(_12874_),
    .B1(net7793),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[31] ),
    .Y(_12875_),
    .A2(net7800));
 sg13g2_nand4_1 _21878_ (.B(_12870_),
    .C(_12871_),
    .A(_12869_),
    .Y(_12876_),
    .D(_12875_));
 sg13g2_nor2b_1 _21879_ (.A(net7686),
    .B_N(_12876_),
    .Y(\soc_I.kianv_I.datapath_unit_I.CSRData[31] ));
 sg13g2_nor2_1 _21880_ (.A(net9244),
    .B(net9292),
    .Y(_12877_));
 sg13g2_nand2_2 _21881_ (.Y(_12878_),
    .A(net9000),
    .B(_10604_));
 sg13g2_nor2_2 _21882_ (.A(\soc_I.spi0_I.ready_xfer ),
    .B(\soc_I.spi0_I.ready_ctrl ),
    .Y(_12879_));
 sg13g2_or2_1 _21883_ (.X(_12880_),
    .B(\soc_I.spi0_I.ready_ctrl ),
    .A(\soc_I.spi0_I.ready_xfer ));
 sg13g2_nor4_1 _21884_ (.A(\soc_I.gpio0_I.ready ),
    .B(net9250),
    .C(_12878_),
    .D(net8960),
    .Y(_12881_));
 sg13g2_and3_1 _21885_ (.X(_12882_),
    .A(_00250_),
    .B(_12877_),
    .C(_12881_));
 sg13g2_nor3_2 _21886_ (.A(_11757_),
    .B(_11758_),
    .C(\soc_I.clint_I.addr[1] ),
    .Y(_12883_));
 sg13g2_nand2_1 _21887_ (.Y(_12884_),
    .A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[2] ),
    .B(net8839));
 sg13g2_a21oi_1 _21888_ (.A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[2] ),
    .A2(net8704),
    .Y(_12885_),
    .B1(net8699));
 sg13g2_o21ai_1 _21889_ (.B1(net8663),
    .Y(_12886_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[2] ),
    .A2(net8693));
 sg13g2_a21oi_1 _21890_ (.A1(_12884_),
    .A2(_12885_),
    .Y(_12887_),
    .B1(_12886_));
 sg13g2_nor2_1 _21891_ (.A(net8707),
    .B(_12887_),
    .Y(_12888_));
 sg13g2_o21ai_1 _21892_ (.B1(_12888_),
    .Y(_12889_),
    .A1(net8662),
    .A2(_11936_));
 sg13g2_a21oi_1 _21893_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[2] ),
    .A2(net8734),
    .Y(_12890_),
    .B1(net8631));
 sg13g2_nor2_2 _21894_ (.A(net8502),
    .B(_12890_),
    .Y(_12891_));
 sg13g2_a22oi_1 _21895_ (.Y(_12892_),
    .B1(_12889_),
    .B2(_12891_),
    .A2(net8377),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[2] ));
 sg13g2_nor2_2 _21896_ (.A(\soc_I.PC[2] ),
    .B(net8576),
    .Y(_12893_));
 sg13g2_a21oi_1 _21897_ (.A1(net8572),
    .A2(net7618),
    .Y(_12894_),
    .B1(_12893_));
 sg13g2_a21o_2 _21898_ (.A2(net7618),
    .A1(net8572),
    .B1(_12893_),
    .X(_12895_));
 sg13g2_nor2_1 _21899_ (.A(\soc_I.PC[3] ),
    .B(net8575),
    .Y(_12896_));
 sg13g2_nand2_1 _21900_ (.Y(_12897_),
    .A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[3] ),
    .B(net8841));
 sg13g2_a21oi_1 _21901_ (.A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[3] ),
    .A2(net8703),
    .Y(_12898_),
    .B1(net8698));
 sg13g2_o21ai_1 _21902_ (.B1(net8657),
    .Y(_12899_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[3] ),
    .A2(net8691));
 sg13g2_a21oi_1 _21903_ (.A1(_12897_),
    .A2(_12898_),
    .Y(_12900_),
    .B1(_12899_));
 sg13g2_nor2_1 _21904_ (.A(net8706),
    .B(_12900_),
    .Y(_12901_));
 sg13g2_o21ai_1 _21905_ (.B1(_12901_),
    .Y(_12902_),
    .A1(net8657),
    .A2(_12376_));
 sg13g2_a21oi_1 _21906_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[3] ),
    .A2(net8733),
    .Y(_12903_),
    .B1(net8630));
 sg13g2_nor2_1 _21907_ (.A(net8501),
    .B(_12903_),
    .Y(_12904_));
 sg13g2_a22oi_1 _21908_ (.Y(_12905_),
    .B1(_12902_),
    .B2(_12904_),
    .A2(net8376),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[3] ));
 sg13g2_a21oi_2 _21909_ (.B1(_12896_),
    .Y(_12906_),
    .A2(_12905_),
    .A1(net8575));
 sg13g2_or2_1 _21910_ (.X(_12907_),
    .B(_12906_),
    .A(net7493));
 sg13g2_inv_1 _21911_ (.Y(_12908_),
    .A(_12907_));
 sg13g2_nor2_1 _21912_ (.A(\soc_I.PC[7] ),
    .B(net8573),
    .Y(_12909_));
 sg13g2_nand2_1 _21913_ (.Y(_12910_),
    .A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[7] ),
    .B(net8838));
 sg13g2_a21oi_2 _21914_ (.B1(net8698),
    .Y(_12911_),
    .A2(net8703),
    .A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[7] ));
 sg13g2_o21ai_1 _21915_ (.B1(net8658),
    .Y(_12912_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[7] ),
    .A2(net8695));
 sg13g2_a21oi_1 _21916_ (.A1(_12910_),
    .A2(_12911_),
    .Y(_12913_),
    .B1(_12912_));
 sg13g2_nor2_1 _21917_ (.A(net8707),
    .B(_12913_),
    .Y(_12914_));
 sg13g2_o21ai_1 _21918_ (.B1(_12914_),
    .Y(_12915_),
    .A1(net8659),
    .A2(_12051_));
 sg13g2_a21oi_1 _21919_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[7] ),
    .A2(net8738),
    .Y(_12916_),
    .B1(net8634));
 sg13g2_nor2_1 _21920_ (.A(net8502),
    .B(_12916_),
    .Y(_12917_));
 sg13g2_a22oi_1 _21921_ (.Y(_12918_),
    .B1(_12915_),
    .B2(_12917_),
    .A2(net8378),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[7] ));
 sg13g2_a21oi_2 _21922_ (.B1(_12909_),
    .Y(_12919_),
    .A2(net7606),
    .A1(net8573));
 sg13g2_nand2_1 _21923_ (.Y(_12920_),
    .A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[5] ),
    .B(net8838));
 sg13g2_a21oi_2 _21924_ (.B1(net8698),
    .Y(_12921_),
    .A2(net8703),
    .A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[5] ));
 sg13g2_o21ai_1 _21925_ (.B1(net8659),
    .Y(_12922_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[5] ),
    .A2(net8690));
 sg13g2_a21oi_1 _21926_ (.A1(_12920_),
    .A2(_12921_),
    .Y(_12923_),
    .B1(_12922_));
 sg13g2_nor2_1 _21927_ (.A(net8706),
    .B(_12923_),
    .Y(_12924_));
 sg13g2_o21ai_1 _21928_ (.B1(_12924_),
    .Y(_12925_),
    .A1(net8659),
    .A2(_12338_));
 sg13g2_a21oi_1 _21929_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[5] ),
    .A2(net8733),
    .Y(_12926_),
    .B1(net8630));
 sg13g2_nor2_1 _21930_ (.A(net8501),
    .B(_12926_),
    .Y(_12927_));
 sg13g2_a22oi_1 _21931_ (.Y(_12928_),
    .B1(_12925_),
    .B2(_12927_),
    .A2(net8376),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[5] ));
 sg13g2_nor2_1 _21932_ (.A(\soc_I.PC[5] ),
    .B(net8576),
    .Y(_12929_));
 sg13g2_a21oi_2 _21933_ (.B1(_12929_),
    .Y(_12930_),
    .A2(_12928_),
    .A1(net8576));
 sg13g2_nand2_1 _21934_ (.Y(_12931_),
    .A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[6] ),
    .B(net8838));
 sg13g2_a21oi_2 _21935_ (.B1(net8700),
    .Y(_12932_),
    .A2(net8705),
    .A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[6] ));
 sg13g2_o21ai_1 _21936_ (.B1(net8658),
    .Y(_12933_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[6] ),
    .A2(net8691));
 sg13g2_a21oi_1 _21937_ (.A1(_12931_),
    .A2(_12932_),
    .Y(_12934_),
    .B1(_12933_));
 sg13g2_nor2_1 _21938_ (.A(net8706),
    .B(_12934_),
    .Y(_12935_));
 sg13g2_o21ai_1 _21939_ (.B1(_12935_),
    .Y(_12936_),
    .A1(net8657),
    .A2(_11893_));
 sg13g2_a21oi_1 _21940_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[6] ),
    .A2(net8733),
    .Y(_12937_),
    .B1(net8631));
 sg13g2_nor2_1 _21941_ (.A(net8501),
    .B(_12937_),
    .Y(_12938_));
 sg13g2_a22oi_1 _21942_ (.Y(_12939_),
    .B1(_12936_),
    .B2(_12938_),
    .A2(net8376),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[6] ));
 sg13g2_nor2_1 _21943_ (.A(\soc_I.PC[6] ),
    .B(net8576),
    .Y(_12940_));
 sg13g2_a21oi_2 _21944_ (.B1(_12940_),
    .Y(_12941_),
    .A2(net7596),
    .A1(net8576));
 sg13g2_nor3_1 _21945_ (.A(_12919_),
    .B(_12930_),
    .C(_12941_),
    .Y(_12942_));
 sg13g2_nand2_1 _21946_ (.Y(_12943_),
    .A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[4] ),
    .B(net8838));
 sg13g2_a21oi_2 _21947_ (.B1(net8698),
    .Y(_12944_),
    .A2(net8703),
    .A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[4] ));
 sg13g2_o21ai_1 _21948_ (.B1(net8659),
    .Y(_12945_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[4] ),
    .A2(net8691));
 sg13g2_a21oi_1 _21949_ (.A1(_12943_),
    .A2(_12944_),
    .Y(_12946_),
    .B1(_12945_));
 sg13g2_nor2_1 _21950_ (.A(net8706),
    .B(_12946_),
    .Y(_12947_));
 sg13g2_o21ai_1 _21951_ (.B1(_12947_),
    .Y(_12948_),
    .A1(net8659),
    .A2(_12416_));
 sg13g2_a21oi_1 _21952_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[4] ),
    .A2(net8735),
    .Y(_12949_),
    .B1(net8630));
 sg13g2_nor2_1 _21953_ (.A(net8501),
    .B(_12949_),
    .Y(_12950_));
 sg13g2_a22oi_1 _21954_ (.Y(_12951_),
    .B1(_12948_),
    .B2(_12950_),
    .A2(net8376),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[4] ));
 sg13g2_nor2_1 _21955_ (.A(\soc_I.PC[4] ),
    .B(net8576),
    .Y(_12952_));
 sg13g2_a21oi_2 _21956_ (.B1(_12952_),
    .Y(_12953_),
    .A2(net7591),
    .A1(net8576));
 sg13g2_nor4_2 _21957_ (.A(_12919_),
    .B(_12930_),
    .C(_12941_),
    .Y(_12954_),
    .D(_12953_));
 sg13g2_nand3_1 _21958_ (.B(_12908_),
    .C(_12954_),
    .A(net7470),
    .Y(_12955_));
 sg13g2_nand2_1 _21959_ (.Y(_12956_),
    .A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[14] ),
    .B(net8836));
 sg13g2_a21oi_1 _21960_ (.A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[14] ),
    .A2(net8701),
    .Y(_12957_),
    .B1(net8696));
 sg13g2_o21ai_1 _21961_ (.B1(net8661),
    .Y(_12958_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[14] ),
    .A2(net8692));
 sg13g2_a21oi_1 _21962_ (.A1(_12956_),
    .A2(_12957_),
    .Y(_12959_),
    .B1(_12958_));
 sg13g2_nor2_1 _21963_ (.A(net8708),
    .B(_12959_),
    .Y(_12960_));
 sg13g2_o21ai_1 _21964_ (.B1(_12960_),
    .Y(_12961_),
    .A1(net8656),
    .A2(_12273_));
 sg13g2_a21oi_1 _21965_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[14] ),
    .A2(net8738),
    .Y(_12962_),
    .B1(net8628));
 sg13g2_nor2_1 _21966_ (.A(net8500),
    .B(_12962_),
    .Y(_12963_));
 sg13g2_a22oi_1 _21967_ (.Y(_12964_),
    .B1(_12961_),
    .B2(_12963_),
    .A2(net8374),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[14] ));
 sg13g2_nor2_1 _21968_ (.A(\soc_I.PC[14] ),
    .B(net8572),
    .Y(_12965_));
 sg13g2_a21oi_1 _21969_ (.A1(net8572),
    .A2(net7582),
    .Y(_12966_),
    .B1(_12965_));
 sg13g2_a21o_1 _21970_ (.A2(net7582),
    .A1(net8572),
    .B1(_12965_),
    .X(_12967_));
 sg13g2_a21o_1 _21971_ (.A2(net8703),
    .A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[9] ),
    .B1(net8698),
    .X(_12968_));
 sg13g2_a21oi_1 _21972_ (.A1(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[9] ),
    .A2(net8838),
    .Y(_12969_),
    .B1(_12968_));
 sg13g2_o21ai_1 _21973_ (.B1(net8657),
    .Y(_12970_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[9] ),
    .A2(net8691));
 sg13g2_o21ai_1 _21974_ (.B1(net8630),
    .Y(_12971_),
    .A1(_12969_),
    .A2(_12970_));
 sg13g2_a21o_1 _21975_ (.A2(_12360_),
    .A1(net8655),
    .B1(_12971_),
    .X(_12972_));
 sg13g2_a21oi_1 _21976_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[9] ),
    .A2(net8733),
    .Y(_12973_),
    .B1(net8630));
 sg13g2_nor2_1 _21977_ (.A(net8501),
    .B(_12973_),
    .Y(_12974_));
 sg13g2_a22oi_1 _21978_ (.Y(_12975_),
    .B1(_12972_),
    .B2(_12974_),
    .A2(net8376),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[9] ));
 sg13g2_nor2_1 _21979_ (.A(\soc_I.PC[9] ),
    .B(net8575),
    .Y(_12976_));
 sg13g2_a21oi_2 _21980_ (.B1(_12976_),
    .Y(_12977_),
    .A2(net7579),
    .A1(net8575));
 sg13g2_nor2_1 _21981_ (.A(\soc_I.PC[11] ),
    .B(net8573),
    .Y(_12978_));
 sg13g2_a21o_1 _21982_ (.A2(net8702),
    .A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[11] ),
    .B1(net8697),
    .X(_12979_));
 sg13g2_a21oi_1 _21983_ (.A1(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[11] ),
    .A2(net8837),
    .Y(_12980_),
    .B1(_12979_));
 sg13g2_o21ai_1 _21984_ (.B1(net8659),
    .Y(_12981_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[11] ),
    .A2(net8690));
 sg13g2_o21ai_1 _21985_ (.B1(net8629),
    .Y(_12982_),
    .A1(_12980_),
    .A2(_12981_));
 sg13g2_a21o_1 _21986_ (.A2(_12026_),
    .A1(net8655),
    .B1(_12982_),
    .X(_12983_));
 sg13g2_a21oi_1 _21987_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[11] ),
    .A2(net8731),
    .Y(_12984_),
    .B1(net8629));
 sg13g2_nor2_1 _21988_ (.A(net8500),
    .B(_12984_),
    .Y(_12985_));
 sg13g2_a22oi_1 _21989_ (.Y(_12986_),
    .B1(_12983_),
    .B2(_12985_),
    .A2(_11760_),
    .A1(net2736));
 sg13g2_a21oi_2 _21990_ (.B1(_12978_),
    .Y(_12987_),
    .A2(net7573),
    .A1(net8573));
 sg13g2_nor2_1 _21991_ (.A(\soc_I.PC[15] ),
    .B(net8573),
    .Y(_12988_));
 sg13g2_nand2_1 _21992_ (.Y(_12989_),
    .A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[15] ),
    .B(net8836));
 sg13g2_a21oi_1 _21993_ (.A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[15] ),
    .A2(net8701),
    .Y(_12990_),
    .B1(net8696));
 sg13g2_o21ai_1 _21994_ (.B1(net8656),
    .Y(_12991_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[15] ),
    .A2(net8690));
 sg13g2_a21oi_1 _21995_ (.A1(_12989_),
    .A2(_12990_),
    .Y(_12992_),
    .B1(_12991_));
 sg13g2_nor2_1 _21996_ (.A(net8708),
    .B(_12992_),
    .Y(_12993_));
 sg13g2_o21ai_1 _21997_ (.B1(_12993_),
    .Y(_12994_),
    .A1(net8664),
    .A2(_12252_));
 sg13g2_a21oi_1 _21998_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[15] ),
    .A2(net8731),
    .Y(_12995_),
    .B1(net8629));
 sg13g2_nor2_1 _21999_ (.A(net8499),
    .B(_12995_),
    .Y(_12996_));
 sg13g2_a22oi_1 _22000_ (.Y(_12997_),
    .B1(_12994_),
    .B2(_12996_),
    .A2(net8374),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[15] ));
 sg13g2_a21oi_2 _22001_ (.B1(_12988_),
    .Y(_12998_),
    .A2(net7567),
    .A1(net8573));
 sg13g2_nor2_1 _22002_ (.A(\soc_I.PC[8] ),
    .B(net8574),
    .Y(_12999_));
 sg13g2_a21o_1 _22003_ (.A2(net8703),
    .A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[8] ),
    .B1(net8698),
    .X(_13000_));
 sg13g2_a21oi_1 _22004_ (.A1(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[8] ),
    .A2(net8841),
    .Y(_13001_),
    .B1(_13000_));
 sg13g2_o21ai_1 _22005_ (.B1(net8658),
    .Y(_13002_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[8] ),
    .A2(net8695));
 sg13g2_o21ai_1 _22006_ (.B1(net8630),
    .Y(_13003_),
    .A1(_13001_),
    .A2(_13002_));
 sg13g2_a21o_1 _22007_ (.A2(_11914_),
    .A1(net8655),
    .B1(_13003_),
    .X(_13004_));
 sg13g2_a21oi_1 _22008_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[8] ),
    .A2(net8733),
    .Y(_13005_),
    .B1(net8630));
 sg13g2_nor2_1 _22009_ (.A(net8501),
    .B(_13005_),
    .Y(_13006_));
 sg13g2_a22oi_1 _22010_ (.Y(_13007_),
    .B1(_13004_),
    .B2(_13006_),
    .A2(net8376),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[8] ));
 sg13g2_a21oi_2 _22011_ (.B1(_12999_),
    .Y(_13008_),
    .A2(_13007_),
    .A1(net8574));
 sg13g2_nor2_1 _22012_ (.A(\soc_I.PC[13] ),
    .B(net8574),
    .Y(_13009_));
 sg13g2_nand2_1 _22013_ (.Y(_13010_),
    .A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[13] ),
    .B(net8838));
 sg13g2_a21oi_1 _22014_ (.A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[13] ),
    .A2(net8703),
    .Y(_13011_),
    .B1(net8698));
 sg13g2_o21ai_1 _22015_ (.B1(net8657),
    .Y(_13012_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[13] ),
    .A2(net8691));
 sg13g2_a21oi_1 _22016_ (.A1(_13010_),
    .A2(_13011_),
    .Y(_13013_),
    .B1(_13012_));
 sg13g2_nor2_1 _22017_ (.A(net8706),
    .B(_13013_),
    .Y(_13014_));
 sg13g2_o21ai_1 _22018_ (.B1(_13014_),
    .Y(_13015_),
    .A1(net8657),
    .A2(_12450_));
 sg13g2_a21oi_1 _22019_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[13] ),
    .A2(net8733),
    .Y(_13016_),
    .B1(net8630));
 sg13g2_nor2_1 _22020_ (.A(net8501),
    .B(_13016_),
    .Y(_13017_));
 sg13g2_a22oi_1 _22021_ (.Y(_13018_),
    .B1(_13015_),
    .B2(_13017_),
    .A2(net8376),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[13] ));
 sg13g2_a21oi_2 _22022_ (.B1(_13009_),
    .Y(_13019_),
    .A2(net7556),
    .A1(_10859_));
 sg13g2_nor2_1 _22023_ (.A(\soc_I.PC[10] ),
    .B(net8574),
    .Y(_13020_));
 sg13g2_nand2_1 _22024_ (.Y(_13021_),
    .A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[10] ),
    .B(net8838));
 sg13g2_a21oi_2 _22025_ (.B1(net8698),
    .Y(_13022_),
    .A2(net8703),
    .A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[10] ));
 sg13g2_o21ai_1 _22026_ (.B1(net8658),
    .Y(_13023_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[10] ),
    .A2(net8691));
 sg13g2_a21oi_1 _22027_ (.A1(_13021_),
    .A2(_13022_),
    .Y(_13024_),
    .B1(_13023_));
 sg13g2_nor2_1 _22028_ (.A(net8706),
    .B(_13024_),
    .Y(_13025_));
 sg13g2_o21ai_1 _22029_ (.B1(_13025_),
    .Y(_13026_),
    .A1(net8657),
    .A2(_12068_));
 sg13g2_a21oi_1 _22030_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[10] ),
    .A2(net8733),
    .Y(_13027_),
    .B1(net8631));
 sg13g2_nor2_1 _22031_ (.A(net8502),
    .B(_13027_),
    .Y(_13028_));
 sg13g2_a22oi_1 _22032_ (.Y(_13029_),
    .B1(_13026_),
    .B2(_13028_),
    .A2(net8378),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[10] ));
 sg13g2_a21oi_2 _22033_ (.B1(_13020_),
    .Y(_13030_),
    .A2(_13029_),
    .A1(net8574));
 sg13g2_nand2_1 _22034_ (.Y(_13031_),
    .A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[12] ),
    .B(net8838));
 sg13g2_a21oi_1 _22035_ (.A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[12] ),
    .A2(net8705),
    .Y(_13032_),
    .B1(net8700));
 sg13g2_o21ai_1 _22036_ (.B1(net8658),
    .Y(_13033_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[12] ),
    .A2(net8691));
 sg13g2_a21oi_1 _22037_ (.A1(_13031_),
    .A2(_13032_),
    .Y(_13034_),
    .B1(_13033_));
 sg13g2_nor2_1 _22038_ (.A(net8706),
    .B(_13034_),
    .Y(_13035_));
 sg13g2_o21ai_1 _22039_ (.B1(_13035_),
    .Y(_13036_),
    .A1(net8657),
    .A2(_12438_));
 sg13g2_a21oi_1 _22040_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[12] ),
    .A2(net8733),
    .Y(_13037_),
    .B1(net8631));
 sg13g2_nor2_1 _22041_ (.A(net8501),
    .B(_13037_),
    .Y(_13038_));
 sg13g2_a22oi_1 _22042_ (.Y(_13039_),
    .B1(_13036_),
    .B2(_13038_),
    .A2(net8376),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[12] ));
 sg13g2_nor2_1 _22043_ (.A(\soc_I.PC[12] ),
    .B(net8574),
    .Y(_13040_));
 sg13g2_a21oi_2 _22044_ (.B1(_13040_),
    .Y(_13041_),
    .A2(net7545),
    .A1(net8574));
 sg13g2_nor3_1 _22045_ (.A(_12998_),
    .B(_13019_),
    .C(_13041_),
    .Y(_13042_));
 sg13g2_nor4_2 _22046_ (.A(_12977_),
    .B(_12987_),
    .C(_13008_),
    .Y(_13043_),
    .D(_13030_));
 sg13g2_and3_2 _22047_ (.X(_13044_),
    .A(_12967_),
    .B(_13042_),
    .C(_13043_));
 sg13g2_nand4_1 _22048_ (.B(_12967_),
    .C(_13042_),
    .A(_12954_),
    .Y(_13045_),
    .D(_13043_));
 sg13g2_nor4_2 _22049_ (.A(\soc_I.clint_I.addr[0] ),
    .B(\soc_I.clint_I.addr[1] ),
    .C(_12907_),
    .Y(_13046_),
    .D(_13045_));
 sg13g2_nand4_1 _22050_ (.B(_12908_),
    .C(_12954_),
    .A(_12883_),
    .Y(_13047_),
    .D(_13044_));
 sg13g2_nor2_1 _22051_ (.A(_12895_),
    .B(_12906_),
    .Y(_13048_));
 sg13g2_and2_2 _22052_ (.A(_12954_),
    .B(_13048_),
    .X(_13049_));
 sg13g2_nand2_2 _22053_ (.Y(_13050_),
    .A(net7470),
    .B(_13049_));
 sg13g2_nand3_1 _22054_ (.B(_13044_),
    .C(_13049_),
    .A(net7470),
    .Y(_13051_));
 sg13g2_nand3_1 _22055_ (.B(_13044_),
    .C(_13049_),
    .A(net7470),
    .Y(_13052_));
 sg13g2_and2_1 _22056_ (.A(_13047_),
    .B(_13051_),
    .X(_13053_));
 sg13g2_nand2_1 _22057_ (.Y(_13054_),
    .A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[17] ),
    .B(net8836));
 sg13g2_a21oi_1 _22058_ (.A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[17] ),
    .A2(net8701),
    .Y(_13055_),
    .B1(net8696));
 sg13g2_o21ai_1 _22059_ (.B1(net8662),
    .Y(_13056_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[17] ),
    .A2(net8690));
 sg13g2_a21oi_1 _22060_ (.A1(_13054_),
    .A2(_13055_),
    .Y(_13057_),
    .B1(_13056_));
 sg13g2_nor2_1 _22061_ (.A(net8708),
    .B(_13057_),
    .Y(_13058_));
 sg13g2_o21ai_1 _22062_ (.B1(_13058_),
    .Y(_13059_),
    .A1(net8656),
    .A2(_12349_));
 sg13g2_a21oi_1 _22063_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[17] ),
    .A2(net8730),
    .Y(_13060_),
    .B1(net8627));
 sg13g2_nor2_1 _22064_ (.A(net8499),
    .B(_13060_),
    .Y(_13061_));
 sg13g2_a22oi_1 _22065_ (.Y(_13062_),
    .B1(_13059_),
    .B2(_13061_),
    .A2(net8374),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[17] ));
 sg13g2_nor2_1 _22066_ (.A(\led[1] ),
    .B(net8570),
    .Y(_13063_));
 sg13g2_a21oi_1 _22067_ (.A1(net8570),
    .A2(net7539),
    .Y(_13064_),
    .B1(_13063_));
 sg13g2_nand2_1 _22068_ (.Y(_13065_),
    .A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[18] ),
    .B(net8836));
 sg13g2_a21oi_1 _22069_ (.A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[18] ),
    .A2(net8701),
    .Y(_13066_),
    .B1(net8696));
 sg13g2_o21ai_1 _22070_ (.B1(net8662),
    .Y(_13067_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[18] ),
    .A2(net8694));
 sg13g2_a21oi_1 _22071_ (.A1(_13065_),
    .A2(_13066_),
    .Y(_13068_),
    .B1(_13067_));
 sg13g2_nor2_1 _22072_ (.A(net8708),
    .B(_13068_),
    .Y(_13069_));
 sg13g2_o21ai_1 _22073_ (.B1(_13069_),
    .Y(_13070_),
    .A1(net8656),
    .A2(_12285_));
 sg13g2_a21oi_1 _22074_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[18] ),
    .A2(net8730),
    .Y(_13071_),
    .B1(net8627));
 sg13g2_nor2_1 _22075_ (.A(net8499),
    .B(_13071_),
    .Y(_13072_));
 sg13g2_a22oi_1 _22076_ (.Y(_13073_),
    .B1(_13070_),
    .B2(_13072_),
    .A2(net8374),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[18] ));
 sg13g2_nor2_1 _22077_ (.A(\led[2] ),
    .B(net8570),
    .Y(_13074_));
 sg13g2_a21oi_1 _22078_ (.A1(net8570),
    .A2(net7533),
    .Y(_13075_),
    .B1(_13074_));
 sg13g2_nand2_1 _22079_ (.Y(_13076_),
    .A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[16] ),
    .B(net8836));
 sg13g2_a21oi_1 _22080_ (.A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[16] ),
    .A2(net8701),
    .Y(_13077_),
    .B1(net8696));
 sg13g2_o21ai_1 _22081_ (.B1(net8656),
    .Y(_13078_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[16] ),
    .A2(net8690));
 sg13g2_a21oi_1 _22082_ (.A1(_13076_),
    .A2(_13077_),
    .Y(_13079_),
    .B1(_13078_));
 sg13g2_nor2_1 _22083_ (.A(net8708),
    .B(_13079_),
    .Y(_13080_));
 sg13g2_o21ai_1 _22084_ (.B1(_13080_),
    .Y(_13081_),
    .A1(net8656),
    .A2(_12427_));
 sg13g2_a21oi_1 _22085_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[16] ),
    .A2(net8730),
    .Y(_13082_),
    .B1(net8627));
 sg13g2_nor2_1 _22086_ (.A(net8499),
    .B(_13082_),
    .Y(_13083_));
 sg13g2_a22oi_1 _22087_ (.Y(_13084_),
    .B1(_13081_),
    .B2(_13083_),
    .A2(net8374),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[16] ));
 sg13g2_nor2_1 _22088_ (.A(\led[0] ),
    .B(net8571),
    .Y(_13085_));
 sg13g2_a21oi_1 _22089_ (.A1(net8570),
    .A2(net7527),
    .Y(_13086_),
    .B1(_13085_));
 sg13g2_nand2_1 _22090_ (.Y(_13087_),
    .A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[19] ),
    .B(net8836));
 sg13g2_a21oi_1 _22091_ (.A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[19] ),
    .A2(net8702),
    .Y(_13088_),
    .B1(net8697));
 sg13g2_o21ai_1 _22092_ (.B1(net8661),
    .Y(_13089_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[19] ),
    .A2(net8694));
 sg13g2_a21oi_1 _22093_ (.A1(_13087_),
    .A2(_13088_),
    .Y(_13090_),
    .B1(_13089_));
 sg13g2_nor2_1 _22094_ (.A(net8708),
    .B(_13090_),
    .Y(_13091_));
 sg13g2_o21ai_1 _22095_ (.B1(_13091_),
    .Y(_13092_),
    .A1(net8656),
    .A2(_12389_));
 sg13g2_a21oi_1 _22096_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[19] ),
    .A2(net8731),
    .Y(_13093_),
    .B1(net8627));
 sg13g2_nor2_1 _22097_ (.A(net8499),
    .B(_13093_),
    .Y(_13094_));
 sg13g2_a22oi_1 _22098_ (.Y(_13095_),
    .B1(_13092_),
    .B2(_13094_),
    .A2(net8375),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[19] ));
 sg13g2_nor2_1 _22099_ (.A(\led[3] ),
    .B(net8572),
    .Y(_13096_));
 sg13g2_a21oi_1 _22100_ (.A1(net8572),
    .A2(_13095_),
    .Y(_13097_),
    .B1(_13096_));
 sg13g2_nor4_2 _22101_ (.A(_13064_),
    .B(_13075_),
    .C(_13086_),
    .Y(_13098_),
    .D(_13097_));
 sg13g2_nor2_1 _22102_ (.A(\soc_I.PC[21] ),
    .B(net8577),
    .Y(_13099_));
 sg13g2_nand2_1 _22103_ (.Y(_13100_),
    .A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[21] ),
    .B(net8840));
 sg13g2_a21oi_1 _22104_ (.A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[21] ),
    .A2(net8704),
    .Y(_13101_),
    .B1(net8699));
 sg13g2_o21ai_1 _22105_ (.B1(net8660),
    .Y(_13102_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[21] ),
    .A2(net8693));
 sg13g2_a21oi_1 _22106_ (.A1(_13100_),
    .A2(_13101_),
    .Y(_13103_),
    .B1(_13102_));
 sg13g2_nor2_1 _22107_ (.A(net8707),
    .B(_13103_),
    .Y(_13104_));
 sg13g2_o21ai_1 _22108_ (.B1(_13104_),
    .Y(_13105_),
    .A1(net8661),
    .A2(_12399_));
 sg13g2_a21oi_1 _22109_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[21] ),
    .A2(net8736),
    .Y(_13106_),
    .B1(net8633));
 sg13g2_nor2_1 _22110_ (.A(net8503),
    .B(_13106_),
    .Y(_13107_));
 sg13g2_a22oi_1 _22111_ (.Y(_13108_),
    .B1(_13105_),
    .B2(_13107_),
    .A2(net8377),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[21] ));
 sg13g2_a21oi_2 _22112_ (.B1(_13099_),
    .Y(_13109_),
    .A2(net7515),
    .A1(net8577));
 sg13g2_nor2_1 _22113_ (.A(\soc_I.PC[20] ),
    .B(net8571),
    .Y(_13110_));
 sg13g2_nand2_1 _22114_ (.Y(_13111_),
    .A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[20] ),
    .B(net8840));
 sg13g2_a21oi_1 _22115_ (.A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[20] ),
    .A2(net8704),
    .Y(_13112_),
    .B1(net8699));
 sg13g2_o21ai_1 _22116_ (.B1(net8660),
    .Y(_13113_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[20] ),
    .A2(net8692));
 sg13g2_a21oi_1 _22117_ (.A1(_13111_),
    .A2(_13112_),
    .Y(_13114_),
    .B1(_13113_));
 sg13g2_nor2_1 _22118_ (.A(net8707),
    .B(_13114_),
    .Y(_13115_));
 sg13g2_o21ai_1 _22119_ (.B1(_13115_),
    .Y(_13116_),
    .A1(net8661),
    .A2(_12179_));
 sg13g2_a21oi_1 _22120_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[20] ),
    .A2(net8737),
    .Y(_13117_),
    .B1(net8633));
 sg13g2_nor2_1 _22121_ (.A(net8503),
    .B(_13117_),
    .Y(_13118_));
 sg13g2_a22oi_1 _22122_ (.Y(_13119_),
    .B1(_13116_),
    .B2(_13118_),
    .A2(net8378),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[20] ));
 sg13g2_a21oi_1 _22123_ (.A1(net8571),
    .A2(net7510),
    .Y(_13120_),
    .B1(_13110_));
 sg13g2_a21o_1 _22124_ (.A2(net7510),
    .A1(net8571),
    .B1(_13110_),
    .X(_13121_));
 sg13g2_nor2_1 _22125_ (.A(_13109_),
    .B(_13121_),
    .Y(_13122_));
 sg13g2_and3_2 _22126_ (.X(_13123_),
    .A(_12467_),
    .B(_13098_),
    .C(_13122_));
 sg13g2_nand2_1 _22127_ (.Y(_13124_),
    .A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[23] ),
    .B(net8839));
 sg13g2_a21oi_1 _22128_ (.A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[23] ),
    .A2(net8704),
    .Y(_13125_),
    .B1(net8699));
 sg13g2_o21ai_1 _22129_ (.B1(net8660),
    .Y(_13126_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[23] ),
    .A2(net8692));
 sg13g2_a21oi_2 _22130_ (.B1(_13126_),
    .Y(_13127_),
    .A2(_13125_),
    .A1(_13124_));
 sg13g2_nor2_2 _22131_ (.A(net8708),
    .B(_13127_),
    .Y(_13128_));
 sg13g2_o21ai_1 _22132_ (.B1(_13128_),
    .Y(_13129_),
    .A1(net8656),
    .A2(_12320_));
 sg13g2_a21oi_1 _22133_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[23] ),
    .A2(net8730),
    .Y(_13130_),
    .B1(net8627));
 sg13g2_nor2_1 _22134_ (.A(net8499),
    .B(_13130_),
    .Y(_13131_));
 sg13g2_a22oi_1 _22135_ (.Y(_13132_),
    .B1(_13129_),
    .B2(_13131_),
    .A2(net8374),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[23] ));
 sg13g2_nor2_2 _22136_ (.A(\soc_I.PC[23] ),
    .B(net8575),
    .Y(_13133_));
 sg13g2_a21oi_2 _22137_ (.B1(_13133_),
    .Y(_13134_),
    .A2(net7503),
    .A1(net8570));
 sg13g2_inv_1 _22138_ (.Y(_13135_),
    .A(_13134_));
 sg13g2_nor2_1 _22139_ (.A(\soc_I.PC[22] ),
    .B(net8577),
    .Y(_13136_));
 sg13g2_nand2_1 _22140_ (.Y(_13137_),
    .A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[22] ),
    .B(net8840));
 sg13g2_a21oi_1 _22141_ (.A1(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[22] ),
    .A2(net8705),
    .Y(_13138_),
    .B1(net8700));
 sg13g2_o21ai_1 _22142_ (.B1(net8660),
    .Y(_13139_),
    .A1(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[22] ),
    .A2(net8692));
 sg13g2_a21oi_1 _22143_ (.A1(_13137_),
    .A2(_13138_),
    .Y(_13140_),
    .B1(_13139_));
 sg13g2_nor2_1 _22144_ (.A(net8707),
    .B(_13140_),
    .Y(_13141_));
 sg13g2_o21ai_1 _22145_ (.B1(_13141_),
    .Y(_13142_),
    .A1(net8662),
    .A2(_12263_));
 sg13g2_a21oi_1 _22146_ (.A1(\soc_I.kianv_I.datapath_unit_I.DataLatched[22] ),
    .A2(net8736),
    .Y(_13143_),
    .B1(net8633));
 sg13g2_nor2_1 _22147_ (.A(net8503),
    .B(_13143_),
    .Y(_13144_));
 sg13g2_a22oi_1 _22148_ (.Y(_13145_),
    .B1(_13142_),
    .B2(_13144_),
    .A2(net8377),
    .A1(\soc_I.kianv_I.datapath_unit_I.ALUOut[22] ));
 sg13g2_a21oi_2 _22149_ (.B1(_13136_),
    .Y(_13146_),
    .A2(_13145_),
    .A1(net8577));
 sg13g2_nand2b_2 _22150_ (.Y(_13147_),
    .B(_13146_),
    .A_N(_13134_));
 sg13g2_and4_1 _22151_ (.A(_12521_),
    .B(_12531_),
    .C(_12540_),
    .D(_12549_),
    .X(_13148_));
 sg13g2_nand4_1 _22152_ (.B(_12531_),
    .C(_12540_),
    .A(_12521_),
    .Y(_13149_),
    .D(_12549_));
 sg13g2_nor2_2 _22153_ (.A(_12500_),
    .B(_13149_),
    .Y(_13150_));
 sg13g2_nand2_2 _22154_ (.Y(_13151_),
    .A(_12511_),
    .B(_13150_));
 sg13g2_nor2_1 _22155_ (.A(_13147_),
    .B(_13151_),
    .Y(_13152_));
 sg13g2_nand2_1 _22156_ (.Y(_13153_),
    .A(_13123_),
    .B(_13152_));
 sg13g2_nor3_2 _22157_ (.A(net8960),
    .B(_13053_),
    .C(_13153_),
    .Y(_13154_));
 sg13g2_and2_2 _22158_ (.A(_12942_),
    .B(_12953_),
    .X(_13155_));
 sg13g2_and4_1 _22159_ (.A(_12883_),
    .B(_12908_),
    .C(_13044_),
    .D(_13155_),
    .X(_13156_));
 sg13g2_nand4_1 _22160_ (.B(_12908_),
    .C(_13044_),
    .A(net7470),
    .Y(_13157_),
    .D(_13155_));
 sg13g2_nor4_2 _22161_ (.A(_13109_),
    .B(_13120_),
    .C(_13134_),
    .Y(_13158_),
    .D(_13146_));
 sg13g2_and2_1 _22162_ (.A(_13098_),
    .B(_13158_),
    .X(_13159_));
 sg13g2_nand2_2 _22163_ (.Y(_13160_),
    .A(_13098_),
    .B(_13158_));
 sg13g2_nand3_1 _22164_ (.B(_13098_),
    .C(_13158_),
    .A(net7480),
    .Y(_13161_));
 sg13g2_nor2_2 _22165_ (.A(_13151_),
    .B(_13161_),
    .Y(_13162_));
 sg13g2_nand3_1 _22166_ (.B(_13156_),
    .C(_13162_),
    .A(net8999),
    .Y(_13163_));
 sg13g2_nor3_1 _22167_ (.A(\soc_I.uart_lsr_rdy ),
    .B(net8666),
    .C(\soc_I.clint_I.addr[1] ),
    .Y(_13164_));
 sg13g2_and3_1 _22168_ (.X(_13165_),
    .A(\soc_I.clint_I.addr[0] ),
    .B(_13044_),
    .C(_13164_));
 sg13g2_nand3_1 _22169_ (.B(_13162_),
    .C(_13165_),
    .A(_13049_),
    .Y(_13166_));
 sg13g2_nand3b_1 _22170_ (.B(_13163_),
    .C(_13166_),
    .Y(_13167_),
    .A_N(_13154_));
 sg13g2_nand2_2 _22171_ (.Y(_13168_),
    .A(_13046_),
    .B(_13162_));
 sg13g2_nor2_2 _22172_ (.A(net9250),
    .B(_13168_),
    .Y(_13169_));
 sg13g2_nor3_2 _22173_ (.A(net5561),
    .B(_13153_),
    .C(_13157_),
    .Y(_13170_));
 sg13g2_nor2_1 _22174_ (.A(net9244),
    .B(_13168_),
    .Y(_13171_));
 sg13g2_nor4_1 _22175_ (.A(_13167_),
    .B(_13169_),
    .C(_13170_),
    .D(_13171_),
    .Y(_13172_));
 sg13g2_nor2_2 _22176_ (.A(net4970),
    .B(net7479),
    .Y(_13173_));
 sg13g2_nand3_1 _22177_ (.B(_13109_),
    .C(_13121_),
    .A(_13098_),
    .Y(_13174_));
 sg13g2_nor3_2 _22178_ (.A(_13147_),
    .B(_13151_),
    .C(_13174_),
    .Y(_13175_));
 sg13g2_nor2b_2 _22179_ (.A(_13051_),
    .B_N(_13175_),
    .Y(_13176_));
 sg13g2_and2_2 _22180_ (.A(_13046_),
    .B(_13175_),
    .X(_13177_));
 sg13g2_nand2_2 _22181_ (.Y(_13178_),
    .A(_12883_),
    .B(_12906_));
 sg13g2_nor3_1 _22182_ (.A(net7493),
    .B(_13045_),
    .C(_13178_),
    .Y(_13179_));
 sg13g2_and2_2 _22183_ (.A(_13175_),
    .B(_13179_),
    .X(_13180_));
 sg13g2_nor3_1 _22184_ (.A(_13176_),
    .B(_13177_),
    .C(_13180_),
    .Y(_13181_));
 sg13g2_nand2b_2 _22185_ (.Y(_13182_),
    .B(_13173_),
    .A_N(_13181_));
 sg13g2_nand3_1 _22186_ (.B(_13042_),
    .C(_13043_),
    .A(_12966_),
    .Y(_13183_));
 sg13g2_nand2_1 _22187_ (.Y(_13184_),
    .A(_12510_),
    .B(_13150_));
 sg13g2_nor2_1 _22188_ (.A(_13160_),
    .B(_13184_),
    .Y(_13185_));
 sg13g2_nor3_2 _22189_ (.A(_13160_),
    .B(_13183_),
    .C(_13184_),
    .Y(_13186_));
 sg13g2_nand2b_2 _22190_ (.Y(_13187_),
    .B(_13186_),
    .A_N(_13050_));
 sg13g2_nand2b_1 _22191_ (.Y(_13188_),
    .B(_13186_),
    .A_N(_12955_));
 sg13g2_nand4_1 _22192_ (.B(_12930_),
    .C(_12941_),
    .A(_12919_),
    .Y(_13189_),
    .D(_12953_));
 sg13g2_nand4_1 _22193_ (.B(_12977_),
    .C(_12987_),
    .A(_12967_),
    .Y(_13190_),
    .D(_12998_));
 sg13g2_nand4_1 _22194_ (.B(_13019_),
    .C(_13030_),
    .A(_13008_),
    .Y(_13191_),
    .D(_13041_));
 sg13g2_nor3_2 _22195_ (.A(_13189_),
    .B(_13190_),
    .C(_13191_),
    .Y(_13192_));
 sg13g2_nand4_1 _22196_ (.B(_12906_),
    .C(_13185_),
    .A(net7470),
    .Y(_13193_),
    .D(_13192_));
 sg13g2_nand2_1 _22197_ (.Y(_13194_),
    .A(_13046_),
    .B(_13185_));
 sg13g2_nand4_1 _22198_ (.B(net7425),
    .C(_13193_),
    .A(_13187_),
    .Y(_13195_),
    .D(_13194_));
 sg13g2_nand2_1 _22199_ (.Y(_13196_),
    .A(net7480),
    .B(_13195_));
 sg13g2_nand3_1 _22200_ (.B(_13182_),
    .C(_13196_),
    .A(_13172_),
    .Y(_13197_));
 sg13g2_nor4_1 _22201_ (.A(_12489_),
    .B(_12510_),
    .C(_13149_),
    .D(_13160_),
    .Y(_13198_));
 sg13g2_a21oi_1 _22202_ (.A1(_13046_),
    .A2(_13198_),
    .Y(_13199_),
    .B1(_13150_));
 sg13g2_a21oi_2 _22203_ (.B1(_13199_),
    .Y(_13200_),
    .A2(_13197_),
    .A1(_12882_));
 sg13g2_nand2b_1 _22204_ (.Y(_13201_),
    .B(_13200_),
    .A_N(net9266));
 sg13g2_nor2_2 _22205_ (.A(\soc_I.uart_lsr_rdy ),
    .B(_13201_),
    .Y(_13202_));
 sg13g2_nand2_1 _22206_ (.Y(_13203_),
    .A(_00108_),
    .B(_12895_));
 sg13g2_a21oi_1 _22207_ (.A1(_00109_),
    .A2(_12894_),
    .Y(_13204_),
    .B1(_12879_));
 sg13g2_and2_2 _22208_ (.A(\soc_I.gpio0_I.ready ),
    .B(_12879_),
    .X(_13205_));
 sg13g2_a221oi_1 _22209_ (.B2(\soc_I.gpio0_I.rdata[0] ),
    .C1(_12878_),
    .B1(_13205_),
    .A1(_13203_),
    .Y(_13206_),
    .A2(_13204_));
 sg13g2_nor2_1 _22210_ (.A(net9254),
    .B(_10604_),
    .Y(_13207_));
 sg13g2_a221oi_1 _22211_ (.B2(_00107_),
    .C1(_13206_),
    .B1(net8834),
    .A1(\soc_I.div_ready ),
    .Y(_13208_),
    .A2(_00106_));
 sg13g2_nand2_1 _22212_ (.Y(_13209_),
    .A(net8993),
    .B(_13208_));
 sg13g2_nor3_1 _22213_ (.A(_12489_),
    .B(_12499_),
    .C(_12511_),
    .Y(_13210_));
 sg13g2_and4_2 _22214_ (.A(_13098_),
    .B(_13148_),
    .C(_13158_),
    .D(_13210_),
    .X(_13211_));
 sg13g2_nand3_1 _22215_ (.B(_13159_),
    .C(_13210_),
    .A(_13148_),
    .Y(_13212_));
 sg13g2_nand2b_1 _22216_ (.Y(_13213_),
    .B(_13211_),
    .A_N(_13183_));
 sg13g2_nor2_1 _22217_ (.A(_12955_),
    .B(net7466),
    .Y(_13214_));
 sg13g2_nor2_1 _22218_ (.A(net7467),
    .B(net7465),
    .Y(_13215_));
 sg13g2_a221oi_1 _22219_ (.B2(_00111_),
    .C1(net8991),
    .B1(net7448),
    .A1(_00110_),
    .Y(_13216_),
    .A2(net7452));
 sg13g2_nand4_1 _22220_ (.B(_12998_),
    .C(_13019_),
    .A(_12967_),
    .Y(_13217_),
    .D(_13041_));
 sg13g2_nand4_1 _22221_ (.B(_12987_),
    .C(_13008_),
    .A(_12977_),
    .Y(_13218_),
    .D(_13030_));
 sg13g2_nor3_2 _22222_ (.A(_13189_),
    .B(_13217_),
    .C(_13218_),
    .Y(_13219_));
 sg13g2_and4_2 _22223_ (.A(net7470),
    .B(_12906_),
    .C(_13211_),
    .D(_13219_),
    .X(_13220_));
 sg13g2_nor2_1 _22224_ (.A(net7450),
    .B(net7445),
    .Y(_13221_));
 sg13g2_a21oi_1 _22225_ (.A1(_12955_),
    .A2(net7467),
    .Y(_13222_),
    .B1(net7466));
 sg13g2_nand2_2 _22226_ (.Y(_13223_),
    .A(_12895_),
    .B(_13220_));
 sg13g2_and2_2 _22227_ (.A(net7492),
    .B(_13220_),
    .X(_13224_));
 sg13g2_nor2_1 _22228_ (.A(net7468),
    .B(_13212_),
    .Y(_13225_));
 sg13g2_and4_2 _22229_ (.A(net7470),
    .B(_12906_),
    .C(_13211_),
    .D(_13219_),
    .X(_13226_));
 sg13g2_a21oi_2 _22230_ (.B1(_13226_),
    .Y(_13227_),
    .A2(_13225_),
    .A1(\soc_I.IRQ3 ));
 sg13g2_and2_1 _22231_ (.A(net7492),
    .B(_13226_),
    .X(_13228_));
 sg13g2_and2_2 _22232_ (.A(_12895_),
    .B(_13226_),
    .X(_13229_));
 sg13g2_nand2_1 _22233_ (.Y(_13230_),
    .A(_12895_),
    .B(_13226_));
 sg13g2_a221oi_1 _22234_ (.B2(_00302_),
    .C1(_13227_),
    .B1(_13229_),
    .A1(_00112_),
    .Y(_13231_),
    .A2(net7443));
 sg13g2_o21ai_1 _22235_ (.B1(_13216_),
    .Y(_13232_),
    .A1(_13222_),
    .A2(_13231_));
 sg13g2_a21oi_1 _22236_ (.A1(_13209_),
    .A2(_13232_),
    .Y(_13233_),
    .B1(net9250));
 sg13g2_nor2_1 _22237_ (.A(net9244),
    .B(_13233_),
    .Y(_13234_));
 sg13g2_nor2_1 _22238_ (.A(\soc_I.rx_uart_i.fifo_i.cnt[1] ),
    .B(net5574),
    .Y(_13235_));
 sg13g2_nor4_2 _22239_ (.A(\soc_I.rx_uart_i.fifo_i.cnt[1] ),
    .B(\soc_I.rx_uart_i.fifo_i.cnt[0] ),
    .C(\soc_I.rx_uart_i.fifo_i.cnt[3] ),
    .Y(_13236_),
    .D(\soc_I.rx_uart_i.fifo_i.cnt[2] ));
 sg13g2_nor2b_2 _22240_ (.A(\soc_I.rx_uart_i.fifo_i.cnt[4] ),
    .B_N(_13236_),
    .Y(_13237_));
 sg13g2_nand2b_2 _22241_ (.Y(_13238_),
    .B(net9240),
    .A_N(_13237_));
 sg13g2_mux2_1 _22242_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[8][0] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[9][0] ),
    .S(net9191),
    .X(_13239_));
 sg13g2_nor2b_1 _22243_ (.A(\soc_I.rx_uart_i.fifo_i.ram[11][0] ),
    .B_N(net9191),
    .Y(_13240_));
 sg13g2_o21ai_1 _22244_ (.B1(net9181),
    .Y(_13241_),
    .A1(net9191),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[10][0] ));
 sg13g2_o21ai_1 _22245_ (.B1(net8981),
    .Y(_13242_),
    .A1(net9188),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[12][0] ));
 sg13g2_a21oi_1 _22246_ (.A1(net9188),
    .A2(_10675_),
    .Y(_13243_),
    .B1(_13242_));
 sg13g2_nor2b_1 _22247_ (.A(\soc_I.rx_uart_i.fifo_i.ram[15][0] ),
    .B_N(net9188),
    .Y(_13244_));
 sg13g2_o21ai_1 _22248_ (.B1(net9182),
    .Y(_13245_),
    .A1(net9188),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[14][0] ));
 sg13g2_mux4_1 _22249_ (.S0(net9194),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[4][0] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[5][0] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[6][0] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[7][0] ),
    .S1(net9180),
    .X(_13246_));
 sg13g2_nor2_1 _22250_ (.A(net9173),
    .B(_13246_),
    .Y(_13247_));
 sg13g2_o21ai_1 _22251_ (.B1(net9174),
    .Y(_13248_),
    .A1(_13244_),
    .A2(_13245_));
 sg13g2_o21ai_1 _22252_ (.B1(net9178),
    .Y(_13249_),
    .A1(_13243_),
    .A2(_13248_));
 sg13g2_nor2_1 _22253_ (.A(_13247_),
    .B(_13249_),
    .Y(_13250_));
 sg13g2_mux4_1 _22254_ (.S0(net9187),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[0][0] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[1][0] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[2][0] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[3][0] ),
    .S1(net9180),
    .X(_13251_));
 sg13g2_nor2_1 _22255_ (.A(net9175),
    .B(_13251_),
    .Y(_13252_));
 sg13g2_o21ai_1 _22256_ (.B1(net9174),
    .Y(_13253_),
    .A1(_13240_),
    .A2(_13241_));
 sg13g2_a21oi_1 _22257_ (.A1(net8981),
    .A2(_13239_),
    .Y(_13254_),
    .B1(_13253_));
 sg13g2_nor3_1 _22258_ (.A(net9177),
    .B(_13252_),
    .C(_13254_),
    .Y(_13255_));
 sg13g2_nor3_2 _22259_ (.A(net8675),
    .B(_13250_),
    .C(_13255_),
    .Y(_13256_));
 sg13g2_nand3b_1 _22260_ (.B(_12511_),
    .C(_13148_),
    .Y(_13257_),
    .A_N(_12500_));
 sg13g2_nor4_2 _22261_ (.A(_12500_),
    .B(_12510_),
    .C(_13147_),
    .Y(_13258_),
    .D(_13149_));
 sg13g2_nand2b_2 _22262_ (.Y(_13259_),
    .B(_13258_),
    .A_N(_13174_));
 sg13g2_nor2_2 _22263_ (.A(_13051_),
    .B(_13259_),
    .Y(_13260_));
 sg13g2_nor2_2 _22264_ (.A(net7468),
    .B(_13259_),
    .Y(_13261_));
 sg13g2_nor4_2 _22265_ (.A(net7493),
    .B(_13045_),
    .C(_13178_),
    .Y(_13262_),
    .D(_13259_));
 sg13g2_or3_1 _22266_ (.A(_13260_),
    .B(_13261_),
    .C(_13262_),
    .X(_13263_));
 sg13g2_nand3b_1 _22267_ (.B(net7480),
    .C(_13159_),
    .Y(_13264_),
    .A_N(_13257_));
 sg13g2_nand3_1 _22268_ (.B(_13123_),
    .C(_13258_),
    .A(_12879_),
    .Y(_13265_));
 sg13g2_a21oi_1 _22269_ (.A1(net7468),
    .A2(_13051_),
    .Y(_13266_),
    .B1(_13265_));
 sg13g2_or4_1 _22270_ (.A(_12489_),
    .B(_12510_),
    .C(_13047_),
    .D(_13160_),
    .X(_13267_));
 sg13g2_nor4_1 _22271_ (.A(net7493),
    .B(_13045_),
    .C(_13178_),
    .D(_13259_),
    .Y(_13268_));
 sg13g2_a21oi_1 _22272_ (.A1(net7468),
    .A2(_13052_),
    .Y(_13269_),
    .B1(_13259_));
 sg13g2_o21ai_1 _22273_ (.B1(_13173_),
    .Y(_13270_),
    .A1(_13268_),
    .A2(_13269_));
 sg13g2_a21o_1 _22274_ (.A2(_13211_),
    .A1(_13046_),
    .B1(_13226_),
    .X(_13271_));
 sg13g2_o21ai_1 _22275_ (.B1(net7480),
    .Y(_13272_),
    .A1(_13222_),
    .A2(_13271_));
 sg13g2_nor2_1 _22276_ (.A(_13161_),
    .B(_13257_),
    .Y(_13273_));
 sg13g2_or2_1 _22277_ (.X(_13274_),
    .B(_13257_),
    .A(_13161_));
 sg13g2_nand3_1 _22278_ (.B(_13165_),
    .C(_13273_),
    .A(_13049_),
    .Y(_13275_));
 sg13g2_nand4_1 _22279_ (.B(_13123_),
    .C(_13156_),
    .A(_10604_),
    .Y(_13276_),
    .D(_13258_));
 sg13g2_and2_1 _22280_ (.A(_13275_),
    .B(_13276_),
    .X(_13277_));
 sg13g2_nor3_1 _22281_ (.A(net9244),
    .B(net7468),
    .C(_13274_),
    .Y(_13278_));
 sg13g2_nor3_1 _22282_ (.A(\soc_I.div_ready ),
    .B(_13157_),
    .C(_13274_),
    .Y(_13279_));
 sg13g2_nor3_1 _22283_ (.A(net9250),
    .B(net7468),
    .C(_13274_),
    .Y(_13280_));
 sg13g2_nor4_1 _22284_ (.A(_13266_),
    .B(_13278_),
    .C(_13279_),
    .D(_13280_),
    .Y(_13281_));
 sg13g2_nand4_1 _22285_ (.B(_13272_),
    .C(_13277_),
    .A(_13270_),
    .Y(_13282_),
    .D(_13281_));
 sg13g2_a221oi_1 _22286_ (.B2(_12882_),
    .C1(_13149_),
    .B1(_13282_),
    .A1(_12500_),
    .Y(_13283_),
    .A2(_13267_));
 sg13g2_nor2_1 _22287_ (.A(net9267),
    .B(\soc_I.uart_lsr_rdy ),
    .Y(_13284_));
 sg13g2_nand2_2 _22288_ (.Y(_13285_),
    .A(_13283_),
    .B(_13284_));
 sg13g2_nor3_1 _22289_ (.A(_13234_),
    .B(_13256_),
    .C(_13285_),
    .Y(_13286_));
 sg13g2_a21o_2 _22290_ (.A2(\soc_I.qqspi_I.rdata[0] ),
    .A1(net9269),
    .B1(_13286_),
    .X(_13287_));
 sg13g2_o21ai_1 _22291_ (.B1(_10952_),
    .Y(_13288_),
    .A1(_00188_),
    .A2(_10925_));
 sg13g2_nor2_2 _22292_ (.A(net9708),
    .B(_10587_),
    .Y(_13289_));
 sg13g2_nand2_2 _22293_ (.Y(_13290_),
    .A(net9702),
    .B(_13289_));
 sg13g2_nand4_1 _22294_ (.B(\soc_I.kianv_I.Instr[2] ),
    .C(\soc_I.kianv_I.Instr[1] ),
    .A(\soc_I.kianv_I.Instr[3] ),
    .Y(_13291_),
    .D(\soc_I.kianv_I.Instr[0] ));
 sg13g2_nor3_1 _22295_ (.A(_11054_),
    .B(_13290_),
    .C(_13291_),
    .Y(_13292_));
 sg13g2_or4_1 _22296_ (.A(net9712),
    .B(_11005_),
    .C(_13290_),
    .D(_13291_),
    .X(_13293_));
 sg13g2_o21ai_1 _22297_ (.B1(_13288_),
    .Y(_13294_),
    .A1(_10903_),
    .A2(_13293_));
 sg13g2_nand2_1 _22298_ (.Y(_13295_),
    .A(_10916_),
    .B(_11001_));
 sg13g2_and2_1 _22299_ (.A(_13294_),
    .B(_13295_),
    .X(_13296_));
 sg13g2_nand2_1 _22300_ (.Y(_13297_),
    .A(_13294_),
    .B(_13295_));
 sg13g2_a21o_2 _22301_ (.A2(_10919_),
    .A1(_00188_),
    .B1(_13294_),
    .X(_13298_));
 sg13g2_nor2b_1 _22302_ (.A(net9707),
    .B_N(_13298_),
    .Y(_13299_));
 sg13g2_nor2_1 _22303_ (.A(net9421),
    .B(net8373),
    .Y(_13300_));
 sg13g2_nor2_1 _22304_ (.A(net8497),
    .B(_13300_),
    .Y(_13301_));
 sg13g2_o21ai_1 _22305_ (.B1(net8494),
    .Y(_13302_),
    .A1(net9422),
    .A2(net8373));
 sg13g2_nor2_2 _22306_ (.A(\soc_I.kianv_I.datapath_unit_I.ADDR_I.q[0] ),
    .B(net9421),
    .Y(_13303_));
 sg13g2_nor2_2 _22307_ (.A(_13302_),
    .B(_13303_),
    .Y(_13304_));
 sg13g2_or2_1 _22308_ (.X(_13305_),
    .B(_13303_),
    .A(_13302_));
 sg13g2_nand2_1 _22309_ (.Y(_13306_),
    .A(_13287_),
    .B(_13305_));
 sg13g2_nand2b_1 _22310_ (.Y(_13307_),
    .B(net7450),
    .A_N(_00075_));
 sg13g2_nor2_1 _22311_ (.A(_00077_),
    .B(net7437),
    .Y(_13308_));
 sg13g2_a221oi_1 _22312_ (.B2(\soc_I.clint_I.mtime[40] ),
    .C1(_13308_),
    .B1(net7440),
    .A1(_10673_),
    .Y(_13309_),
    .A2(net7445));
 sg13g2_nand3_1 _22313_ (.B(_13307_),
    .C(_13309_),
    .A(net9290),
    .Y(_13310_));
 sg13g2_a22oi_1 _22314_ (.Y(_13311_),
    .B1(net8832),
    .B2(\soc_I.spi0_I.div[8] ),
    .A2(_10672_),
    .A1(net9254));
 sg13g2_a21oi_1 _22315_ (.A1(net8989),
    .A2(_13311_),
    .Y(_13312_),
    .B1(net9247));
 sg13g2_a21o_2 _22316_ (.A2(_13312_),
    .A1(_13310_),
    .B1(net9240),
    .X(_13313_));
 sg13g2_a21o_1 _22317_ (.A2(_13313_),
    .A1(net8676),
    .B1(\soc_I.uart_lsr_rdy ),
    .X(_13314_));
 sg13g2_a21oi_1 _22318_ (.A1(\soc_I.uart_lsr_rdy ),
    .A2(_13237_),
    .Y(_13315_),
    .B1(_13201_));
 sg13g2_nand2b_1 _22319_ (.Y(_13316_),
    .B(_13283_),
    .A_N(net9267));
 sg13g2_a22oi_1 _22320_ (.Y(_13317_),
    .B1(_13314_),
    .B2(_13315_),
    .A2(\soc_I.qqspi_I.rdata[8] ),
    .A1(net9266));
 sg13g2_and2_2 _22321_ (.A(\soc_I.kianv_I.datapath_unit_I.ADDR_I.q[0] ),
    .B(_13299_),
    .X(_13318_));
 sg13g2_nand2_1 _22322_ (.Y(_13319_),
    .A(\soc_I.kianv_I.datapath_unit_I.ADDR_I.q[0] ),
    .B(net8373));
 sg13g2_nor3_1 _22323_ (.A(net9421),
    .B(_13317_),
    .C(_13319_),
    .Y(_13320_));
 sg13g2_o21ai_1 _22324_ (.B1(net9292),
    .Y(_13321_),
    .A1(_00016_),
    .A2(net7425));
 sg13g2_inv_1 _22325_ (.Y(_13322_),
    .A(_13321_));
 sg13g2_nor2_1 _22326_ (.A(_00018_),
    .B(net7438),
    .Y(_13323_));
 sg13g2_a221oi_1 _22327_ (.B2(\soc_I.clint_I.mtime[56] ),
    .C1(_13323_),
    .B1(net7442),
    .A1(_10655_),
    .Y(_13324_),
    .A2(net7447));
 sg13g2_a22oi_1 _22328_ (.Y(_13325_),
    .B1(net8833),
    .B2(\soc_I.spi_div_reg[24] ),
    .A2(\soc_I.div_ready ),
    .A1(_10598_));
 sg13g2_a221oi_1 _22329_ (.B2(net8992),
    .C1(net9249),
    .B1(_13325_),
    .A1(_13322_),
    .Y(_13326_),
    .A2(_13324_));
 sg13g2_or2_1 _22330_ (.X(_13327_),
    .B(_13326_),
    .A(net9244));
 sg13g2_nor2b_1 _22331_ (.A(_13285_),
    .B_N(net8676),
    .Y(_13328_));
 sg13g2_nand3_1 _22332_ (.B(_13283_),
    .C(_13284_),
    .A(net8676),
    .Y(_13329_));
 sg13g2_a22oi_1 _22333_ (.Y(_13330_),
    .B1(_13327_),
    .B2(net7361),
    .A2(\soc_I.qqspi_I.rdata[24] ),
    .A1(net9267));
 sg13g2_nand2_1 _22334_ (.Y(_13331_),
    .A(net9422),
    .B(_13318_));
 sg13g2_o21ai_1 _22335_ (.B1(net9291),
    .Y(_13332_),
    .A1(_00013_),
    .A2(net7424));
 sg13g2_nor2_1 _22336_ (.A(_00015_),
    .B(net7437),
    .Y(_13333_));
 sg13g2_a221oi_1 _22337_ (.B2(\soc_I.clint_I.mtime[48] ),
    .C1(_13333_),
    .B1(net7441),
    .A1(_10654_),
    .Y(_13334_),
    .A2(net7446));
 sg13g2_nand2b_1 _22338_ (.Y(_13335_),
    .B(_13334_),
    .A_N(_13332_));
 sg13g2_o21ai_1 _22339_ (.B1(net8992),
    .Y(_13336_),
    .A1(net8999),
    .A2(_00012_));
 sg13g2_a21oi_1 _22340_ (.A1(\soc_I.spi_div_reg[16] ),
    .A2(net8833),
    .Y(_13337_),
    .B1(_13336_));
 sg13g2_nor2_1 _22341_ (.A(net9249),
    .B(_13337_),
    .Y(_13338_));
 sg13g2_a21o_1 _22342_ (.A2(_13338_),
    .A1(_13335_),
    .B1(net9244),
    .X(_13339_));
 sg13g2_a22oi_1 _22343_ (.Y(_13340_),
    .B1(net7362),
    .B2(_13339_),
    .A2(\soc_I.qqspi_I.rdata[16] ),
    .A1(net9269));
 sg13g2_nand2b_2 _22344_ (.Y(_13341_),
    .B(net9422),
    .A_N(_13299_));
 sg13g2_nor2_2 _22345_ (.A(_10647_),
    .B(_13318_),
    .Y(_13342_));
 sg13g2_nand2b_1 _22346_ (.Y(_13343_),
    .B(_13342_),
    .A_N(_13340_));
 sg13g2_o21ai_1 _22347_ (.B1(_13343_),
    .Y(_13344_),
    .A1(_13330_),
    .A2(_13331_));
 sg13g2_o21ai_1 _22348_ (.B1(net8493),
    .Y(_13345_),
    .A1(_13320_),
    .A2(_13344_));
 sg13g2_nand2_1 _22349_ (.Y(\soc_I.kianv_I.datapath_unit_I.Data[0] ),
    .A(_13306_),
    .B(_13345_));
 sg13g2_nand2_1 _22350_ (.Y(_13346_),
    .A(net9266),
    .B(\soc_I.qqspi_I.rdata[1] ));
 sg13g2_nand2b_1 _22351_ (.Y(_13347_),
    .B(net9190),
    .A_N(\soc_I.rx_uart_i.fifo_i.ram[9][1] ));
 sg13g2_o21ai_1 _22352_ (.B1(_13347_),
    .Y(_13348_),
    .A1(net9190),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[8][1] ));
 sg13g2_mux2_1 _22353_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[10][1] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[11][1] ),
    .S(net9191),
    .X(_13349_));
 sg13g2_o21ai_1 _22354_ (.B1(net8981),
    .Y(_13350_),
    .A1(net9186),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[12][1] ));
 sg13g2_a21oi_1 _22355_ (.A1(net9186),
    .A2(_10677_),
    .Y(_13351_),
    .B1(_13350_));
 sg13g2_nor2b_1 _22356_ (.A(\soc_I.rx_uart_i.fifo_i.ram[15][1] ),
    .B_N(net9185),
    .Y(_13352_));
 sg13g2_o21ai_1 _22357_ (.B1(net9179),
    .Y(_13353_),
    .A1(net9184),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[14][1] ));
 sg13g2_mux4_1 _22358_ (.S0(net9184),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[4][1] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[5][1] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[6][1] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[7][1] ),
    .S1(net9179),
    .X(_13354_));
 sg13g2_nor2_1 _22359_ (.A(net9172),
    .B(_13354_),
    .Y(_13355_));
 sg13g2_o21ai_1 _22360_ (.B1(net9172),
    .Y(_13356_),
    .A1(_13352_),
    .A2(_13353_));
 sg13g2_o21ai_1 _22361_ (.B1(net9178),
    .Y(_13357_),
    .A1(_13351_),
    .A2(_13356_));
 sg13g2_nor2_2 _22362_ (.A(_13355_),
    .B(_13357_),
    .Y(_13358_));
 sg13g2_mux4_1 _22363_ (.S0(net9193),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[0][1] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[1][1] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[2][1] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[3][1] ),
    .S1(net9183),
    .X(_13359_));
 sg13g2_a21oi_1 _22364_ (.A1(net9182),
    .A2(_13349_),
    .Y(_13360_),
    .B1(_10676_));
 sg13g2_o21ai_1 _22365_ (.B1(_13360_),
    .Y(_13361_),
    .A1(net9181),
    .A2(_13348_));
 sg13g2_o21ai_1 _22366_ (.B1(_13361_),
    .Y(_13362_),
    .A1(net9175),
    .A2(_13359_));
 sg13g2_nor2_1 _22367_ (.A(net8675),
    .B(_13358_),
    .Y(_13363_));
 sg13g2_o21ai_1 _22368_ (.B1(_13363_),
    .Y(_13364_),
    .A1(net9177),
    .A2(_13362_));
 sg13g2_o21ai_1 _22369_ (.B1(net9291),
    .Y(_13365_),
    .A1(_00115_),
    .A2(net7424));
 sg13g2_nor3_1 _22370_ (.A(_00116_),
    .B(net7467),
    .C(net7465),
    .Y(_13366_));
 sg13g2_nand2_1 _22371_ (.Y(_13367_),
    .A(\soc_I.clint_I.mtime[33] ),
    .B(net7444));
 sg13g2_o21ai_1 _22372_ (.B1(_13367_),
    .Y(_13368_),
    .A1(_00117_),
    .A2(net7439));
 sg13g2_nor3_1 _22373_ (.A(_13365_),
    .B(_13366_),
    .C(_13368_),
    .Y(_13369_));
 sg13g2_nand3_1 _22374_ (.B(net8960),
    .C(net7491),
    .A(\soc_I.spi0_I.rx_data[1] ),
    .Y(_13370_));
 sg13g2_a21oi_1 _22375_ (.A1(\soc_I.gpio0_I.rdata[1] ),
    .A2(_13205_),
    .Y(_13371_),
    .B1(net9253));
 sg13g2_a22oi_1 _22376_ (.Y(_13372_),
    .B1(_13370_),
    .B2(_13371_),
    .A2(_00114_),
    .A1(net9253));
 sg13g2_o21ai_1 _22377_ (.B1(net8991),
    .Y(_13373_),
    .A1(net8996),
    .A2(_00113_));
 sg13g2_a21oi_1 _22378_ (.A1(net8998),
    .A2(_13372_),
    .Y(_13374_),
    .B1(_13373_));
 sg13g2_nor3_1 _22379_ (.A(net9248),
    .B(_13369_),
    .C(_13374_),
    .Y(_13375_));
 sg13g2_o21ai_1 _22380_ (.B1(_13364_),
    .Y(_13376_),
    .A1(net9242),
    .A2(_13375_));
 sg13g2_o21ai_1 _22381_ (.B1(_13346_),
    .Y(_13377_),
    .A1(_13285_),
    .A2(_13376_));
 sg13g2_o21ai_1 _22382_ (.B1(net9292),
    .Y(_13378_),
    .A1(_00024_),
    .A2(net7425));
 sg13g2_nor2_1 _22383_ (.A(_00026_),
    .B(net7438),
    .Y(_13379_));
 sg13g2_a221oi_1 _22384_ (.B2(\soc_I.clint_I.mtime[57] ),
    .C1(_13379_),
    .B1(net7442),
    .A1(_10658_),
    .Y(_13380_),
    .A2(net7447));
 sg13g2_nand2b_1 _22385_ (.Y(_13381_),
    .B(_13380_),
    .A_N(_13378_));
 sg13g2_o21ai_1 _22386_ (.B1(net8993),
    .Y(_13382_),
    .A1(net9000),
    .A2(_00023_));
 sg13g2_a21oi_1 _22387_ (.A1(\soc_I.spi_div_reg[25] ),
    .A2(net8834),
    .Y(_13383_),
    .B1(_13382_));
 sg13g2_nor2_1 _22388_ (.A(net9250),
    .B(_13383_),
    .Y(_13384_));
 sg13g2_a21oi_1 _22389_ (.A1(_13381_),
    .A2(_13384_),
    .Y(_13385_),
    .B1(net9245));
 sg13g2_inv_1 _22390_ (.Y(_13386_),
    .A(_13385_));
 sg13g2_a22oi_1 _22391_ (.Y(_13387_),
    .B1(net7361),
    .B2(_13386_),
    .A2(\soc_I.qqspi_I.rdata[25] ),
    .A1(net9268));
 sg13g2_and2_1 _22392_ (.A(net9421),
    .B(_13387_),
    .X(_13388_));
 sg13g2_nand2b_1 _22393_ (.Y(_13389_),
    .B(net7445),
    .A_N(_00080_));
 sg13g2_nand2b_1 _22394_ (.Y(_13390_),
    .B(net7450),
    .A_N(_00079_));
 sg13g2_a22oi_1 _22395_ (.Y(_13391_),
    .B1(_13229_),
    .B2(_10682_),
    .A2(net7440),
    .A1(\soc_I.clint_I.mtime[41] ));
 sg13g2_nand4_1 _22396_ (.B(_13389_),
    .C(_13390_),
    .A(net9290),
    .Y(_13392_),
    .D(_13391_));
 sg13g2_o21ai_1 _22397_ (.B1(net8988),
    .Y(_13393_),
    .A1(net8997),
    .A2(_00078_));
 sg13g2_a21oi_1 _22398_ (.A1(\soc_I.spi0_I.div[9] ),
    .A2(net8832),
    .Y(_13394_),
    .B1(_13393_));
 sg13g2_nor2_1 _22399_ (.A(net9247),
    .B(_13394_),
    .Y(_13395_));
 sg13g2_a21o_2 _22400_ (.A2(_13395_),
    .A1(_13392_),
    .B1(net9240),
    .X(_13396_));
 sg13g2_a22oi_1 _22401_ (.Y(_13397_),
    .B1(net7362),
    .B2(_13396_),
    .A2(\soc_I.qqspi_I.rdata[9] ),
    .A1(net9270));
 sg13g2_a21oi_1 _22402_ (.A1(_10647_),
    .A2(_13397_),
    .Y(_13398_),
    .B1(_13388_));
 sg13g2_nand2_1 _22403_ (.Y(_13399_),
    .A(_13318_),
    .B(_13398_));
 sg13g2_nand2_1 _22404_ (.Y(_13400_),
    .A(net9269),
    .B(\soc_I.qqspi_I.rdata[17] ));
 sg13g2_nand2b_1 _22405_ (.Y(_13401_),
    .B(net7451),
    .A_N(_00020_));
 sg13g2_nor2_1 _22406_ (.A(_00022_),
    .B(net7437),
    .Y(_13402_));
 sg13g2_a221oi_1 _22407_ (.B2(\soc_I.clint_I.mtime[49] ),
    .C1(_13402_),
    .B1(net7441),
    .A1(_10657_),
    .Y(_13403_),
    .A2(net7446));
 sg13g2_nand3_1 _22408_ (.B(_13401_),
    .C(_13403_),
    .A(net9291),
    .Y(_13404_));
 sg13g2_o21ai_1 _22409_ (.B1(net8992),
    .Y(_13405_),
    .A1(net8999),
    .A2(_00019_));
 sg13g2_a21oi_1 _22410_ (.A1(\soc_I.spi_div_reg[17] ),
    .A2(net8833),
    .Y(_13406_),
    .B1(_13405_));
 sg13g2_nor2_1 _22411_ (.A(net9249),
    .B(_13406_),
    .Y(_13407_));
 sg13g2_a21oi_1 _22412_ (.A1(_13404_),
    .A2(_13407_),
    .Y(_13408_),
    .B1(net9244));
 sg13g2_o21ai_1 _22413_ (.B1(_13400_),
    .Y(_13409_),
    .A1(_13329_),
    .A2(_13408_));
 sg13g2_inv_1 _22414_ (.Y(_13410_),
    .A(_13409_));
 sg13g2_nand2_1 _22415_ (.Y(_13411_),
    .A(_13342_),
    .B(_13409_));
 sg13g2_a21oi_1 _22416_ (.A1(_13399_),
    .A2(_13411_),
    .Y(_13412_),
    .B1(net8498));
 sg13g2_a21o_2 _22417_ (.A2(_13377_),
    .A1(_13305_),
    .B1(_13412_),
    .X(\soc_I.kianv_I.datapath_unit_I.Data[1] ));
 sg13g2_mux2_1 _22418_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[8][2] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[9][2] ),
    .S(net9190),
    .X(_13413_));
 sg13g2_nand2_1 _22419_ (.Y(_13414_),
    .A(net8982),
    .B(_13413_));
 sg13g2_mux2_1 _22420_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[10][2] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[11][2] ),
    .S(net9190),
    .X(_13415_));
 sg13g2_mux2_1 _22421_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[12][2] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[13][2] ),
    .S(net9188),
    .X(_13416_));
 sg13g2_nand2_1 _22422_ (.Y(_13417_),
    .A(net8982),
    .B(_13416_));
 sg13g2_mux2_1 _22423_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[14][2] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[15][2] ),
    .S(net9186),
    .X(_13418_));
 sg13g2_mux4_1 _22424_ (.S0(net9193),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[0][2] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[1][2] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[2][2] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[3][2] ),
    .S1(net9183),
    .X(_13419_));
 sg13g2_a21oi_1 _22425_ (.A1(net9181),
    .A2(_13415_),
    .Y(_13420_),
    .B1(_10676_));
 sg13g2_a21oi_1 _22426_ (.A1(_13414_),
    .A2(_13420_),
    .Y(_13421_),
    .B1(net9177));
 sg13g2_o21ai_1 _22427_ (.B1(_13421_),
    .Y(_13422_),
    .A1(net9174),
    .A2(_13419_));
 sg13g2_a21oi_1 _22428_ (.A1(net9182),
    .A2(_13418_),
    .Y(_13423_),
    .B1(_10676_));
 sg13g2_mux4_1 _22429_ (.S0(net9185),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[4][2] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[5][2] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[6][2] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[7][2] ),
    .S1(net9179),
    .X(_13424_));
 sg13g2_o21ai_1 _22430_ (.B1(net9178),
    .Y(_13425_),
    .A1(net9172),
    .A2(_13424_));
 sg13g2_a21oi_2 _22431_ (.B1(_13425_),
    .Y(_13426_),
    .A2(_13423_),
    .A1(_13417_));
 sg13g2_nor2_1 _22432_ (.A(net8675),
    .B(_13426_),
    .Y(_13427_));
 sg13g2_a21oi_1 _22433_ (.A1(_10686_),
    .A2(net7451),
    .Y(_13428_),
    .B1(net8991));
 sg13g2_o21ai_1 _22434_ (.B1(_13428_),
    .Y(_13429_),
    .A1(_00122_),
    .A2(_13223_));
 sg13g2_a221oi_1 _22435_ (.B2(\soc_I.clint_I.mtime[34] ),
    .C1(_13429_),
    .B1(_13224_),
    .A1(_10685_),
    .Y(_13430_),
    .A2(net7446));
 sg13g2_nand3_1 _22436_ (.B(net8960),
    .C(net7491),
    .A(\soc_I.spi0_I.rx_data[2] ),
    .Y(_13431_));
 sg13g2_a21oi_1 _22437_ (.A1(\soc_I.gpio0_I.rdata[2] ),
    .A2(_13205_),
    .Y(_13432_),
    .B1(net9253));
 sg13g2_a22oi_1 _22438_ (.Y(_13433_),
    .B1(_13431_),
    .B2(_13432_),
    .A2(_00119_),
    .A1(net9252));
 sg13g2_o21ai_1 _22439_ (.B1(net8989),
    .Y(_13434_),
    .A1(net8996),
    .A2(_00118_));
 sg13g2_a21oi_1 _22440_ (.A1(net8995),
    .A2(_13433_),
    .Y(_13435_),
    .B1(_13434_));
 sg13g2_nor3_1 _22441_ (.A(net9246),
    .B(_13430_),
    .C(_13435_),
    .Y(_13436_));
 sg13g2_nor2_1 _22442_ (.A(net9240),
    .B(_13436_),
    .Y(_13437_));
 sg13g2_a21oi_2 _22443_ (.B1(_13437_),
    .Y(_13438_),
    .A2(_13427_),
    .A1(_13422_));
 sg13g2_a22oi_1 _22444_ (.Y(_13439_),
    .B1(_13202_),
    .B2(_13438_),
    .A2(\soc_I.qqspi_I.rdata[2] ),
    .A1(net9266));
 sg13g2_nand2_1 _22445_ (.Y(_13440_),
    .A(net9267),
    .B(\soc_I.qqspi_I.rdata[26] ));
 sg13g2_o21ai_1 _22446_ (.B1(net9293),
    .Y(_13441_),
    .A1(_00032_),
    .A2(net7425));
 sg13g2_nor3_1 _22447_ (.A(_00033_),
    .B(_13050_),
    .C(net7466),
    .Y(_13442_));
 sg13g2_nand2_1 _22448_ (.Y(_13443_),
    .A(\soc_I.clint_I.mtime[58] ),
    .B(net7442));
 sg13g2_o21ai_1 _22449_ (.B1(_13443_),
    .Y(_13444_),
    .A1(_00034_),
    .A2(net7438));
 sg13g2_nor3_1 _22450_ (.A(_13441_),
    .B(_13442_),
    .C(_13444_),
    .Y(_13445_));
 sg13g2_o21ai_1 _22451_ (.B1(net8993),
    .Y(_13446_),
    .A1(net8999),
    .A2(_00031_));
 sg13g2_a21oi_2 _22452_ (.B1(_13446_),
    .Y(_13447_),
    .A2(net8834),
    .A1(\soc_I.spi_div_reg[26] ));
 sg13g2_nor3_1 _22453_ (.A(net9249),
    .B(_13445_),
    .C(_13447_),
    .Y(_13448_));
 sg13g2_nor2_1 _22454_ (.A(net9243),
    .B(_13448_),
    .Y(_13449_));
 sg13g2_o21ai_1 _22455_ (.B1(_13440_),
    .Y(_13450_),
    .A1(_13329_),
    .A2(_13449_));
 sg13g2_inv_2 _22456_ (.Y(_13451_),
    .A(_13450_));
 sg13g2_nor2_1 _22457_ (.A(_10647_),
    .B(_13450_),
    .Y(_13452_));
 sg13g2_nand2b_1 _22458_ (.Y(_13453_),
    .B(net7445),
    .A_N(_00084_));
 sg13g2_nand2b_1 _22459_ (.Y(_13454_),
    .B(net7450),
    .A_N(_00083_));
 sg13g2_a22oi_1 _22460_ (.Y(_13455_),
    .B1(_13229_),
    .B2(_10683_),
    .A2(net7440),
    .A1(\soc_I.clint_I.mtime[42] ));
 sg13g2_nand4_1 _22461_ (.B(_13453_),
    .C(_13454_),
    .A(net9290),
    .Y(_13456_),
    .D(_13455_));
 sg13g2_o21ai_1 _22462_ (.B1(net8988),
    .Y(_13457_),
    .A1(net8996),
    .A2(_00082_));
 sg13g2_a21oi_1 _22463_ (.A1(\soc_I.spi0_I.div[10] ),
    .A2(net8832),
    .Y(_13458_),
    .B1(_13457_));
 sg13g2_nor2_1 _22464_ (.A(net9247),
    .B(_13458_),
    .Y(_13459_));
 sg13g2_a21o_2 _22465_ (.A2(_13459_),
    .A1(_13456_),
    .B1(net9240),
    .X(_13460_));
 sg13g2_a22oi_1 _22466_ (.Y(_13461_),
    .B1(net7362),
    .B2(_13460_),
    .A2(\soc_I.qqspi_I.rdata[10] ),
    .A1(net9270));
 sg13g2_a21oi_1 _22467_ (.A1(_10647_),
    .A2(_13461_),
    .Y(_13462_),
    .B1(_13452_));
 sg13g2_nand2_1 _22468_ (.Y(_13463_),
    .A(net9270),
    .B(\soc_I.qqspi_I.rdata[18] ));
 sg13g2_nand2b_1 _22469_ (.Y(_13464_),
    .B(net7451),
    .A_N(_00028_));
 sg13g2_nand2b_1 _22470_ (.Y(_13465_),
    .B(net7446),
    .A_N(_00029_));
 sg13g2_a22oi_1 _22471_ (.Y(_13466_),
    .B1(_13229_),
    .B2(_10659_),
    .A2(net7441),
    .A1(\soc_I.clint_I.mtime[50] ));
 sg13g2_nand4_1 _22472_ (.B(_13464_),
    .C(_13465_),
    .A(net9291),
    .Y(_13467_),
    .D(_13466_));
 sg13g2_o21ai_1 _22473_ (.B1(net8994),
    .Y(_13468_),
    .A1(net8998),
    .A2(_00027_));
 sg13g2_a21oi_1 _22474_ (.A1(\soc_I.spi_div_reg[18] ),
    .A2(net8832),
    .Y(_13469_),
    .B1(_13468_));
 sg13g2_nor2_2 _22475_ (.A(net9248),
    .B(_13469_),
    .Y(_13470_));
 sg13g2_a21oi_2 _22476_ (.B1(net9242),
    .Y(_13471_),
    .A2(_13470_),
    .A1(_13467_));
 sg13g2_o21ai_1 _22477_ (.B1(_13463_),
    .Y(_13472_),
    .A1(_13329_),
    .A2(_13471_));
 sg13g2_inv_1 _22478_ (.Y(_13473_),
    .A(_13472_));
 sg13g2_a22oi_1 _22479_ (.Y(_13474_),
    .B1(_13472_),
    .B2(_13342_),
    .A2(_13462_),
    .A1(_13318_));
 sg13g2_or2_1 _22480_ (.X(_13475_),
    .B(_13474_),
    .A(net8498));
 sg13g2_o21ai_1 _22481_ (.B1(_13475_),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[2] ),
    .A1(_13304_),
    .A2(_13439_));
 sg13g2_a22oi_1 _22482_ (.Y(_13476_),
    .B1(_13224_),
    .B2(\soc_I.clint_I.mtime[35] ),
    .A2(net7449),
    .A1(_10687_));
 sg13g2_nand2b_1 _22483_ (.Y(_13477_),
    .B(net7451),
    .A_N(_00125_));
 sg13g2_or2_1 _22484_ (.X(_13478_),
    .B(_13223_),
    .A(_00127_));
 sg13g2_nand4_1 _22485_ (.B(_13476_),
    .C(_13477_),
    .A(net9290),
    .Y(_13479_),
    .D(_13478_));
 sg13g2_nand3_1 _22486_ (.B(net8960),
    .C(net7491),
    .A(\soc_I.spi0_I.rx_data[3] ),
    .Y(_13480_));
 sg13g2_a21oi_1 _22487_ (.A1(\soc_I.gpio0_I.rdata[3] ),
    .A2(_13205_),
    .Y(_13481_),
    .B1(net9252));
 sg13g2_a22oi_1 _22488_ (.Y(_13482_),
    .B1(_13480_),
    .B2(_13481_),
    .A2(_00124_),
    .A1(net9252));
 sg13g2_o21ai_1 _22489_ (.B1(net8989),
    .Y(_13483_),
    .A1(net8995),
    .A2(_00123_));
 sg13g2_a21oi_1 _22490_ (.A1(net8995),
    .A2(_13482_),
    .Y(_13484_),
    .B1(_13483_));
 sg13g2_nor2_1 _22491_ (.A(net9247),
    .B(_13484_),
    .Y(_13485_));
 sg13g2_a21oi_1 _22492_ (.A1(_13479_),
    .A2(_13485_),
    .Y(_13486_),
    .B1(net9241));
 sg13g2_mux2_1 _22493_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[8][3] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[9][3] ),
    .S(net9189),
    .X(_13487_));
 sg13g2_nor2b_1 _22494_ (.A(\soc_I.rx_uart_i.fifo_i.ram[11][3] ),
    .B_N(net9189),
    .Y(_13488_));
 sg13g2_o21ai_1 _22495_ (.B1(net9182),
    .Y(_13489_),
    .A1(net9189),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[10][3] ));
 sg13g2_o21ai_1 _22496_ (.B1(net8981),
    .Y(_13490_),
    .A1(net9184),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[12][3] ));
 sg13g2_a21oi_1 _22497_ (.A1(net9184),
    .A2(_10678_),
    .Y(_13491_),
    .B1(_13490_));
 sg13g2_nor2b_1 _22498_ (.A(\soc_I.rx_uart_i.fifo_i.ram[15][3] ),
    .B_N(net9184),
    .Y(_13492_));
 sg13g2_o21ai_1 _22499_ (.B1(net9179),
    .Y(_13493_),
    .A1(net9184),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[14][3] ));
 sg13g2_mux4_1 _22500_ (.S0(net9187),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[0][3] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[1][3] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[2][3] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[3][3] ),
    .S1(net9180),
    .X(_13494_));
 sg13g2_nor2_1 _22501_ (.A(net9173),
    .B(_13494_),
    .Y(_13495_));
 sg13g2_o21ai_1 _22502_ (.B1(net9172),
    .Y(_13496_),
    .A1(_13488_),
    .A2(_13489_));
 sg13g2_a21oi_2 _22503_ (.B1(_13496_),
    .Y(_13497_),
    .A2(_13487_),
    .A1(net8981));
 sg13g2_nor3_1 _22504_ (.A(net9178),
    .B(_13495_),
    .C(_13497_),
    .Y(_13498_));
 sg13g2_mux4_1 _22505_ (.S0(net9187),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[4][3] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[5][3] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[6][3] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[7][3] ),
    .S1(net9180),
    .X(_13499_));
 sg13g2_nor2_1 _22506_ (.A(net9173),
    .B(_13499_),
    .Y(_13500_));
 sg13g2_o21ai_1 _22507_ (.B1(net9172),
    .Y(_13501_),
    .A1(_13492_),
    .A2(_13493_));
 sg13g2_o21ai_1 _22508_ (.B1(net9178),
    .Y(_13502_),
    .A1(_13491_),
    .A2(_13501_));
 sg13g2_nor2_1 _22509_ (.A(_13500_),
    .B(_13502_),
    .Y(_13503_));
 sg13g2_nor3_2 _22510_ (.A(net8675),
    .B(_13498_),
    .C(_13503_),
    .Y(_13504_));
 sg13g2_nor2_2 _22511_ (.A(_13486_),
    .B(_13504_),
    .Y(_13505_));
 sg13g2_a22oi_1 _22512_ (.Y(_13506_),
    .B1(_13202_),
    .B2(_13505_),
    .A2(\soc_I.qqspi_I.rdata[3] ),
    .A1(net9266));
 sg13g2_nand2b_1 _22513_ (.Y(_13507_),
    .B(net7452),
    .A_N(_00040_));
 sg13g2_nor2_1 _22514_ (.A(_00042_),
    .B(net7438),
    .Y(_13508_));
 sg13g2_a221oi_1 _22515_ (.B2(\soc_I.clint_I.mtime[59] ),
    .C1(_13508_),
    .B1(net7443),
    .A1(_10661_),
    .Y(_13509_),
    .A2(net7448));
 sg13g2_nand3_1 _22516_ (.B(_13507_),
    .C(_13509_),
    .A(net9292),
    .Y(_13510_));
 sg13g2_o21ai_1 _22517_ (.B1(net8993),
    .Y(_13511_),
    .A1(net9000),
    .A2(_00039_));
 sg13g2_a21oi_1 _22518_ (.A1(\soc_I.spi_div_reg[27] ),
    .A2(net8834),
    .Y(_13512_),
    .B1(_13511_));
 sg13g2_nor2_1 _22519_ (.A(net9249),
    .B(_13512_),
    .Y(_13513_));
 sg13g2_a21oi_1 _22520_ (.A1(_13510_),
    .A2(_13513_),
    .Y(_13514_),
    .B1(net9245));
 sg13g2_inv_1 _22521_ (.Y(_13515_),
    .A(_13514_));
 sg13g2_a22oi_1 _22522_ (.Y(_13516_),
    .B1(net7361),
    .B2(_13515_),
    .A2(\soc_I.qqspi_I.rdata[27] ),
    .A1(net9268));
 sg13g2_and2_1 _22523_ (.A(net9421),
    .B(_13516_),
    .X(_13517_));
 sg13g2_o21ai_1 _22524_ (.B1(net9290),
    .Y(_13518_),
    .A1(_00087_),
    .A2(net7424));
 sg13g2_nor3_1 _22525_ (.A(_00088_),
    .B(net7467),
    .C(net7465),
    .Y(_13519_));
 sg13g2_nand2_1 _22526_ (.Y(_13520_),
    .A(\soc_I.clint_I.mtime[43] ),
    .B(net7440));
 sg13g2_o21ai_1 _22527_ (.B1(_13520_),
    .Y(_13521_),
    .A1(_00089_),
    .A2(net7439));
 sg13g2_nor3_1 _22528_ (.A(_13518_),
    .B(_13519_),
    .C(_13521_),
    .Y(_13522_));
 sg13g2_o21ai_1 _22529_ (.B1(net8988),
    .Y(_13523_),
    .A1(net8997),
    .A2(_00086_));
 sg13g2_a21oi_2 _22530_ (.B1(_13523_),
    .Y(_13524_),
    .A2(net8832),
    .A1(\soc_I.spi0_I.div[11] ));
 sg13g2_nor3_1 _22531_ (.A(net9246),
    .B(_13522_),
    .C(_13524_),
    .Y(_13525_));
 sg13g2_or2_2 _22532_ (.X(_13526_),
    .B(_13525_),
    .A(net9240));
 sg13g2_a22oi_1 _22533_ (.Y(_13527_),
    .B1(net7362),
    .B2(_13526_),
    .A2(\soc_I.qqspi_I.rdata[11] ),
    .A1(net9270));
 sg13g2_a21oi_1 _22534_ (.A1(_10647_),
    .A2(_13527_),
    .Y(_13528_),
    .B1(_13517_));
 sg13g2_nand2_1 _22535_ (.Y(_13529_),
    .A(net9270),
    .B(\soc_I.qqspi_I.rdata[19] ));
 sg13g2_o21ai_1 _22536_ (.B1(net9290),
    .Y(_13530_),
    .A1(_00036_),
    .A2(net7424));
 sg13g2_nor2_1 _22537_ (.A(_00038_),
    .B(net7438),
    .Y(_13531_));
 sg13g2_a221oi_1 _22538_ (.B2(\soc_I.clint_I.mtime[51] ),
    .C1(_13531_),
    .B1(net7444),
    .A1(_10660_),
    .Y(_13532_),
    .A2(net7448));
 sg13g2_nand2b_1 _22539_ (.Y(_13533_),
    .B(_13532_),
    .A_N(_13530_));
 sg13g2_o21ai_1 _22540_ (.B1(net8992),
    .Y(_13534_),
    .A1(net8999),
    .A2(_00035_));
 sg13g2_a21oi_1 _22541_ (.A1(\soc_I.spi_div_reg[19] ),
    .A2(net8833),
    .Y(_13535_),
    .B1(_13534_));
 sg13g2_nor2_1 _22542_ (.A(net9251),
    .B(_13535_),
    .Y(_13536_));
 sg13g2_a21oi_2 _22543_ (.B1(net9245),
    .Y(_13537_),
    .A2(_13536_),
    .A1(_13533_));
 sg13g2_o21ai_1 _22544_ (.B1(_13529_),
    .Y(_13538_),
    .A1(_13329_),
    .A2(_13537_));
 sg13g2_inv_1 _22545_ (.Y(_13539_),
    .A(_13538_));
 sg13g2_a22oi_1 _22546_ (.Y(_13540_),
    .B1(_13538_),
    .B2(_13342_),
    .A2(_13528_),
    .A1(_13318_));
 sg13g2_or2_1 _22547_ (.X(_13541_),
    .B(_13540_),
    .A(net8498));
 sg13g2_o21ai_1 _22548_ (.B1(_13541_),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[3] ),
    .A1(_13304_),
    .A2(_13506_));
 sg13g2_nand2_1 _22549_ (.Y(_13542_),
    .A(net9267),
    .B(\soc_I.qqspi_I.rdata[4] ));
 sg13g2_a21oi_1 _22550_ (.A1(_10689_),
    .A2(net7450),
    .Y(_13543_),
    .B1(net8988));
 sg13g2_o21ai_1 _22551_ (.B1(_13543_),
    .Y(_13544_),
    .A1(_00132_),
    .A2(_13223_));
 sg13g2_a221oi_1 _22552_ (.B2(\soc_I.clint_I.mtime[36] ),
    .C1(_13544_),
    .B1(_13224_),
    .A1(_10688_),
    .Y(_13545_),
    .A2(net7446));
 sg13g2_nand3_1 _22553_ (.B(net8960),
    .C(net7491),
    .A(\soc_I.spi0_I.rx_data[4] ),
    .Y(_13546_));
 sg13g2_a21oi_1 _22554_ (.A1(\soc_I.gpio0_I.rdata[4] ),
    .A2(_13205_),
    .Y(_13547_),
    .B1(net9253));
 sg13g2_a22oi_1 _22555_ (.Y(_13548_),
    .B1(_13546_),
    .B2(_13547_),
    .A2(_00129_),
    .A1(net9252));
 sg13g2_o21ai_1 _22556_ (.B1(net8989),
    .Y(_13549_),
    .A1(net8995),
    .A2(_00128_));
 sg13g2_a21oi_1 _22557_ (.A1(net8995),
    .A2(_13548_),
    .Y(_13550_),
    .B1(_13549_));
 sg13g2_nor3_1 _22558_ (.A(net9247),
    .B(_13545_),
    .C(_13550_),
    .Y(_13551_));
 sg13g2_nand2b_1 _22559_ (.Y(_13552_),
    .B(net9190),
    .A_N(\soc_I.rx_uart_i.fifo_i.ram[9][4] ));
 sg13g2_o21ai_1 _22560_ (.B1(_13552_),
    .Y(_13553_),
    .A1(net9190),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[8][4] ));
 sg13g2_mux2_1 _22561_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[10][4] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[11][4] ),
    .S(net9190),
    .X(_13554_));
 sg13g2_o21ai_1 _22562_ (.B1(net8982),
    .Y(_13555_),
    .A1(net9188),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[12][4] ));
 sg13g2_a21oi_1 _22563_ (.A1(net9188),
    .A2(_10679_),
    .Y(_13556_),
    .B1(_13555_));
 sg13g2_nor2b_1 _22564_ (.A(\soc_I.rx_uart_i.fifo_i.ram[15][4] ),
    .B_N(net9192),
    .Y(_13557_));
 sg13g2_o21ai_1 _22565_ (.B1(net9182),
    .Y(_13558_),
    .A1(net9192),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[14][4] ));
 sg13g2_mux4_1 _22566_ (.S0(net9187),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[4][4] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[5][4] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[6][4] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[7][4] ),
    .S1(net9180),
    .X(_13559_));
 sg13g2_nor2_1 _22567_ (.A(net9173),
    .B(_13559_),
    .Y(_13560_));
 sg13g2_o21ai_1 _22568_ (.B1(net9175),
    .Y(_13561_),
    .A1(_13557_),
    .A2(_13558_));
 sg13g2_o21ai_1 _22569_ (.B1(_00002_),
    .Y(_13562_),
    .A1(_13556_),
    .A2(_13561_));
 sg13g2_nor2_1 _22570_ (.A(_13560_),
    .B(_13562_),
    .Y(_13563_));
 sg13g2_mux4_1 _22571_ (.S0(net9187),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[0][4] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[1][4] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[2][4] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[3][4] ),
    .S1(net9183),
    .X(_13564_));
 sg13g2_a21oi_1 _22572_ (.A1(net9181),
    .A2(_13554_),
    .Y(_13565_),
    .B1(_10676_));
 sg13g2_o21ai_1 _22573_ (.B1(_13565_),
    .Y(_13566_),
    .A1(net9181),
    .A2(_13553_));
 sg13g2_o21ai_1 _22574_ (.B1(_13566_),
    .Y(_13567_),
    .A1(net9175),
    .A2(_13564_));
 sg13g2_nor2_1 _22575_ (.A(net8675),
    .B(_13563_),
    .Y(_13568_));
 sg13g2_o21ai_1 _22576_ (.B1(_13568_),
    .Y(_13569_),
    .A1(net9177),
    .A2(_13567_));
 sg13g2_o21ai_1 _22577_ (.B1(_13569_),
    .Y(_13570_),
    .A1(net9241),
    .A2(_13551_));
 sg13g2_o21ai_1 _22578_ (.B1(_13542_),
    .Y(_13571_),
    .A1(_13285_),
    .A2(_13570_));
 sg13g2_o21ai_1 _22579_ (.B1(net9292),
    .Y(_13572_),
    .A1(_00046_),
    .A2(net7424));
 sg13g2_nor2_1 _22580_ (.A(_00048_),
    .B(net7438),
    .Y(_13573_));
 sg13g2_a221oi_1 _22581_ (.B2(\soc_I.clint_I.mtime[60] ),
    .C1(_13573_),
    .B1(net7443),
    .A1(_10663_),
    .Y(_13574_),
    .A2(net7448));
 sg13g2_nand2b_1 _22582_ (.Y(_13575_),
    .B(_13574_),
    .A_N(_13572_));
 sg13g2_a22oi_1 _22583_ (.Y(_13576_),
    .B1(net8835),
    .B2(\soc_I.spi_div_reg[28] ),
    .A2(net9254),
    .A1(_10599_));
 sg13g2_a21oi_2 _22584_ (.B1(net9251),
    .Y(_13577_),
    .A2(_13576_),
    .A1(net8994));
 sg13g2_a21oi_2 _22585_ (.B1(net9242),
    .Y(_13578_),
    .A2(_13577_),
    .A1(_13575_));
 sg13g2_inv_2 _22586_ (.Y(_13579_),
    .A(_13578_));
 sg13g2_a22oi_1 _22587_ (.Y(_13580_),
    .B1(net7361),
    .B2(_13579_),
    .A2(\soc_I.qqspi_I.rdata[28] ),
    .A1(net9271));
 sg13g2_and2_1 _22588_ (.A(net9421),
    .B(_13580_),
    .X(_13581_));
 sg13g2_o21ai_1 _22589_ (.B1(net9290),
    .Y(_13582_),
    .A1(_00091_),
    .A2(net7424));
 sg13g2_nor3_1 _22590_ (.A(_00092_),
    .B(net7467),
    .C(net7465),
    .Y(_13583_));
 sg13g2_nand2_1 _22591_ (.Y(_13584_),
    .A(\soc_I.clint_I.mtime[44] ),
    .B(net7440));
 sg13g2_o21ai_1 _22592_ (.B1(_13584_),
    .Y(_13585_),
    .A1(_00093_),
    .A2(net7437));
 sg13g2_nor3_1 _22593_ (.A(_13582_),
    .B(_13583_),
    .C(_13585_),
    .Y(_13586_));
 sg13g2_o21ai_1 _22594_ (.B1(net8988),
    .Y(_13587_),
    .A1(net8996),
    .A2(_00090_));
 sg13g2_a21oi_2 _22595_ (.B1(_13587_),
    .Y(_13588_),
    .A2(net8832),
    .A1(\soc_I.spi0_I.div[12] ));
 sg13g2_nor3_1 _22596_ (.A(net9246),
    .B(_13586_),
    .C(_13588_),
    .Y(_13589_));
 sg13g2_or2_2 _22597_ (.X(_13590_),
    .B(_13589_),
    .A(net9241));
 sg13g2_a22oi_1 _22598_ (.Y(_13591_),
    .B1(net7362),
    .B2(_13590_),
    .A2(\soc_I.qqspi_I.rdata[12] ),
    .A1(net9269));
 sg13g2_a21oi_1 _22599_ (.A1(_10647_),
    .A2(_13591_),
    .Y(_13592_),
    .B1(_13581_));
 sg13g2_nand2_1 _22600_ (.Y(_13593_),
    .A(_13318_),
    .B(_13592_));
 sg13g2_nand2_1 _22601_ (.Y(_13594_),
    .A(net9270),
    .B(\soc_I.qqspi_I.rdata[20] ));
 sg13g2_nand2b_1 _22602_ (.Y(_13595_),
    .B(net7448),
    .A_N(_00044_));
 sg13g2_nand2b_1 _22603_ (.Y(_13596_),
    .B(net7452),
    .A_N(_00043_));
 sg13g2_a22oi_1 _22604_ (.Y(_13597_),
    .B1(_13229_),
    .B2(_10662_),
    .A2(net7442),
    .A1(\soc_I.clint_I.mtime[52] ));
 sg13g2_nand4_1 _22605_ (.B(_13595_),
    .C(_13596_),
    .A(net9292),
    .Y(_13598_),
    .D(_13597_));
 sg13g2_a22oi_1 _22606_ (.Y(_13599_),
    .B1(net8833),
    .B2(\soc_I.spi_div_reg[20] ),
    .A2(net9254),
    .A1(_10597_));
 sg13g2_a21oi_1 _22607_ (.A1(net8992),
    .A2(_13599_),
    .Y(_13600_),
    .B1(net9249));
 sg13g2_a21oi_1 _22608_ (.A1(_13598_),
    .A2(_13600_),
    .Y(_13601_),
    .B1(net9243));
 sg13g2_o21ai_1 _22609_ (.B1(_13594_),
    .Y(_13602_),
    .A1(_13329_),
    .A2(_13601_));
 sg13g2_inv_1 _22610_ (.Y(_13603_),
    .A(_13602_));
 sg13g2_nand2_1 _22611_ (.Y(_13604_),
    .A(_13342_),
    .B(_13602_));
 sg13g2_a21oi_1 _22612_ (.A1(_13593_),
    .A2(_13604_),
    .Y(_13605_),
    .B1(net8497));
 sg13g2_a21o_2 _22613_ (.A2(_13571_),
    .A1(_13305_),
    .B1(_13605_),
    .X(\soc_I.kianv_I.datapath_unit_I.Data[4] ));
 sg13g2_mux2_1 _22614_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[8][5] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[9][5] ),
    .S(net9192),
    .X(_13606_));
 sg13g2_nand2_1 _22615_ (.Y(_13607_),
    .A(net8982),
    .B(_13606_));
 sg13g2_mux2_1 _22616_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[10][5] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[11][5] ),
    .S(net9190),
    .X(_13608_));
 sg13g2_mux2_1 _22617_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[12][5] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[13][5] ),
    .S(net9189),
    .X(_13609_));
 sg13g2_nand2_1 _22618_ (.Y(_13610_),
    .A(net8982),
    .B(_13609_));
 sg13g2_mux2_1 _22619_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[14][5] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[15][5] ),
    .S(net9188),
    .X(_13611_));
 sg13g2_mux4_1 _22620_ (.S0(net9193),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[0][5] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[1][5] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[2][5] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[3][5] ),
    .S1(net9183),
    .X(_13612_));
 sg13g2_a21oi_1 _22621_ (.A1(net9182),
    .A2(_13608_),
    .Y(_13613_),
    .B1(_10676_));
 sg13g2_a21oi_1 _22622_ (.A1(_13607_),
    .A2(_13613_),
    .Y(_13614_),
    .B1(net9177));
 sg13g2_o21ai_1 _22623_ (.B1(_13614_),
    .Y(_13615_),
    .A1(net9174),
    .A2(_13612_));
 sg13g2_a21oi_1 _22624_ (.A1(net9181),
    .A2(_13611_),
    .Y(_13616_),
    .B1(_10676_));
 sg13g2_mux4_1 _22625_ (.S0(net9185),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[4][5] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[5][5] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[6][5] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[7][5] ),
    .S1(net9179),
    .X(_13617_));
 sg13g2_o21ai_1 _22626_ (.B1(net9177),
    .Y(_13618_),
    .A1(net9174),
    .A2(_13617_));
 sg13g2_a21oi_2 _22627_ (.B1(_13618_),
    .Y(_13619_),
    .A2(_13616_),
    .A1(_13610_));
 sg13g2_nor2_1 _22628_ (.A(net8675),
    .B(_13619_),
    .Y(_13620_));
 sg13g2_o21ai_1 _22629_ (.B1(net9290),
    .Y(_13621_),
    .A1(_00135_),
    .A2(net7424));
 sg13g2_nor3_1 _22630_ (.A(_00136_),
    .B(net7467),
    .C(net7465),
    .Y(_13622_));
 sg13g2_nand2_1 _22631_ (.Y(_13623_),
    .A(\soc_I.clint_I.mtime[37] ),
    .B(net7441));
 sg13g2_o21ai_1 _22632_ (.B1(_13623_),
    .Y(_13624_),
    .A1(_00137_),
    .A2(net7437));
 sg13g2_nor3_1 _22633_ (.A(_13621_),
    .B(_13622_),
    .C(_13624_),
    .Y(_13625_));
 sg13g2_nand3_1 _22634_ (.B(net8960),
    .C(net7491),
    .A(\soc_I.spi0_I.rx_data[5] ),
    .Y(_13626_));
 sg13g2_a21oi_1 _22635_ (.A1(\soc_I.gpio0_I.rdata[5] ),
    .A2(_13205_),
    .Y(_13627_),
    .B1(net9252));
 sg13g2_a22oi_1 _22636_ (.Y(_13628_),
    .B1(_13626_),
    .B2(_13627_),
    .A2(_00134_),
    .A1(net9252));
 sg13g2_o21ai_1 _22637_ (.B1(net8989),
    .Y(_13629_),
    .A1(net8995),
    .A2(_00133_));
 sg13g2_a21oi_1 _22638_ (.A1(net8995),
    .A2(_13628_),
    .Y(_13630_),
    .B1(_13629_));
 sg13g2_nor3_1 _22639_ (.A(net9246),
    .B(_13625_),
    .C(_13630_),
    .Y(_13631_));
 sg13g2_nor2_1 _22640_ (.A(net9240),
    .B(_13631_),
    .Y(_13632_));
 sg13g2_a21oi_2 _22641_ (.B1(_13632_),
    .Y(_13633_),
    .A2(_13620_),
    .A1(_13615_));
 sg13g2_a22oi_1 _22642_ (.Y(_13634_),
    .B1(_13202_),
    .B2(_13633_),
    .A2(\soc_I.qqspi_I.rdata[5] ),
    .A1(net9266));
 sg13g2_nand2b_1 _22643_ (.Y(_13635_),
    .B(net7452),
    .A_N(_00054_));
 sg13g2_nor2_1 _22644_ (.A(_00056_),
    .B(net7438),
    .Y(_13636_));
 sg13g2_a221oi_1 _22645_ (.B2(\soc_I.clint_I.mtime[61] ),
    .C1(_13636_),
    .B1(net7442),
    .A1(_10665_),
    .Y(_13637_),
    .A2(net7447));
 sg13g2_nand3_1 _22646_ (.B(_13635_),
    .C(_13637_),
    .A(net9292),
    .Y(_13638_));
 sg13g2_o21ai_1 _22647_ (.B1(net8994),
    .Y(_13639_),
    .A1(net9000),
    .A2(_00053_));
 sg13g2_a21oi_1 _22648_ (.A1(\soc_I.spi_div_reg[29] ),
    .A2(net8835),
    .Y(_13640_),
    .B1(_13639_));
 sg13g2_nor2_1 _22649_ (.A(net9251),
    .B(_13640_),
    .Y(_13641_));
 sg13g2_a21o_1 _22650_ (.A2(_13641_),
    .A1(_13638_),
    .B1(net9245),
    .X(_13642_));
 sg13g2_a22oi_1 _22651_ (.Y(_13643_),
    .B1(net7361),
    .B2(_13642_),
    .A2(\soc_I.qqspi_I.rdata[29] ),
    .A1(net9271));
 sg13g2_nand2_1 _22652_ (.Y(_13644_),
    .A(net9269),
    .B(\soc_I.qqspi_I.rdata[21] ));
 sg13g2_nand2b_1 _22653_ (.Y(_13645_),
    .B(net7453),
    .A_N(_00050_));
 sg13g2_nand2b_1 _22654_ (.Y(_13646_),
    .B(net7447),
    .A_N(_00051_));
 sg13g2_a22oi_1 _22655_ (.Y(_13647_),
    .B1(_13229_),
    .B2(_10664_),
    .A2(net7442),
    .A1(\soc_I.clint_I.mtime[53] ));
 sg13g2_nand4_1 _22656_ (.B(_13645_),
    .C(_13646_),
    .A(net9292),
    .Y(_13648_),
    .D(_13647_));
 sg13g2_o21ai_1 _22657_ (.B1(net8992),
    .Y(_13649_),
    .A1(net8999),
    .A2(_00049_));
 sg13g2_a21oi_1 _22658_ (.A1(\soc_I.spi_div_reg[21] ),
    .A2(net8833),
    .Y(_13650_),
    .B1(_13649_));
 sg13g2_nor2_1 _22659_ (.A(net9249),
    .B(_13650_),
    .Y(_13651_));
 sg13g2_a21oi_1 _22660_ (.A1(_13648_),
    .A2(_13651_),
    .Y(_13652_),
    .B1(net9243));
 sg13g2_o21ai_1 _22661_ (.B1(_13644_),
    .Y(_13653_),
    .A1(_13329_),
    .A2(_13652_));
 sg13g2_inv_1 _22662_ (.Y(_13654_),
    .A(_13653_));
 sg13g2_nor3_1 _22663_ (.A(_00096_),
    .B(net7467),
    .C(net7465),
    .Y(_13655_));
 sg13g2_nor3_1 _22664_ (.A(_00095_),
    .B(_12955_),
    .C(net7465),
    .Y(_13656_));
 sg13g2_nand2_1 _22665_ (.Y(_13657_),
    .A(\soc_I.clint_I.mtime[45] ),
    .B(net7440));
 sg13g2_o21ai_1 _22666_ (.B1(_13657_),
    .Y(_13658_),
    .A1(_00097_),
    .A2(net7437));
 sg13g2_nor4_1 _22667_ (.A(net8990),
    .B(_13655_),
    .C(_13656_),
    .D(_13658_),
    .Y(_13659_));
 sg13g2_o21ai_1 _22668_ (.B1(net8989),
    .Y(_13660_),
    .A1(net8996),
    .A2(_00094_));
 sg13g2_a21oi_2 _22669_ (.B1(_13660_),
    .Y(_13661_),
    .A2(net8832),
    .A1(\soc_I.spi0_I.div[13] ));
 sg13g2_nor3_2 _22670_ (.A(net9246),
    .B(_13659_),
    .C(_13661_),
    .Y(_13662_));
 sg13g2_o21ai_1 _22671_ (.B1(net8676),
    .Y(_13663_),
    .A1(net9243),
    .A2(_13662_));
 sg13g2_nand2b_1 _22672_ (.Y(_13664_),
    .B(_13663_),
    .A_N(\soc_I.uart_lsr_rdy ));
 sg13g2_nor2_1 _22673_ (.A(\soc_I.tx_uart_i.state[1] ),
    .B(\soc_I.tx_uart_i.state[0] ),
    .Y(_13665_));
 sg13g2_or2_2 _22674_ (.X(_13666_),
    .B(\soc_I.tx_uart_i.state[0] ),
    .A(\soc_I.tx_uart_i.state[1] ));
 sg13g2_a21oi_1 _22675_ (.A1(\soc_I.uart_lsr_rdy ),
    .A2(_13666_),
    .Y(_13667_),
    .B1(_13316_));
 sg13g2_a22oi_1 _22676_ (.Y(_13668_),
    .B1(_13664_),
    .B2(_13667_),
    .A2(\soc_I.qqspi_I.rdata[13] ),
    .A1(net9269));
 sg13g2_nor3_1 _22677_ (.A(net9421),
    .B(_13319_),
    .C(_13668_),
    .Y(_13669_));
 sg13g2_a21oi_1 _22678_ (.A1(_13342_),
    .A2(_13653_),
    .Y(_13670_),
    .B1(_13669_));
 sg13g2_o21ai_1 _22679_ (.B1(_13670_),
    .Y(_13671_),
    .A1(_13331_),
    .A2(_13643_));
 sg13g2_nand2_1 _22680_ (.Y(_13672_),
    .A(net8496),
    .B(_13671_));
 sg13g2_o21ai_1 _22681_ (.B1(_13672_),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[5] ),
    .A1(_13304_),
    .A2(_13634_));
 sg13g2_a21oi_1 _22682_ (.A1(_10691_),
    .A2(net7450),
    .Y(_13673_),
    .B1(net8988));
 sg13g2_o21ai_1 _22683_ (.B1(_13673_),
    .Y(_13674_),
    .A1(_00142_),
    .A2(_13223_));
 sg13g2_a221oi_1 _22684_ (.B2(\soc_I.clint_I.mtime[38] ),
    .C1(_13674_),
    .B1(_13224_),
    .A1(_10690_),
    .Y(_13675_),
    .A2(net7445));
 sg13g2_nand3_1 _22685_ (.B(net8960),
    .C(net7491),
    .A(\soc_I.spi0_I.rx_data[6] ),
    .Y(_13676_));
 sg13g2_a21oi_1 _22686_ (.A1(\soc_I.gpio0_I.rdata[6] ),
    .A2(_13205_),
    .Y(_13677_),
    .B1(net9252));
 sg13g2_a22oi_1 _22687_ (.Y(_13678_),
    .B1(_13676_),
    .B2(_13677_),
    .A2(_00139_),
    .A1(net9252));
 sg13g2_o21ai_1 _22688_ (.B1(net8988),
    .Y(_13679_),
    .A1(net8996),
    .A2(_00138_));
 sg13g2_a21oi_2 _22689_ (.B1(_13679_),
    .Y(_13680_),
    .A2(_13678_),
    .A1(net8995));
 sg13g2_nor3_1 _22690_ (.A(net9246),
    .B(_13675_),
    .C(_13680_),
    .Y(_13681_));
 sg13g2_nor2_1 _22691_ (.A(net9240),
    .B(_13681_),
    .Y(_13682_));
 sg13g2_mux2_1 _22692_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[8][6] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[9][6] ),
    .S(net9191),
    .X(_13683_));
 sg13g2_nor2b_1 _22693_ (.A(\soc_I.rx_uart_i.fifo_i.ram[11][6] ),
    .B_N(net9189),
    .Y(_13684_));
 sg13g2_o21ai_1 _22694_ (.B1(net9181),
    .Y(_13685_),
    .A1(net9189),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[10][6] ));
 sg13g2_o21ai_1 _22695_ (.B1(net8981),
    .Y(_13686_),
    .A1(net9185),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[12][6] ));
 sg13g2_a21oi_1 _22696_ (.A1(net9185),
    .A2(_10680_),
    .Y(_13687_),
    .B1(_13686_));
 sg13g2_nor2b_1 _22697_ (.A(\soc_I.rx_uart_i.fifo_i.ram[15][6] ),
    .B_N(net9185),
    .Y(_13688_));
 sg13g2_o21ai_1 _22698_ (.B1(net9179),
    .Y(_13689_),
    .A1(net9185),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[14][6] ));
 sg13g2_mux4_1 _22699_ (.S0(net9193),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[0][6] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[1][6] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[2][6] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[3][6] ),
    .S1(net9183),
    .X(_13690_));
 sg13g2_nor2_1 _22700_ (.A(net9175),
    .B(_13690_),
    .Y(_13691_));
 sg13g2_o21ai_1 _22701_ (.B1(net9174),
    .Y(_13692_),
    .A1(_13684_),
    .A2(_13685_));
 sg13g2_a21oi_1 _22702_ (.A1(net8981),
    .A2(_13683_),
    .Y(_13693_),
    .B1(_13692_));
 sg13g2_nor3_1 _22703_ (.A(net9177),
    .B(_13691_),
    .C(_13693_),
    .Y(_13694_));
 sg13g2_mux4_1 _22704_ (.S0(net9185),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[4][6] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[5][6] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[6][6] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[7][6] ),
    .S1(net9179),
    .X(_13695_));
 sg13g2_nor2_1 _22705_ (.A(net9172),
    .B(_13695_),
    .Y(_13696_));
 sg13g2_o21ai_1 _22706_ (.B1(net9172),
    .Y(_13697_),
    .A1(_13688_),
    .A2(_13689_));
 sg13g2_o21ai_1 _22707_ (.B1(net9178),
    .Y(_13698_),
    .A1(_13687_),
    .A2(_13697_));
 sg13g2_nor2_2 _22708_ (.A(_13696_),
    .B(_13698_),
    .Y(_13699_));
 sg13g2_nor3_2 _22709_ (.A(net8675),
    .B(_13694_),
    .C(_13699_),
    .Y(_13700_));
 sg13g2_nor2_2 _22710_ (.A(_13682_),
    .B(_13700_),
    .Y(_13701_));
 sg13g2_a22oi_1 _22711_ (.Y(_13702_),
    .B1(_13202_),
    .B2(_13701_),
    .A2(\soc_I.qqspi_I.rdata[6] ),
    .A1(net9267));
 sg13g2_nand2_1 _22712_ (.Y(_13703_),
    .A(net9270),
    .B(\soc_I.qqspi_I.rdata[22] ));
 sg13g2_nand2b_1 _22713_ (.Y(_13704_),
    .B(net7447),
    .A_N(_00059_));
 sg13g2_nand2b_1 _22714_ (.Y(_13705_),
    .B(net7453),
    .A_N(_00058_));
 sg13g2_a22oi_1 _22715_ (.Y(_13706_),
    .B1(_13229_),
    .B2(_10666_),
    .A2(net7442),
    .A1(\soc_I.clint_I.mtime[54] ));
 sg13g2_nand4_1 _22716_ (.B(_13704_),
    .C(_13705_),
    .A(net9293),
    .Y(_13707_),
    .D(_13706_));
 sg13g2_o21ai_1 _22717_ (.B1(net8992),
    .Y(_13708_),
    .A1(net8999),
    .A2(_00057_));
 sg13g2_a21oi_1 _22718_ (.A1(\soc_I.spi_div_reg[22] ),
    .A2(net8833),
    .Y(_13709_),
    .B1(_13708_));
 sg13g2_nor2_1 _22719_ (.A(net9249),
    .B(_13709_),
    .Y(_13710_));
 sg13g2_a21oi_1 _22720_ (.A1(_13707_),
    .A2(_13710_),
    .Y(_13711_),
    .B1(net9243));
 sg13g2_o21ai_1 _22721_ (.B1(_13703_),
    .Y(_13712_),
    .A1(_13329_),
    .A2(_13711_));
 sg13g2_inv_2 _22722_ (.Y(_13713_),
    .A(_13712_));
 sg13g2_and2_1 _22723_ (.A(_13342_),
    .B(_13712_),
    .X(_13714_));
 sg13g2_o21ai_1 _22724_ (.B1(_13221_),
    .Y(_13715_),
    .A1(_00101_),
    .A2(_13223_));
 sg13g2_a21oi_1 _22725_ (.A1(\soc_I.clint_I.mtime[46] ),
    .A2(_13224_),
    .Y(_13716_),
    .B1(_13715_));
 sg13g2_a221oi_1 _22726_ (.B2(_00100_),
    .C1(_13716_),
    .B1(net7445),
    .A1(_00099_),
    .Y(_13717_),
    .A2(net7450));
 sg13g2_nor2_1 _22727_ (.A(net8990),
    .B(_13717_),
    .Y(_13718_));
 sg13g2_o21ai_1 _22728_ (.B1(net8988),
    .Y(_13719_),
    .A1(net8996),
    .A2(_00098_));
 sg13g2_a21oi_2 _22729_ (.B1(_13719_),
    .Y(_13720_),
    .A2(net8832),
    .A1(\soc_I.spi0_I.div[14] ));
 sg13g2_nor3_2 _22730_ (.A(net9246),
    .B(_13718_),
    .C(_13720_),
    .Y(_13721_));
 sg13g2_o21ai_1 _22731_ (.B1(net8676),
    .Y(_13722_),
    .A1(net9243),
    .A2(_13721_));
 sg13g2_nand2b_1 _22732_ (.Y(_13723_),
    .B(_13722_),
    .A_N(\soc_I.uart_lsr_rdy ));
 sg13g2_a22oi_1 _22733_ (.Y(_13724_),
    .B1(_13667_),
    .B2(_13723_),
    .A2(\soc_I.qqspi_I.rdata[14] ),
    .A1(net9269));
 sg13g2_or3_1 _22734_ (.A(net9422),
    .B(_13319_),
    .C(_13724_),
    .X(_13725_));
 sg13g2_a21oi_1 _22735_ (.A1(_10668_),
    .A2(net7452),
    .Y(_13726_),
    .B1(net8994));
 sg13g2_a22oi_1 _22736_ (.Y(_13727_),
    .B1(_13229_),
    .B2(_00064_),
    .A2(net7492),
    .A1(_10400_));
 sg13g2_a22oi_1 _22737_ (.Y(_13728_),
    .B1(_13226_),
    .B2(_13727_),
    .A2(net7449),
    .A1(_10667_));
 sg13g2_o21ai_1 _22738_ (.B1(net8994),
    .Y(_13729_),
    .A1(net9000),
    .A2(_00061_));
 sg13g2_a21oi_1 _22739_ (.A1(\soc_I.spi_div_reg[30] ),
    .A2(net8835),
    .Y(_13730_),
    .B1(_13729_));
 sg13g2_or2_1 _22740_ (.X(_13731_),
    .B(_13730_),
    .A(net9251));
 sg13g2_a21oi_2 _22741_ (.B1(_13731_),
    .Y(_13732_),
    .A2(_13728_),
    .A1(_13726_));
 sg13g2_or2_1 _22742_ (.X(_13733_),
    .B(_13732_),
    .A(net9243));
 sg13g2_a22oi_1 _22743_ (.Y(_13734_),
    .B1(net7361),
    .B2(_13733_),
    .A2(\soc_I.qqspi_I.rdata[30] ),
    .A1(net9266));
 sg13g2_o21ai_1 _22744_ (.B1(_13725_),
    .Y(_13735_),
    .A1(_13331_),
    .A2(_13734_));
 sg13g2_o21ai_1 _22745_ (.B1(net8494),
    .Y(_13736_),
    .A1(_13714_),
    .A2(_13735_));
 sg13g2_o21ai_1 _22746_ (.B1(_13736_),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[6] ),
    .A1(_13304_),
    .A2(_13702_));
 sg13g2_nand2_1 _22747_ (.Y(_13737_),
    .A(net9266),
    .B(\soc_I.qqspi_I.rdata[7] ));
 sg13g2_mux2_1 _22748_ (.A0(\soc_I.rx_uart_i.fifo_i.ram[8][7] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[9][7] ),
    .S(net9191),
    .X(_13738_));
 sg13g2_nor2b_1 _22749_ (.A(\soc_I.rx_uart_i.fifo_i.ram[11][7] ),
    .B_N(net9191),
    .Y(_13739_));
 sg13g2_o21ai_1 _22750_ (.B1(net9181),
    .Y(_13740_),
    .A1(net9191),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[10][7] ));
 sg13g2_o21ai_1 _22751_ (.B1(net8981),
    .Y(_13741_),
    .A1(net9184),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[12][7] ));
 sg13g2_a21oi_1 _22752_ (.A1(net9184),
    .A2(_10681_),
    .Y(_13742_),
    .B1(_13741_));
 sg13g2_nor2b_1 _22753_ (.A(\soc_I.rx_uart_i.fifo_i.ram[15][7] ),
    .B_N(net9189),
    .Y(_13743_));
 sg13g2_o21ai_1 _22754_ (.B1(net9182),
    .Y(_13744_),
    .A1(net9189),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[14][7] ));
 sg13g2_mux4_1 _22755_ (.S0(net9187),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[0][7] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[1][7] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[2][7] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[3][7] ),
    .S1(net9180),
    .X(_13745_));
 sg13g2_nor2_1 _22756_ (.A(net9173),
    .B(_13745_),
    .Y(_13746_));
 sg13g2_o21ai_1 _22757_ (.B1(net9174),
    .Y(_13747_),
    .A1(_13739_),
    .A2(_13740_));
 sg13g2_a21oi_2 _22758_ (.B1(_13747_),
    .Y(_13748_),
    .A2(_13738_),
    .A1(net8982));
 sg13g2_nor3_1 _22759_ (.A(net9177),
    .B(_13746_),
    .C(_13748_),
    .Y(_13749_));
 sg13g2_mux4_1 _22760_ (.S0(net9194),
    .A0(\soc_I.rx_uart_i.fifo_i.ram[4][7] ),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[5][7] ),
    .A2(\soc_I.rx_uart_i.fifo_i.ram[6][7] ),
    .A3(\soc_I.rx_uart_i.fifo_i.ram[7][7] ),
    .S1(net9183),
    .X(_13750_));
 sg13g2_nor2_1 _22761_ (.A(net9175),
    .B(_13750_),
    .Y(_13751_));
 sg13g2_o21ai_1 _22762_ (.B1(net9172),
    .Y(_13752_),
    .A1(_13743_),
    .A2(_13744_));
 sg13g2_o21ai_1 _22763_ (.B1(net9178),
    .Y(_13753_),
    .A1(_13742_),
    .A2(_13752_));
 sg13g2_nor2_1 _22764_ (.A(_13751_),
    .B(_13753_),
    .Y(_13754_));
 sg13g2_or3_1 _22765_ (.A(net8675),
    .B(_13749_),
    .C(_13754_),
    .X(_13755_));
 sg13g2_a21oi_1 _22766_ (.A1(_00146_),
    .A2(net7446),
    .Y(_13756_),
    .B1(net7451));
 sg13g2_a21oi_1 _22767_ (.A1(\soc_I.clint_I.mtime[39] ),
    .A2(net7440),
    .Y(_13757_),
    .B1(net7445));
 sg13g2_o21ai_1 _22768_ (.B1(_13757_),
    .Y(_13758_),
    .A1(_00147_),
    .A2(net7437));
 sg13g2_a221oi_1 _22769_ (.B2(_13758_),
    .C1(net8990),
    .B1(_13756_),
    .A1(_10692_),
    .Y(_13759_),
    .A2(net7450));
 sg13g2_nand2_1 _22770_ (.Y(_13760_),
    .A(\soc_I.gpio0_I.rdata[7] ),
    .B(_13205_));
 sg13g2_nand3_1 _22771_ (.B(_12880_),
    .C(net7492),
    .A(\soc_I.spi0_I.rx_data[7] ),
    .Y(_13761_));
 sg13g2_a21oi_2 _22772_ (.B1(_12878_),
    .Y(_13762_),
    .A2(_13761_),
    .A1(_13760_));
 sg13g2_o21ai_1 _22773_ (.B1(net8989),
    .Y(_13763_),
    .A1(net8996),
    .A2(_00143_));
 sg13g2_nor3_1 _22774_ (.A(net9254),
    .B(_10604_),
    .C(_00144_),
    .Y(_13764_));
 sg13g2_nor3_2 _22775_ (.A(_13762_),
    .B(_13763_),
    .C(_13764_),
    .Y(_13765_));
 sg13g2_nor3_1 _22776_ (.A(net9246),
    .B(_13759_),
    .C(_13765_),
    .Y(_13766_));
 sg13g2_o21ai_1 _22777_ (.B1(_13755_),
    .Y(_13767_),
    .A1(net9241),
    .A2(_13766_));
 sg13g2_o21ai_1 _22778_ (.B1(_13737_),
    .Y(_13768_),
    .A1(_13285_),
    .A2(_13767_));
 sg13g2_a21oi_1 _22779_ (.A1(_00067_),
    .A2(net7447),
    .Y(_13769_),
    .B1(net7453));
 sg13g2_a21oi_1 _22780_ (.A1(\soc_I.clint_I.mtime[55] ),
    .A2(net7442),
    .Y(_13770_),
    .B1(net7448));
 sg13g2_o21ai_1 _22781_ (.B1(_13770_),
    .Y(_13771_),
    .A1(_00068_),
    .A2(net7438));
 sg13g2_a221oi_1 _22782_ (.B2(_13771_),
    .C1(net8993),
    .B1(_13769_),
    .A1(_10669_),
    .Y(_13772_),
    .A2(net7452));
 sg13g2_o21ai_1 _22783_ (.B1(net8992),
    .Y(_13773_),
    .A1(net8999),
    .A2(_00065_));
 sg13g2_a21oi_1 _22784_ (.A1(\soc_I.spi_div_reg[23] ),
    .A2(net8833),
    .Y(_13774_),
    .B1(_13773_));
 sg13g2_nor3_1 _22785_ (.A(net9250),
    .B(_13772_),
    .C(_13774_),
    .Y(_13775_));
 sg13g2_or2_1 _22786_ (.X(_13776_),
    .B(_13775_),
    .A(net9243));
 sg13g2_a22oi_1 _22787_ (.Y(_13777_),
    .B1(net7361),
    .B2(_13776_),
    .A2(\soc_I.qqspi_I.rdata[23] ),
    .A1(net9270));
 sg13g2_nand2_1 _22788_ (.Y(_13778_),
    .A(net9269),
    .B(\soc_I.qqspi_I.rdata[15] ));
 sg13g2_a21oi_1 _22789_ (.A1(_00104_),
    .A2(net7446),
    .Y(_13779_),
    .B1(net7451));
 sg13g2_a21oi_1 _22790_ (.A1(\soc_I.clint_I.mtime[47] ),
    .A2(net7440),
    .Y(_13780_),
    .B1(net7445));
 sg13g2_o21ai_1 _22791_ (.B1(_13780_),
    .Y(_13781_),
    .A1(_00105_),
    .A2(net7437));
 sg13g2_a221oi_1 _22792_ (.B2(_13781_),
    .C1(net8991),
    .B1(_13779_),
    .A1(_10684_),
    .Y(_13782_),
    .A2(net7451));
 sg13g2_o21ai_1 _22793_ (.B1(net8991),
    .Y(_13783_),
    .A1(net8998),
    .A2(_00102_));
 sg13g2_a21oi_2 _22794_ (.B1(_13783_),
    .Y(_13784_),
    .A2(_13207_),
    .A1(\soc_I.spi0_I.div[15] ));
 sg13g2_nor3_1 _22795_ (.A(net9248),
    .B(_13782_),
    .C(_13784_),
    .Y(_13785_));
 sg13g2_nor2_2 _22796_ (.A(net9242),
    .B(_13785_),
    .Y(_13786_));
 sg13g2_o21ai_1 _22797_ (.B1(_13778_),
    .Y(_13787_),
    .A1(_13329_),
    .A2(_13786_));
 sg13g2_o21ai_1 _22798_ (.B1(\soc_I.kianv_I.datapath_unit_I.ADDR_I.q[0] ),
    .Y(_13788_),
    .A1(net9421),
    .A2(_13787_));
 sg13g2_o21ai_1 _22799_ (.B1(_13788_),
    .Y(_13789_),
    .A1(_10647_),
    .A2(_13777_));
 sg13g2_a21oi_1 _22800_ (.A1(_00072_),
    .A2(net7447),
    .Y(_13790_),
    .B1(net7453));
 sg13g2_a21oi_1 _22801_ (.A1(\soc_I.clint_I.mtime[63] ),
    .A2(net7443),
    .Y(_13791_),
    .B1(net7448));
 sg13g2_o21ai_1 _22802_ (.B1(_13791_),
    .Y(_13792_),
    .A1(_00073_),
    .A2(net7439));
 sg13g2_a221oi_1 _22803_ (.B2(_13792_),
    .C1(net8994),
    .B1(_13790_),
    .A1(_10671_),
    .Y(_13793_),
    .A2(net7452));
 sg13g2_or4_2 _22804_ (.A(\soc_I.spi0_I.xfer_cycles[3] ),
    .B(\soc_I.spi0_I.xfer_cycles[2] ),
    .C(\soc_I.spi0_I.xfer_cycles[1] ),
    .D(\soc_I.spi0_I.xfer_cycles[0] ),
    .X(_13794_));
 sg13g2_nor3_2 _22805_ (.A(net4823),
    .B(net4292),
    .C(_13794_),
    .Y(_13795_));
 sg13g2_or3_1 _22806_ (.A(\soc_I.spi0_I.xfer_cycles[5] ),
    .B(\soc_I.spi0_I.xfer_cycles[4] ),
    .C(_13794_),
    .X(_13796_));
 sg13g2_nor4_2 _22807_ (.A(_12878_),
    .B(_12879_),
    .C(net7491),
    .Y(_13797_),
    .D(_13795_));
 sg13g2_o21ai_1 _22808_ (.B1(net8993),
    .Y(_13798_),
    .A1(net9000),
    .A2(_00069_));
 sg13g2_nor3_1 _22809_ (.A(net9254),
    .B(_10604_),
    .C(_00070_),
    .Y(_13799_));
 sg13g2_nor3_2 _22810_ (.A(_13797_),
    .B(_13798_),
    .C(_13799_),
    .Y(_13800_));
 sg13g2_nor3_1 _22811_ (.A(net9251),
    .B(_13793_),
    .C(_13800_),
    .Y(_13801_));
 sg13g2_or2_1 _22812_ (.X(_13802_),
    .B(_13801_),
    .A(net9245));
 sg13g2_a22oi_1 _22813_ (.Y(_13803_),
    .B1(net7361),
    .B2(_13802_),
    .A2(\soc_I.qqspi_I.rdata[31] ),
    .A1(net9268));
 sg13g2_nand3_1 _22814_ (.B(net9422),
    .C(_13803_),
    .A(\soc_I.kianv_I.datapath_unit_I.ADDR_I.q[0] ),
    .Y(_13804_));
 sg13g2_a22oi_1 _22815_ (.Y(_13805_),
    .B1(_13789_),
    .B2(_13804_),
    .A2(_13768_),
    .A1(_13303_));
 sg13g2_nand2b_1 _22816_ (.Y(_13806_),
    .B(_13299_),
    .A_N(_13805_));
 sg13g2_o21ai_1 _22817_ (.B1(_13806_),
    .Y(_13807_),
    .A1(_13341_),
    .A2(_13777_));
 sg13g2_a22oi_1 _22818_ (.Y(_13808_),
    .B1(_13807_),
    .B2(net8496),
    .A2(_13768_),
    .A1(_13302_));
 sg13g2_inv_1 _22819_ (.Y(\soc_I.kianv_I.datapath_unit_I.Data[7] ),
    .A(_13808_));
 sg13g2_nor2b_1 _22820_ (.A(_13805_),
    .B_N(_13289_),
    .Y(_13809_));
 sg13g2_nor2_1 _22821_ (.A(_13330_),
    .B(_13341_),
    .Y(_13810_));
 sg13g2_o21ai_1 _22822_ (.B1(net8493),
    .Y(_13811_),
    .A1(net7336),
    .A2(_13810_));
 sg13g2_o21ai_1 _22823_ (.B1(_13811_),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[8] ),
    .A1(_13301_),
    .A2(_13317_));
 sg13g2_nor2b_1 _22824_ (.A(net8373),
    .B_N(_13398_),
    .Y(_13812_));
 sg13g2_nor3_1 _22825_ (.A(net8498),
    .B(net7336),
    .C(_13812_),
    .Y(_13813_));
 sg13g2_a21oi_2 _22826_ (.B1(_13813_),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[9] ),
    .A2(_13397_),
    .A1(net8498));
 sg13g2_nor2b_1 _22827_ (.A(net8373),
    .B_N(_13462_),
    .Y(_13814_));
 sg13g2_nor3_1 _22828_ (.A(net8498),
    .B(net7336),
    .C(_13814_),
    .Y(_13815_));
 sg13g2_a21oi_2 _22829_ (.B1(_13815_),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[10] ),
    .A2(_13461_),
    .A1(net8497));
 sg13g2_nor2b_1 _22830_ (.A(net8373),
    .B_N(_13528_),
    .Y(_13816_));
 sg13g2_nor3_1 _22831_ (.A(net8497),
    .B(net7336),
    .C(_13816_),
    .Y(_13817_));
 sg13g2_a21oi_1 _22832_ (.A1(net8497),
    .A2(_13527_),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[11] ),
    .B1(_13817_));
 sg13g2_nor2b_1 _22833_ (.A(net8373),
    .B_N(_13592_),
    .Y(_13818_));
 sg13g2_nor3_1 _22834_ (.A(net8497),
    .B(net7336),
    .C(_13818_),
    .Y(_13819_));
 sg13g2_a21oi_2 _22835_ (.B1(_13819_),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[12] ),
    .A2(_13591_),
    .A1(net8497));
 sg13g2_nor2_1 _22836_ (.A(_13341_),
    .B(_13643_),
    .Y(_13820_));
 sg13g2_o21ai_1 _22837_ (.B1(net8494),
    .Y(_13821_),
    .A1(net7336),
    .A2(_13820_));
 sg13g2_o21ai_1 _22838_ (.B1(_13821_),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[13] ),
    .A1(_13301_),
    .A2(_13668_));
 sg13g2_nor2_1 _22839_ (.A(_13341_),
    .B(_13734_),
    .Y(_13822_));
 sg13g2_o21ai_1 _22840_ (.B1(net8494),
    .Y(_13823_),
    .A1(net7336),
    .A2(_13822_));
 sg13g2_o21ai_1 _22841_ (.B1(_13823_),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[14] ),
    .A1(_13301_),
    .A2(_13724_));
 sg13g2_nand2_1 _22842_ (.Y(_13824_),
    .A(_13300_),
    .B(_13787_));
 sg13g2_o21ai_1 _22843_ (.B1(_13824_),
    .Y(_13825_),
    .A1(_13341_),
    .A2(_13803_));
 sg13g2_nor3_1 _22844_ (.A(net8497),
    .B(net7336),
    .C(_13825_),
    .Y(_13826_));
 sg13g2_nor2_1 _22845_ (.A(net8493),
    .B(_13787_),
    .Y(_13827_));
 sg13g2_nor2_1 _22846_ (.A(_13826_),
    .B(_13827_),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[15] ));
 sg13g2_and2_1 _22847_ (.A(_13298_),
    .B(_13825_),
    .X(_13828_));
 sg13g2_o21ai_1 _22848_ (.B1(net8493),
    .Y(_13829_),
    .A1(_13809_),
    .A2(_13828_));
 sg13g2_o21ai_1 _22849_ (.B1(net7335),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[16] ),
    .A1(net8493),
    .A2(_13340_));
 sg13g2_o21ai_1 _22850_ (.B1(net7335),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[17] ),
    .A1(net8493),
    .A2(_13410_));
 sg13g2_o21ai_1 _22851_ (.B1(net7335),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[18] ),
    .A1(net8493),
    .A2(_13473_));
 sg13g2_o21ai_1 _22852_ (.B1(net7335),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[19] ),
    .A1(net8494),
    .A2(_13539_));
 sg13g2_o21ai_1 _22853_ (.B1(net7334),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[20] ),
    .A1(net8495),
    .A2(_13603_));
 sg13g2_o21ai_1 _22854_ (.B1(net7334),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[21] ),
    .A1(net8495),
    .A2(_13654_));
 sg13g2_o21ai_1 _22855_ (.B1(net7334),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[22] ),
    .A1(net8495),
    .A2(_13713_));
 sg13g2_o21ai_1 _22856_ (.B1(net7335),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[23] ),
    .A1(net8494),
    .A2(_13777_));
 sg13g2_o21ai_1 _22857_ (.B1(net7334),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[24] ),
    .A1(net8495),
    .A2(_13330_));
 sg13g2_o21ai_1 _22858_ (.B1(net7334),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[25] ),
    .A1(net8495),
    .A2(_13387_));
 sg13g2_o21ai_1 _22859_ (.B1(net7334),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[26] ),
    .A1(net8495),
    .A2(_13451_));
 sg13g2_o21ai_1 _22860_ (.B1(net7334),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[27] ),
    .A1(net8495),
    .A2(_13516_));
 sg13g2_o21ai_1 _22861_ (.B1(_13829_),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[28] ),
    .A1(net8496),
    .A2(_13580_));
 sg13g2_o21ai_1 _22862_ (.B1(net7334),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[29] ),
    .A1(net8495),
    .A2(_13643_));
 sg13g2_o21ai_1 _22863_ (.B1(net7335),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[30] ),
    .A1(net8496),
    .A2(_13734_));
 sg13g2_o21ai_1 _22864_ (.B1(net7335),
    .Y(\soc_I.kianv_I.datapath_unit_I.Data[31] ),
    .A1(net8493),
    .A2(_13803_));
 sg13g2_nor2_2 _22865_ (.A(_10841_),
    .B(_10861_),
    .Y(_13830_));
 sg13g2_nor2_2 _22866_ (.A(_10841_),
    .B(_10871_),
    .Y(_13831_));
 sg13g2_o21ai_1 _22867_ (.B1(_10874_),
    .Y(_13832_),
    .A1(net9702),
    .A2(_10587_));
 sg13g2_nand2_2 _22868_ (.Y(_13833_),
    .A(_13831_),
    .B(_13832_));
 sg13g2_nor2_1 _22869_ (.A(net9705),
    .B(net9707),
    .Y(_13834_));
 sg13g2_or2_1 _22870_ (.X(_13835_),
    .B(net9707),
    .A(net9705));
 sg13g2_nand2_2 _22871_ (.Y(_13836_),
    .A(_00188_),
    .B(net8959));
 sg13g2_mux2_2 _22872_ (.A0(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[0] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[32] ),
    .S(net8825),
    .X(_13837_));
 sg13g2_nor2_2 _22873_ (.A(net8623),
    .B(_13837_),
    .Y(_13838_));
 sg13g2_nor2_1 _22874_ (.A(_10517_),
    .B(net8963),
    .Y(_13839_));
 sg13g2_a21oi_1 _22875_ (.A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[0] ),
    .A2(net8963),
    .Y(_13840_),
    .B1(_13839_));
 sg13g2_a21oi_2 _22876_ (.B1(_13838_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[0] ),
    .A2(_13840_),
    .A1(net8614));
 sg13g2_nand2_1 _22877_ (.Y(_13841_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[33] ),
    .B(net8820));
 sg13g2_o21ai_1 _22878_ (.B1(_13841_),
    .Y(_13842_),
    .A1(_10619_),
    .A2(net8820));
 sg13g2_nor2_1 _22879_ (.A(net8624),
    .B(_13842_),
    .Y(_13843_));
 sg13g2_nor2_1 _22880_ (.A(_10516_),
    .B(net8967),
    .Y(_13844_));
 sg13g2_a21oi_1 _22881_ (.A1(net5414),
    .A2(net8967),
    .Y(_13845_),
    .B1(_13844_));
 sg13g2_a21oi_1 _22882_ (.A1(net8616),
    .A2(_13845_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[1] ),
    .B1(_13843_));
 sg13g2_nor2_1 _22883_ (.A(_10620_),
    .B(net8820),
    .Y(_13846_));
 sg13g2_a21oi_2 _22884_ (.B1(_13846_),
    .Y(_13847_),
    .A2(net8821),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[34] ));
 sg13g2_mux2_1 _22885_ (.A0(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[2] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[2] ),
    .S(net8967),
    .X(_13848_));
 sg13g2_nand2_1 _22886_ (.Y(_13849_),
    .A(net8616),
    .B(_13848_));
 sg13g2_o21ai_1 _22887_ (.B1(_13849_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[2] ),
    .A1(net8618),
    .A2(_13847_));
 sg13g2_nor2_1 _22888_ (.A(_10621_),
    .B(net8822),
    .Y(_13850_));
 sg13g2_a21oi_2 _22889_ (.B1(_13850_),
    .Y(_13851_),
    .A2(net8822),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[35] ));
 sg13g2_mux2_1 _22890_ (.A0(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[3] ),
    .A1(net5325),
    .S(net8967),
    .X(_13852_));
 sg13g2_nand2_1 _22891_ (.Y(_13853_),
    .A(net8616),
    .B(_13852_));
 sg13g2_o21ai_1 _22892_ (.B1(_13853_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[3] ),
    .A1(net8617),
    .A2(_13851_));
 sg13g2_nor2_1 _22893_ (.A(_10622_),
    .B(net8822),
    .Y(_13854_));
 sg13g2_a21oi_2 _22894_ (.B1(_13854_),
    .Y(_13855_),
    .A2(net8822),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[36] ));
 sg13g2_mux2_1 _22895_ (.A0(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[4] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[4] ),
    .S(net8967),
    .X(_13856_));
 sg13g2_nand2_1 _22896_ (.Y(_13857_),
    .A(net8616),
    .B(_13856_));
 sg13g2_o21ai_1 _22897_ (.B1(_13857_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[4] ),
    .A1(net8616),
    .A2(_13855_));
 sg13g2_mux2_2 _22898_ (.A0(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[5] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[37] ),
    .S(net8820),
    .X(_13858_));
 sg13g2_nor2_1 _22899_ (.A(net8619),
    .B(_13858_),
    .Y(_13859_));
 sg13g2_nor2b_1 _22900_ (.A(net8966),
    .B_N(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[5] ),
    .Y(_13860_));
 sg13g2_a21oi_1 _22901_ (.A1(net5447),
    .A2(net8965),
    .Y(_13861_),
    .B1(_13860_));
 sg13g2_a21oi_1 _22902_ (.A1(net8616),
    .A2(_13861_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[5] ),
    .B1(_13859_));
 sg13g2_mux2_2 _22903_ (.A0(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[6] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[38] ),
    .S(net8820),
    .X(_13862_));
 sg13g2_nor2_1 _22904_ (.A(net8619),
    .B(_13862_),
    .Y(_13863_));
 sg13g2_nor2b_1 _22905_ (.A(net8966),
    .B_N(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[6] ),
    .Y(_13864_));
 sg13g2_a21oi_1 _22906_ (.A1(net5256),
    .A2(net8965),
    .Y(_13865_),
    .B1(_13864_));
 sg13g2_a21oi_1 _22907_ (.A1(net8617),
    .A2(_13865_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[6] ),
    .B1(_13863_));
 sg13g2_mux2_2 _22908_ (.A0(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[7] ),
    .A1(net9206),
    .S(net8820),
    .X(_13866_));
 sg13g2_nor2_1 _22909_ (.A(net8619),
    .B(_13866_),
    .Y(_13867_));
 sg13g2_nor2_1 _22910_ (.A(_10515_),
    .B(net8966),
    .Y(_13868_));
 sg13g2_a21oi_1 _22911_ (.A1(net5283),
    .A2(net8965),
    .Y(_13869_),
    .B1(_13868_));
 sg13g2_a21oi_1 _22912_ (.A1(net8617),
    .A2(_13869_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[7] ),
    .B1(_13867_));
 sg13g2_mux2_2 _22913_ (.A0(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[8] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[40] ),
    .S(net8820),
    .X(_13870_));
 sg13g2_nor2_1 _22914_ (.A(net8619),
    .B(_13870_),
    .Y(_13871_));
 sg13g2_nor2b_1 _22915_ (.A(net8965),
    .B_N(net5310),
    .Y(_13872_));
 sg13g2_a21oi_1 _22916_ (.A1(net5230),
    .A2(net8965),
    .Y(_13873_),
    .B1(_13872_));
 sg13g2_a21oi_1 _22917_ (.A1(net8617),
    .A2(_13873_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[8] ),
    .B1(_13871_));
 sg13g2_nor2_1 _22918_ (.A(_10625_),
    .B(net8821),
    .Y(_13874_));
 sg13g2_a21oi_2 _22919_ (.B1(_13874_),
    .Y(_13875_),
    .A2(net8820),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[41] ));
 sg13g2_mux2_1 _22920_ (.A0(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[9] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[9] ),
    .S(net8967),
    .X(_13876_));
 sg13g2_nand2_1 _22921_ (.Y(_13877_),
    .A(net8616),
    .B(_13876_));
 sg13g2_o21ai_1 _22922_ (.B1(_13877_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[9] ),
    .A1(net8616),
    .A2(_13875_));
 sg13g2_mux2_2 _22923_ (.A0(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[10] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[42] ),
    .S(net8821),
    .X(_13878_));
 sg13g2_nor2_1 _22924_ (.A(net8619),
    .B(_13878_),
    .Y(_13879_));
 sg13g2_nor2b_1 _22925_ (.A(net8966),
    .B_N(net5235),
    .Y(_13880_));
 sg13g2_a21oi_1 _22926_ (.A1(net5224),
    .A2(net8965),
    .Y(_13881_),
    .B1(_13880_));
 sg13g2_a21oi_1 _22927_ (.A1(net8617),
    .A2(_13881_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[10] ),
    .B1(_13879_));
 sg13g2_nor2_1 _22928_ (.A(_10626_),
    .B(net8822),
    .Y(_13882_));
 sg13g2_a21oi_2 _22929_ (.B1(_13882_),
    .Y(_13883_),
    .A2(net8821),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[43] ));
 sg13g2_mux2_1 _22930_ (.A0(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[11] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[11] ),
    .S(net8966),
    .X(_13884_));
 sg13g2_nand2_1 _22931_ (.Y(_13885_),
    .A(net8618),
    .B(_13884_));
 sg13g2_o21ai_1 _22932_ (.B1(_13885_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[11] ),
    .A1(net8618),
    .A2(_13883_));
 sg13g2_nor2_1 _22933_ (.A(_10627_),
    .B(net8821),
    .Y(_13886_));
 sg13g2_a21oi_2 _22934_ (.B1(_13886_),
    .Y(_13887_),
    .A2(net8821),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[44] ));
 sg13g2_mux2_1 _22935_ (.A0(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[12] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[12] ),
    .S(net8965),
    .X(_13888_));
 sg13g2_nand2_1 _22936_ (.Y(_13889_),
    .A(net8624),
    .B(_13888_));
 sg13g2_o21ai_1 _22937_ (.B1(_13889_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[12] ),
    .A1(net8619),
    .A2(_13887_));
 sg13g2_mux2_2 _22938_ (.A0(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[13] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[45] ),
    .S(net8821),
    .X(_13890_));
 sg13g2_nor2_1 _22939_ (.A(net8618),
    .B(_13890_),
    .Y(_13891_));
 sg13g2_nor2b_2 _22940_ (.A(net8968),
    .B_N(net5543),
    .Y(_13892_));
 sg13g2_a21oi_1 _22941_ (.A1(net5520),
    .A2(net8965),
    .Y(_13893_),
    .B1(_13892_));
 sg13g2_a21oi_1 _22942_ (.A1(net8617),
    .A2(_13893_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[13] ),
    .B1(_13891_));
 sg13g2_mux2_2 _22943_ (.A0(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[14] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[46] ),
    .S(net8825),
    .X(_13894_));
 sg13g2_nor2_1 _22944_ (.A(net8623),
    .B(_13894_),
    .Y(_13895_));
 sg13g2_nor2b_1 _22945_ (.A(net8968),
    .B_N(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[14] ),
    .Y(_13896_));
 sg13g2_a21oi_1 _22946_ (.A1(net5573),
    .A2(net8968),
    .Y(_13897_),
    .B1(_13896_));
 sg13g2_a21oi_2 _22947_ (.B1(_13895_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[14] ),
    .A2(_13897_),
    .A1(net8625));
 sg13g2_nor2_1 _22948_ (.A(_10628_),
    .B(net8825),
    .Y(_13898_));
 sg13g2_a21oi_2 _22949_ (.B1(_13898_),
    .Y(_13899_),
    .A2(net8825),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[47] ));
 sg13g2_mux2_1 _22950_ (.A0(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[15] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[15] ),
    .S(net8968),
    .X(_13900_));
 sg13g2_nand2_1 _22951_ (.Y(_13901_),
    .A(net8622),
    .B(_13900_));
 sg13g2_o21ai_1 _22952_ (.B1(_13901_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[15] ),
    .A1(net8622),
    .A2(_13899_));
 sg13g2_mux2_2 _22953_ (.A0(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[16] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[48] ),
    .S(net8825),
    .X(_13902_));
 sg13g2_nor2_1 _22954_ (.A(net8623),
    .B(_13902_),
    .Y(_13903_));
 sg13g2_nor2b_1 _22955_ (.A(net8969),
    .B_N(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[16] ),
    .Y(_13904_));
 sg13g2_a21oi_1 _22956_ (.A1(net5572),
    .A2(net8969),
    .Y(_13905_),
    .B1(_13904_));
 sg13g2_a21oi_2 _22957_ (.B1(_13903_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[16] ),
    .A2(_13905_),
    .A1(net8615));
 sg13g2_nor2_1 _22958_ (.A(_10629_),
    .B(net8825),
    .Y(_13906_));
 sg13g2_a21oi_2 _22959_ (.B1(_13906_),
    .Y(_13907_),
    .A2(net8825),
    .A1(net4367));
 sg13g2_mux2_1 _22960_ (.A0(net5138),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[17] ),
    .S(net8968),
    .X(_13908_));
 sg13g2_nand2_1 _22961_ (.Y(_13909_),
    .A(net8620),
    .B(_13908_));
 sg13g2_o21ai_1 _22962_ (.B1(_13909_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[17] ),
    .A1(net8622),
    .A2(_13907_));
 sg13g2_mux2_1 _22963_ (.A0(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[18] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[50] ),
    .S(net8825),
    .X(_13910_));
 sg13g2_nor2_1 _22964_ (.A(net8623),
    .B(_13910_),
    .Y(_13911_));
 sg13g2_nor2b_1 _22965_ (.A(net8968),
    .B_N(net4999),
    .Y(_13912_));
 sg13g2_a21oi_1 _22966_ (.A1(net5360),
    .A2(net8968),
    .Y(_13913_),
    .B1(_13912_));
 sg13g2_a21oi_1 _22967_ (.A1(net8622),
    .A2(_13913_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[18] ),
    .B1(_13911_));
 sg13g2_mux2_1 _22968_ (.A0(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[19] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[51] ),
    .S(net8824),
    .X(_13914_));
 sg13g2_nor2_1 _22969_ (.A(net8621),
    .B(_13914_),
    .Y(_13915_));
 sg13g2_nor2b_1 _22970_ (.A(net8968),
    .B_N(net5057),
    .Y(_13916_));
 sg13g2_a21oi_1 _22971_ (.A1(net5212),
    .A2(net8969),
    .Y(_13917_),
    .B1(_13916_));
 sg13g2_a21oi_1 _22972_ (.A1(net8621),
    .A2(_13917_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[19] ),
    .B1(_13915_));
 sg13g2_mux2_1 _22973_ (.A0(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[20] ),
    .A1(net4928),
    .S(net8824),
    .X(_13918_));
 sg13g2_nor2_1 _22974_ (.A(net8620),
    .B(_13918_),
    .Y(_13919_));
 sg13g2_nor2b_1 _22975_ (.A(net8970),
    .B_N(net5171),
    .Y(_13920_));
 sg13g2_a21oi_1 _22976_ (.A1(net5463),
    .A2(net8970),
    .Y(_13921_),
    .B1(_13920_));
 sg13g2_a21oi_1 _22977_ (.A1(net8620),
    .A2(_13921_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[20] ),
    .B1(_13919_));
 sg13g2_nor2_1 _22978_ (.A(_10630_),
    .B(net8824),
    .Y(_13922_));
 sg13g2_a21oi_1 _22979_ (.A1(net3860),
    .A2(net8824),
    .Y(_13923_),
    .B1(_13922_));
 sg13g2_mux2_1 _22980_ (.A0(net5420),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[21] ),
    .S(net8969),
    .X(_13924_));
 sg13g2_nand2_1 _22981_ (.Y(_13925_),
    .A(net8615),
    .B(_13924_));
 sg13g2_o21ai_1 _22982_ (.B1(_13925_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[21] ),
    .A1(net8620),
    .A2(_13923_));
 sg13g2_mux2_1 _22983_ (.A0(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[22] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[54] ),
    .S(net8823),
    .X(_13926_));
 sg13g2_nor2_1 _22984_ (.A(net8620),
    .B(_13926_),
    .Y(_13927_));
 sg13g2_nor2b_1 _22985_ (.A(net8970),
    .B_N(net5081),
    .Y(_13928_));
 sg13g2_a21oi_1 _22986_ (.A1(net5248),
    .A2(net8970),
    .Y(_13929_),
    .B1(_13928_));
 sg13g2_a21oi_1 _22987_ (.A1(net8615),
    .A2(_13929_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[22] ),
    .B1(_13927_));
 sg13g2_nor2_1 _22988_ (.A(_10631_),
    .B(net8823),
    .Y(_13930_));
 sg13g2_a21oi_2 _22989_ (.B1(_13930_),
    .Y(_13931_),
    .A2(net8823),
    .A1(net4658));
 sg13g2_mux2_1 _22990_ (.A0(net4408),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[23] ),
    .S(net8970),
    .X(_13932_));
 sg13g2_nand2_1 _22991_ (.Y(_13933_),
    .A(net8615),
    .B(_13932_));
 sg13g2_o21ai_1 _22992_ (.B1(_13933_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[23] ),
    .A1(net8615),
    .A2(_13931_));
 sg13g2_mux2_1 _22993_ (.A0(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[24] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[56] ),
    .S(net8823),
    .X(_13934_));
 sg13g2_nor2_2 _22994_ (.A(net8621),
    .B(_13934_),
    .Y(_13935_));
 sg13g2_nor2b_1 _22995_ (.A(net8963),
    .B_N(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[24] ),
    .Y(_13936_));
 sg13g2_a21oi_1 _22996_ (.A1(net5373),
    .A2(net8963),
    .Y(_13937_),
    .B1(_13936_));
 sg13g2_a21oi_2 _22997_ (.B1(_13935_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[24] ),
    .A2(_13937_),
    .A1(net8614));
 sg13g2_mux2_1 _22998_ (.A0(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[25] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[57] ),
    .S(net8823),
    .X(_13938_));
 sg13g2_nor2_2 _22999_ (.A(net8620),
    .B(_13938_),
    .Y(_13939_));
 sg13g2_nor2b_1 _23000_ (.A(net8963),
    .B_N(net4768),
    .Y(_13940_));
 sg13g2_a21oi_1 _23001_ (.A1(net5315),
    .A2(net8963),
    .Y(_13941_),
    .B1(_13940_));
 sg13g2_a21oi_2 _23002_ (.B1(_13939_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[25] ),
    .A2(_13941_),
    .A1(net8614));
 sg13g2_mux2_1 _23003_ (.A0(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[26] ),
    .A1(net4887),
    .S(net8823),
    .X(_13942_));
 sg13g2_nor2_1 _23004_ (.A(net8621),
    .B(_13942_),
    .Y(_13943_));
 sg13g2_nor2b_1 _23005_ (.A(net8963),
    .B_N(net5545),
    .Y(_13944_));
 sg13g2_a21oi_2 _23006_ (.B1(_13944_),
    .Y(_13945_),
    .A2(net8963),
    .A1(net5504));
 sg13g2_a21oi_1 _23007_ (.A1(net8621),
    .A2(_13945_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[26] ),
    .B1(_13943_));
 sg13g2_mux2_1 _23008_ (.A0(net9205),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[59] ),
    .S(net8823),
    .X(_13946_));
 sg13g2_nor2_2 _23009_ (.A(net8620),
    .B(_13946_),
    .Y(_13947_));
 sg13g2_nor2b_1 _23010_ (.A(net8964),
    .B_N(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[27] ),
    .Y(_13948_));
 sg13g2_a21oi_1 _23011_ (.A1(net5245),
    .A2(net8964),
    .Y(_13949_),
    .B1(_13948_));
 sg13g2_a21oi_2 _23012_ (.B1(_13947_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[27] ),
    .A2(_13949_),
    .A1(net8614));
 sg13g2_mux2_1 _23013_ (.A0(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[28] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[60] ),
    .S(net8823),
    .X(_13950_));
 sg13g2_nor2_2 _23014_ (.A(net8620),
    .B(_13950_),
    .Y(_13951_));
 sg13g2_nor2b_1 _23015_ (.A(net8964),
    .B_N(net4872),
    .Y(_13952_));
 sg13g2_a21oi_1 _23016_ (.A1(net5222),
    .A2(net8964),
    .Y(_13953_),
    .B1(_13952_));
 sg13g2_a21oi_2 _23017_ (.B1(_13951_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[28] ),
    .A2(_13953_),
    .A1(net8614));
 sg13g2_nor2_1 _23018_ (.A(_10632_),
    .B(net8826),
    .Y(_13954_));
 sg13g2_a21oi_2 _23019_ (.B1(_13954_),
    .Y(_13955_),
    .A2(net8824),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[61] ));
 sg13g2_mux2_1 _23020_ (.A0(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[29] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[29] ),
    .S(net8964),
    .X(_13956_));
 sg13g2_nand2_1 _23021_ (.Y(_13957_),
    .A(net8614),
    .B(_13956_));
 sg13g2_o21ai_1 _23022_ (.B1(_13957_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[29] ),
    .A1(net8614),
    .A2(_13955_));
 sg13g2_mux2_2 _23023_ (.A0(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[30] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[62] ),
    .S(net8826),
    .X(_13958_));
 sg13g2_nor2_2 _23024_ (.A(net8615),
    .B(_13958_),
    .Y(_13959_));
 sg13g2_nor2_1 _23025_ (.A(_10514_),
    .B(net8964),
    .Y(_13960_));
 sg13g2_a21oi_1 _23026_ (.A1(net5261),
    .A2(net8971),
    .Y(_13961_),
    .B1(_13960_));
 sg13g2_a21oi_2 _23027_ (.B1(_13959_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[30] ),
    .A2(_13961_),
    .A1(net8625));
 sg13g2_nor2_1 _23028_ (.A(_10634_),
    .B(net8826),
    .Y(_13962_));
 sg13g2_a21oi_2 _23029_ (.B1(_13962_),
    .Y(_13963_),
    .A2(net8826),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[63] ));
 sg13g2_mux2_1 _23030_ (.A0(net5568),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[31] ),
    .S(net8964),
    .X(_13964_));
 sg13g2_nand2_1 _23031_ (.Y(_13965_),
    .A(net8614),
    .B(_13964_));
 sg13g2_o21ai_1 _23032_ (.B1(_13965_),
    .Y(\soc_I.kianv_I.datapath_unit_I.MULExtResult[31] ),
    .A1(net8615),
    .A2(_13963_));
 sg13g2_mux2_2 _23033_ (.A0(\soc_I.spi0_I.cen ),
    .A1(\gpio_uo_out[0] ),
    .S(\gpio_uo_en[0] ),
    .X(uo_out[0]));
 sg13g2_mux2_2 _23034_ (.A0(\soc_I.spi0_I.sclk ),
    .A1(\gpio_uo_out[1] ),
    .S(\gpio_uo_en[1] ),
    .X(uo_out[1]));
 sg13g2_nand2_1 _23035_ (.Y(_13966_),
    .A(\gpio_uo_en[2] ),
    .B(\gpio_uo_out[2] ));
 sg13g2_o21ai_1 _23036_ (.B1(_13966_),
    .Y(uo_out[2]),
    .A1(_10398_),
    .A2(\gpio_uo_en[2] ));
 sg13g2_nand2_1 _23037_ (.Y(_13967_),
    .A(\gpio_uo_en[3] ),
    .B(\gpio_uo_out[3] ));
 sg13g2_o21ai_1 _23038_ (.B1(_13967_),
    .Y(uo_out[3]),
    .A1(\gpio_uo_en[3] ),
    .A2(_10457_));
 sg13g2_mux2_2 _23039_ (.A0(\soc_I.tx_uart_i.tx_out ),
    .A1(\gpio_uo_out[4] ),
    .S(\gpio_uo_en[4] ),
    .X(uo_out[4]));
 sg13g2_nand2_1 _23040_ (.Y(_13968_),
    .A(\gpio_uo_en[5] ),
    .B(\gpio_uo_out[5] ));
 sg13g2_o21ai_1 _23041_ (.B1(_13968_),
    .Y(uo_out[5]),
    .A1(\gpio_uo_en[5] ),
    .A2(_10456_));
 sg13g2_nand2_1 _23042_ (.Y(_13969_),
    .A(\gpio_uo_en[6] ),
    .B(\gpio_uo_out[6] ));
 sg13g2_o21ai_1 _23043_ (.B1(_13969_),
    .Y(uo_out[6]),
    .A1(\gpio_uo_en[6] ),
    .A2(_10455_));
 sg13g2_nand2_1 _23044_ (.Y(_13970_),
    .A(\gpio_uo_en[7] ),
    .B(\gpio_uo_out[7] ));
 sg13g2_o21ai_1 _23045_ (.B1(_13970_),
    .Y(uo_out[7]),
    .A1(\gpio_uo_en[7] ),
    .A2(_10454_));
 sg13g2_nand2b_2 _23046_ (.Y(_13971_),
    .B(net8958),
    .A_N(\soc_I.clint_I.addr[0] ));
 sg13g2_o21ai_1 _23047_ (.B1(net8667),
    .Y(_13972_),
    .A1(net9705),
    .A2(net7668));
 sg13g2_nand2b_2 _23048_ (.Y(_13973_),
    .B(_13971_),
    .A_N(_13972_));
 sg13g2_mux2_2 _23049_ (.A0(_00211_),
    .A1(_00210_),
    .S(net8740),
    .X(_13974_));
 sg13g2_nand2_1 _23050_ (.Y(_13975_),
    .A(net8957),
    .B(_13974_));
 sg13g2_and2_2 _23051_ (.A(_00209_),
    .B(net8734),
    .X(_13976_));
 sg13g2_a21oi_2 _23052_ (.B1(_13976_),
    .Y(_13977_),
    .A2(net8739),
    .A1(_00208_));
 sg13g2_a21o_2 _23053_ (.A2(net8739),
    .A1(_00208_),
    .B1(_13976_),
    .X(_13978_));
 sg13g2_o21ai_1 _23054_ (.B1(_13975_),
    .Y(_13979_),
    .A1(net8957),
    .A2(_13977_));
 sg13g2_nand2_1 _23055_ (.Y(_13980_),
    .A(net7480),
    .B(net7447));
 sg13g2_nor2_2 _23056_ (.A(_13973_),
    .B(_13980_),
    .Y(_13981_));
 sg13g2_nand2_1 _23057_ (.Y(_13982_),
    .A(_13979_),
    .B(net7405));
 sg13g2_o21ai_1 _23058_ (.B1(_13982_),
    .Y(_13983_),
    .A1(net4553),
    .A2(net7405));
 sg13g2_nor2_1 _23059_ (.A(net9003),
    .B(_13983_),
    .Y(_00306_));
 sg13g2_mux2_2 _23060_ (.A0(_00207_),
    .A1(_00206_),
    .S(net8742),
    .X(_13984_));
 sg13g2_nand2_1 _23061_ (.Y(_13985_),
    .A(net8956),
    .B(_13984_));
 sg13g2_mux2_2 _23062_ (.A0(_00205_),
    .A1(_00204_),
    .S(net8743),
    .X(_13986_));
 sg13g2_nand2_1 _23063_ (.Y(_13987_),
    .A(net8958),
    .B(net8613));
 sg13g2_nand2_2 _23064_ (.Y(_13988_),
    .A(_13985_),
    .B(_13987_));
 sg13g2_o21ai_1 _23065_ (.B1(net9308),
    .Y(_13989_),
    .A1(net4386),
    .A2(net7405));
 sg13g2_a21oi_1 _23066_ (.A1(net7405),
    .A2(_13988_),
    .Y(_00307_),
    .B1(_13989_));
 sg13g2_o21ai_1 _23067_ (.B1(net9300),
    .Y(_13990_),
    .A1(net4758),
    .A2(net7405));
 sg13g2_mux2_2 _23068_ (.A0(_00203_),
    .A1(_00202_),
    .S(net8741),
    .X(_13991_));
 sg13g2_mux2_2 _23069_ (.A0(_00201_),
    .A1(_00200_),
    .S(net8740),
    .X(_13992_));
 sg13g2_and2_1 _23070_ (.A(net8958),
    .B(net8611),
    .X(_13993_));
 sg13g2_a21oi_2 _23071_ (.B1(_13993_),
    .Y(_13994_),
    .A2(_13991_),
    .A1(net8956));
 sg13g2_a21o_2 _23072_ (.A2(_13991_),
    .A1(net8956),
    .B1(_13993_),
    .X(_13995_));
 sg13g2_a21oi_1 _23073_ (.A1(net7405),
    .A2(_13995_),
    .Y(_00308_),
    .B1(_13990_));
 sg13g2_o21ai_1 _23074_ (.B1(net9308),
    .Y(_13996_),
    .A1(net4974),
    .A2(net7405));
 sg13g2_and2_1 _23075_ (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[3] ),
    .B(net8742),
    .X(_13997_));
 sg13g2_a21oi_2 _23076_ (.B1(_13997_),
    .Y(_13998_),
    .A2(net8735),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[3] ));
 sg13g2_nand2_1 _23077_ (.Y(_13999_),
    .A(net8959),
    .B(net8550));
 sg13g2_mux2_1 _23078_ (.A0(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[11] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[11] ),
    .S(net8729),
    .X(_14000_));
 sg13g2_o21ai_1 _23079_ (.B1(_13999_),
    .Y(_14001_),
    .A1(net8959),
    .A2(_14000_));
 sg13g2_inv_1 _23080_ (.Y(_14002_),
    .A(_14001_));
 sg13g2_a21oi_1 _23081_ (.A1(net7405),
    .A2(_14001_),
    .Y(_00309_),
    .B1(_13996_));
 sg13g2_mux2_2 _23082_ (.A0(_00199_),
    .A1(_00198_),
    .S(net8740),
    .X(_14003_));
 sg13g2_mux2_1 _23083_ (.A0(_00197_),
    .A1(_00196_),
    .S(net8740),
    .X(_14004_));
 sg13g2_and2_1 _23084_ (.A(net8959),
    .B(net8609),
    .X(_14005_));
 sg13g2_a21oi_2 _23085_ (.B1(_14005_),
    .Y(_14006_),
    .A2(_14003_),
    .A1(net8956));
 sg13g2_a21o_2 _23086_ (.A2(_14003_),
    .A1(net8957),
    .B1(_14005_),
    .X(_14007_));
 sg13g2_nand2_1 _23087_ (.Y(_14008_),
    .A(net7406),
    .B(_14007_));
 sg13g2_o21ai_1 _23088_ (.B1(_14008_),
    .Y(_14009_),
    .A1(net4944),
    .A2(net7406));
 sg13g2_nor2_1 _23089_ (.A(net9004),
    .B(_14009_),
    .Y(_00310_));
 sg13g2_mux2_2 _23090_ (.A0(_00195_),
    .A1(_00194_),
    .S(net8740),
    .X(_14010_));
 sg13g2_mux2_2 _23091_ (.A0(_00193_),
    .A1(_00192_),
    .S(net8741),
    .X(_14011_));
 sg13g2_and2_1 _23092_ (.A(net8959),
    .B(net8607),
    .X(_14012_));
 sg13g2_a21oi_2 _23093_ (.B1(_14012_),
    .Y(_14013_),
    .A2(_14010_),
    .A1(net8956));
 sg13g2_a21o_2 _23094_ (.A2(_14010_),
    .A1(net8956),
    .B1(_14012_),
    .X(_14014_));
 sg13g2_o21ai_1 _23095_ (.B1(net9300),
    .Y(_14015_),
    .A1(net5019),
    .A2(net7406));
 sg13g2_a21oi_1 _23096_ (.A1(net7406),
    .A2(_14014_),
    .Y(_00311_),
    .B1(_14015_));
 sg13g2_mux2_2 _23097_ (.A0(_00191_),
    .A1(_00190_),
    .S(net8744),
    .X(_14016_));
 sg13g2_mux2_2 _23098_ (.A0(_00187_),
    .A1(_00186_),
    .S(net8741),
    .X(_14017_));
 sg13g2_and2_1 _23099_ (.A(net8958),
    .B(net8605),
    .X(_14018_));
 sg13g2_a21oi_2 _23100_ (.B1(_14018_),
    .Y(_14019_),
    .A2(_14016_),
    .A1(net8956));
 sg13g2_a21o_2 _23101_ (.A2(_14016_),
    .A1(net8956),
    .B1(_14018_),
    .X(_14020_));
 sg13g2_nand2_1 _23102_ (.Y(_14021_),
    .A(net7406),
    .B(_14020_));
 sg13g2_o21ai_1 _23103_ (.B1(_14021_),
    .Y(_14022_),
    .A1(net4707),
    .A2(net7406));
 sg13g2_nor2_1 _23104_ (.A(net9004),
    .B(_14022_),
    .Y(_00312_));
 sg13g2_and2_1 _23105_ (.A(\soc_I.kianv_I.datapath_unit_I.A2[7] ),
    .B(net8729),
    .X(_14023_));
 sg13g2_a21oi_2 _23106_ (.B1(_14023_),
    .Y(_14024_),
    .A2(net8739),
    .A1(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[7] ));
 sg13g2_a21o_2 _23107_ (.A2(net8739),
    .A1(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[7] ),
    .B1(_14023_),
    .X(_14025_));
 sg13g2_nor2_1 _23108_ (.A(net8957),
    .B(_14025_),
    .Y(_14026_));
 sg13g2_inv_1 _23109_ (.Y(_14027_),
    .A(_14026_));
 sg13g2_mux2_2 _23110_ (.A0(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[15] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[15] ),
    .S(net8729),
    .X(_14028_));
 sg13g2_o21ai_1 _23111_ (.B1(_14027_),
    .Y(_14029_),
    .A1(net8958),
    .A2(_14028_));
 sg13g2_inv_1 _23112_ (.Y(_14030_),
    .A(_14029_));
 sg13g2_o21ai_1 _23113_ (.B1(net9300),
    .Y(_14031_),
    .A1(net4930),
    .A2(net7406));
 sg13g2_a21oi_1 _23114_ (.A1(net7406),
    .A2(_14029_),
    .Y(_00313_),
    .B1(_14031_));
 sg13g2_o21ai_1 _23115_ (.B1(net8666),
    .Y(_14032_),
    .A1(net9700),
    .A2(\soc_I.clint_I.addr[1] ));
 sg13g2_nand2b_2 _23116_ (.Y(_14033_),
    .B(_13971_),
    .A_N(_14032_));
 sg13g2_nor2_1 _23117_ (.A(_13980_),
    .B(_14033_),
    .Y(_14034_));
 sg13g2_o21ai_1 _23118_ (.B1(net9700),
    .Y(_14035_),
    .A1(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[16] ),
    .A2(net8729));
 sg13g2_a21oi_1 _23119_ (.A1(_10591_),
    .A2(net8732),
    .Y(_14036_),
    .B1(_14035_));
 sg13g2_a21oi_2 _23120_ (.B1(_14036_),
    .Y(_14037_),
    .A2(_13977_),
    .A1(_10465_));
 sg13g2_o21ai_1 _23121_ (.B1(net9315),
    .Y(_14038_),
    .A1(net4710),
    .A2(net7399));
 sg13g2_a21oi_1 _23122_ (.A1(net7399),
    .A2(_14037_),
    .Y(_00314_),
    .B1(_14038_));
 sg13g2_and2_1 _23123_ (.A(\soc_I.kianv_I.datapath_unit_I.A2[17] ),
    .B(net8729),
    .X(_14039_));
 sg13g2_a21oi_2 _23124_ (.B1(_14039_),
    .Y(_14040_),
    .A2(net8739),
    .A1(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[17] ));
 sg13g2_mux2_2 _23125_ (.A0(net8613),
    .A1(_14040_),
    .S(net9700),
    .X(_14041_));
 sg13g2_nand2_1 _23126_ (.Y(_14042_),
    .A(net7399),
    .B(_14041_));
 sg13g2_o21ai_1 _23127_ (.B1(_14042_),
    .Y(_14043_),
    .A1(net4692),
    .A2(net7399));
 sg13g2_nor2_1 _23128_ (.A(net9009),
    .B(_14043_),
    .Y(_00315_));
 sg13g2_and2_1 _23129_ (.A(\soc_I.kianv_I.datapath_unit_I.A2[18] ),
    .B(net8729),
    .X(_14044_));
 sg13g2_a21oi_1 _23130_ (.A1(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[18] ),
    .A2(net8739),
    .Y(_14045_),
    .B1(_14044_));
 sg13g2_mux2_2 _23131_ (.A0(net8611),
    .A1(_14045_),
    .S(net9701),
    .X(_14046_));
 sg13g2_o21ai_1 _23132_ (.B1(net9315),
    .Y(_14047_),
    .A1(net4922),
    .A2(net7399));
 sg13g2_a21oi_1 _23133_ (.A1(net7399),
    .A2(_14046_),
    .Y(_00316_),
    .B1(_14047_));
 sg13g2_nand2_1 _23134_ (.Y(_14048_),
    .A(\soc_I.kianv_I.datapath_unit_I.A2[19] ),
    .B(net8731));
 sg13g2_a21oi_1 _23135_ (.A1(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[19] ),
    .A2(net8739),
    .Y(_14049_),
    .B1(_10465_));
 sg13g2_a22oi_1 _23136_ (.Y(_14050_),
    .B1(_14048_),
    .B2(_14049_),
    .A2(net8550),
    .A1(_10465_));
 sg13g2_inv_4 _23137_ (.A(_14050_),
    .Y(_14051_));
 sg13g2_nand2_1 _23138_ (.Y(_14052_),
    .A(net7399),
    .B(_14051_));
 sg13g2_o21ai_1 _23139_ (.B1(_14052_),
    .Y(_14053_),
    .A1(net4749),
    .A2(net7399));
 sg13g2_nor2_1 _23140_ (.A(net9009),
    .B(_14053_),
    .Y(_00317_));
 sg13g2_and2_1 _23141_ (.A(\soc_I.kianv_I.datapath_unit_I.A2[20] ),
    .B(net8734),
    .X(_14054_));
 sg13g2_a21oi_1 _23142_ (.A1(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[20] ),
    .A2(net8740),
    .Y(_14055_),
    .B1(_14054_));
 sg13g2_mux2_2 _23143_ (.A0(net8609),
    .A1(_14055_),
    .S(net9703),
    .X(_14056_));
 sg13g2_o21ai_1 _23144_ (.B1(net9318),
    .Y(_14057_),
    .A1(net4859),
    .A2(net7401));
 sg13g2_a21oi_1 _23145_ (.A1(net7404),
    .A2(_14056_),
    .Y(_00318_),
    .B1(_14057_));
 sg13g2_and2_1 _23146_ (.A(\soc_I.kianv_I.datapath_unit_I.A2[21] ),
    .B(net8734),
    .X(_14058_));
 sg13g2_a21oi_2 _23147_ (.B1(_14058_),
    .Y(_14059_),
    .A2(net8740),
    .A1(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[21] ));
 sg13g2_mux2_2 _23148_ (.A0(net8607),
    .A1(_14059_),
    .S(net9701),
    .X(_14060_));
 sg13g2_nand2_1 _23149_ (.Y(_14061_),
    .A(net7400),
    .B(_14060_));
 sg13g2_o21ai_1 _23150_ (.B1(_14061_),
    .Y(_14062_),
    .A1(net5030),
    .A2(net7400));
 sg13g2_nor2_1 _23151_ (.A(net9012),
    .B(_14062_),
    .Y(_00319_));
 sg13g2_and2_1 _23152_ (.A(\soc_I.kianv_I.datapath_unit_I.A2[22] ),
    .B(net8734),
    .X(_14063_));
 sg13g2_a21oi_1 _23153_ (.A1(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[22] ),
    .A2(net8740),
    .Y(_14064_),
    .B1(_14063_));
 sg13g2_mux2_2 _23154_ (.A0(_14017_),
    .A1(_14064_),
    .S(net9703),
    .X(_14065_));
 sg13g2_o21ai_1 _23155_ (.B1(net9319),
    .Y(_14066_),
    .A1(net5032),
    .A2(net7400));
 sg13g2_a21oi_1 _23156_ (.A1(net7400),
    .A2(_14065_),
    .Y(_00320_),
    .B1(_14066_));
 sg13g2_nand2_1 _23157_ (.Y(_14067_),
    .A(\soc_I.kianv_I.datapath_unit_I.A2[23] ),
    .B(net8729));
 sg13g2_a21oi_2 _23158_ (.B1(_10465_),
    .Y(_14068_),
    .A2(net8739),
    .A1(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[23] ));
 sg13g2_a22oi_1 _23159_ (.Y(_14069_),
    .B1(_14067_),
    .B2(_14068_),
    .A2(_14024_),
    .A1(_10465_));
 sg13g2_inv_4 _23160_ (.A(_14069_),
    .Y(_14070_));
 sg13g2_nand2_1 _23161_ (.Y(_14071_),
    .A(net7400),
    .B(_14070_));
 sg13g2_o21ai_1 _23162_ (.B1(_14071_),
    .Y(_14072_),
    .A1(net4849),
    .A2(net7401));
 sg13g2_nor2_1 _23163_ (.A(net9010),
    .B(_14072_),
    .Y(_00321_));
 sg13g2_and2_1 _23164_ (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[24] ),
    .B(net8742),
    .X(_14073_));
 sg13g2_a21oi_2 _23165_ (.B1(_14073_),
    .Y(_14074_),
    .A2(net8735),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[24] ));
 sg13g2_a22oi_1 _23166_ (.Y(_14075_),
    .B1(_14074_),
    .B2(net9705),
    .A2(_13974_),
    .A1(_10915_));
 sg13g2_o21ai_1 _23167_ (.B1(_14075_),
    .Y(_14076_),
    .A1(net8957),
    .A2(_13977_));
 sg13g2_nand2_1 _23168_ (.Y(_14077_),
    .A(net7400),
    .B(_14076_));
 sg13g2_o21ai_1 _23169_ (.B1(_14077_),
    .Y(_14078_),
    .A1(net4694),
    .A2(net7401));
 sg13g2_nor2_1 _23170_ (.A(net9010),
    .B(_14078_),
    .Y(_00322_));
 sg13g2_and2_1 _23171_ (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[25] ),
    .B(net8741),
    .X(_14079_));
 sg13g2_a21oi_2 _23172_ (.B1(_14079_),
    .Y(_14080_),
    .A2(net8737),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[25] ));
 sg13g2_a22oi_1 _23173_ (.Y(_14081_),
    .B1(_14080_),
    .B2(net9705),
    .A2(_13984_),
    .A1(net8962));
 sg13g2_nand2_2 _23174_ (.Y(_14082_),
    .A(_13987_),
    .B(_14081_));
 sg13g2_o21ai_1 _23175_ (.B1(net9319),
    .Y(_14083_),
    .A1(net5101),
    .A2(net7400));
 sg13g2_a21oi_1 _23176_ (.A1(net7400),
    .A2(_14082_),
    .Y(_00323_),
    .B1(_14083_));
 sg13g2_o21ai_1 _23177_ (.B1(net9328),
    .Y(_14084_),
    .A1(net4919),
    .A2(net7403));
 sg13g2_and2_1 _23178_ (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[26] ),
    .B(net8741),
    .X(_14085_));
 sg13g2_a21oi_2 _23179_ (.B1(_14085_),
    .Y(_14086_),
    .A2(net8736),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[26] ));
 sg13g2_a22oi_1 _23180_ (.Y(_14087_),
    .B1(_14086_),
    .B2(net9700),
    .A2(_13991_),
    .A1(net8962));
 sg13g2_nand2b_2 _23181_ (.Y(_14088_),
    .B(_14087_),
    .A_N(_13993_));
 sg13g2_a21oi_1 _23182_ (.A1(net7402),
    .A2(_14088_),
    .Y(_00324_),
    .B1(_14084_));
 sg13g2_and2_1 _23183_ (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[27] ),
    .B(net8743),
    .X(_14089_));
 sg13g2_a21oi_2 _23184_ (.B1(_14089_),
    .Y(_14090_),
    .A2(net8738),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[27] ));
 sg13g2_o21ai_1 _23185_ (.B1(_13999_),
    .Y(_14091_),
    .A1(_10916_),
    .A2(_14000_));
 sg13g2_a21o_2 _23186_ (.A2(_14090_),
    .A1(net9701),
    .B1(_14091_),
    .X(_14092_));
 sg13g2_nand2_1 _23187_ (.Y(_14093_),
    .A(net7402),
    .B(_14092_));
 sg13g2_o21ai_1 _23188_ (.B1(_14093_),
    .Y(_14094_),
    .A1(net4831),
    .A2(net7403));
 sg13g2_nor2_1 _23189_ (.A(net9010),
    .B(_14094_),
    .Y(_00325_));
 sg13g2_o21ai_1 _23190_ (.B1(net9327),
    .Y(_14095_),
    .A1(net4829),
    .A2(net7402));
 sg13g2_and2_1 _23191_ (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[28] ),
    .B(net8743),
    .X(_14096_));
 sg13g2_a21oi_2 _23192_ (.B1(_14096_),
    .Y(_14097_),
    .A2(net8735),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[28] ));
 sg13g2_a22oi_1 _23193_ (.Y(_14098_),
    .B1(_14097_),
    .B2(net9700),
    .A2(_14003_),
    .A1(net8962));
 sg13g2_nand2b_2 _23194_ (.Y(_14099_),
    .B(_14098_),
    .A_N(_14005_));
 sg13g2_a21oi_1 _23195_ (.A1(net7402),
    .A2(_14099_),
    .Y(_00326_),
    .B1(_14095_));
 sg13g2_nand2_1 _23196_ (.Y(_14100_),
    .A(\soc_I.kianv_I.datapath_unit_I.A2[29] ),
    .B(net8735));
 sg13g2_nand2_1 _23197_ (.Y(_14101_),
    .A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[29] ),
    .B(net8742));
 sg13g2_nand3_1 _23198_ (.B(_14100_),
    .C(_14101_),
    .A(net9703),
    .Y(_14102_));
 sg13g2_a21oi_1 _23199_ (.A1(net8962),
    .A2(_14010_),
    .Y(_14103_),
    .B1(_14012_));
 sg13g2_nand2_2 _23200_ (.Y(_14104_),
    .A(_14102_),
    .B(_14103_));
 sg13g2_inv_1 _23201_ (.Y(_14105_),
    .A(_14104_));
 sg13g2_nand2_1 _23202_ (.Y(_14106_),
    .A(net7402),
    .B(_14104_));
 sg13g2_o21ai_1 _23203_ (.B1(_14106_),
    .Y(_14107_),
    .A1(net4916),
    .A2(net7402));
 sg13g2_nor2_1 _23204_ (.A(net9011),
    .B(_14107_),
    .Y(_00327_));
 sg13g2_and2_1 _23205_ (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[30] ),
    .B(net8744),
    .X(_14108_));
 sg13g2_a21oi_2 _23206_ (.B1(_14108_),
    .Y(_14109_),
    .A2(net8730),
    .A1(\soc_I.kianv_I.datapath_unit_I.A2[30] ));
 sg13g2_a22oi_1 _23207_ (.Y(_14110_),
    .B1(_14109_),
    .B2(net9700),
    .A2(_14016_),
    .A1(net8962));
 sg13g2_nand2b_2 _23208_ (.Y(_14111_),
    .B(_14110_),
    .A_N(_14018_));
 sg13g2_o21ai_1 _23209_ (.B1(net9328),
    .Y(_14112_),
    .A1(net5055),
    .A2(net7403));
 sg13g2_a21oi_1 _23210_ (.A1(net7403),
    .A2(_14111_),
    .Y(_00328_),
    .B1(_14112_));
 sg13g2_o21ai_1 _23211_ (.B1(net9701),
    .Y(_14113_),
    .A1(_10507_),
    .A2(net8729));
 sg13g2_a21oi_1 _23212_ (.A1(\soc_I.kianv_I.datapath_unit_I.A2[31] ),
    .A2(net8732),
    .Y(_14114_),
    .B1(_14113_));
 sg13g2_nor2_1 _23213_ (.A(_10916_),
    .B(_14028_),
    .Y(_14115_));
 sg13g2_or3_2 _23214_ (.A(_14026_),
    .B(_14114_),
    .C(_14115_),
    .X(_14116_));
 sg13g2_nand2_1 _23215_ (.Y(_14117_),
    .A(net7402),
    .B(_14116_));
 sg13g2_o21ai_1 _23216_ (.B1(_14117_),
    .Y(_14118_),
    .A1(net5137),
    .A2(net7402));
 sg13g2_nor2_1 _23217_ (.A(net9013),
    .B(_14118_),
    .Y(_00329_));
 sg13g2_nand2_1 _23218_ (.Y(_14119_),
    .A(net5106),
    .B(_13236_));
 sg13g2_a21oi_1 _23219_ (.A1(\soc_I.rx_uart_i.fifo_i.cnt[4] ),
    .A2(_13236_),
    .Y(_14120_),
    .B1(_10397_));
 sg13g2_nand2_2 _23220_ (.Y(_14121_),
    .A(\soc_I.rx_uart_i.ready ),
    .B(_14119_));
 sg13g2_nor3_2 _23221_ (.A(\soc_I.rx_uart_i.fifo_i.wr_ptr[1] ),
    .B(\soc_I.rx_uart_i.fifo_i.wr_ptr[0] ),
    .C(_14121_),
    .Y(_14122_));
 sg13g2_nor2b_2 _23222_ (.A(\soc_I.rx_uart_i.fifo_i.wr_ptr[3] ),
    .B_N(\soc_I.rx_uart_i.fifo_i.wr_ptr[2] ),
    .Y(_14123_));
 sg13g2_nand2_1 _23223_ (.Y(_14124_),
    .A(_14122_),
    .B(_14123_));
 sg13g2_nand2_1 _23224_ (.Y(_14125_),
    .A(net2652),
    .B(net8548));
 sg13g2_o21ai_1 _23225_ (.B1(_14125_),
    .Y(_00330_),
    .A1(net9170),
    .A2(net8548));
 sg13g2_mux2_1 _23226_ (.A0(net9289),
    .A1(net4136),
    .S(net8548),
    .X(_00331_));
 sg13g2_mux2_1 _23227_ (.A0(net9287),
    .A1(net3941),
    .S(net8548),
    .X(_00332_));
 sg13g2_mux2_1 _23228_ (.A0(net9284),
    .A1(net4074),
    .S(net8548),
    .X(_00333_));
 sg13g2_mux2_1 _23229_ (.A0(net9283),
    .A1(net4082),
    .S(_14124_),
    .X(_00334_));
 sg13g2_mux2_1 _23230_ (.A0(net9281),
    .A1(net3921),
    .S(net8548),
    .X(_00335_));
 sg13g2_mux2_1 _23231_ (.A0(net9277),
    .A1(net4253),
    .S(net8548),
    .X(_00336_));
 sg13g2_mux2_1 _23232_ (.A0(net9276),
    .A1(net4182),
    .S(net8548),
    .X(_00337_));
 sg13g2_nor2_2 _23233_ (.A(_10467_),
    .B(\soc_I.kianv_I.Instr[7] ),
    .Y(_14126_));
 sg13g2_nor2_2 _23234_ (.A(net9709),
    .B(_00185_),
    .Y(_14127_));
 sg13g2_nor2_2 _23235_ (.A(_10984_),
    .B(_12465_),
    .Y(_14128_));
 sg13g2_a21oi_1 _23236_ (.A1(_12607_),
    .A2(net8961),
    .Y(_14129_),
    .B1(_14128_));
 sg13g2_nor3_2 _23237_ (.A(net9709),
    .B(net9710),
    .C(_00185_),
    .Y(_14130_));
 sg13g2_nand3_1 _23238_ (.B(net8371),
    .C(_14130_),
    .A(_14126_),
    .Y(_14131_));
 sg13g2_nand2_1 _23239_ (.Y(_14132_),
    .A(net2769),
    .B(net8243));
 sg13g2_o21ai_1 _23240_ (.B1(_14132_),
    .Y(_00338_),
    .A1(net7488),
    .A2(net8243));
 sg13g2_nand2_1 _23241_ (.Y(_14133_),
    .A(net2832),
    .B(net8243));
 sg13g2_o21ai_1 _23242_ (.B1(_14133_),
    .Y(_00339_),
    .A1(net7667),
    .A2(net8243));
 sg13g2_nand2_1 _23243_ (.Y(_14134_),
    .A(net3232),
    .B(net8243));
 sg13g2_o21ai_1 _23244_ (.B1(_14134_),
    .Y(_00340_),
    .A1(net7613),
    .A2(net8243));
 sg13g2_nand2_1 _23245_ (.Y(_14135_),
    .A(net2916),
    .B(net8241));
 sg13g2_o21ai_1 _23246_ (.B1(_14135_),
    .Y(_00341_),
    .A1(net7611),
    .A2(net8241));
 sg13g2_nand2_1 _23247_ (.Y(_14136_),
    .A(net2770),
    .B(net8238));
 sg13g2_o21ai_1 _23248_ (.B1(_14136_),
    .Y(_00342_),
    .A1(net7586),
    .A2(net8238));
 sg13g2_nand2_1 _23249_ (.Y(_14137_),
    .A(net2743),
    .B(net8238));
 sg13g2_o21ai_1 _23250_ (.B1(_14137_),
    .Y(_00343_),
    .A1(net7598),
    .A2(net8238));
 sg13g2_nand2_1 _23251_ (.Y(_14138_),
    .A(net2788),
    .B(net8240));
 sg13g2_o21ai_1 _23252_ (.B1(_14138_),
    .Y(_00344_),
    .A1(net7594),
    .A2(net8240));
 sg13g2_nand2_1 _23253_ (.Y(_14139_),
    .A(net2765),
    .B(net8233));
 sg13g2_o21ai_1 _23254_ (.B1(_14139_),
    .Y(_00345_),
    .A1(net7602),
    .A2(net8233));
 sg13g2_nand2_1 _23255_ (.Y(_14140_),
    .A(net2810),
    .B(net8239));
 sg13g2_o21ai_1 _23256_ (.B1(_14140_),
    .Y(_00346_),
    .A1(net7562),
    .A2(net8239));
 sg13g2_nand2_1 _23257_ (.Y(_14141_),
    .A(net2762),
    .B(net8242));
 sg13g2_o21ai_1 _23258_ (.B1(_14141_),
    .Y(_00347_),
    .A1(net7576),
    .A2(net8242));
 sg13g2_nand2_1 _23259_ (.Y(_14142_),
    .A(net2980),
    .B(net8240));
 sg13g2_o21ai_1 _23260_ (.B1(_14142_),
    .Y(_00348_),
    .A1(net7550),
    .A2(net8240));
 sg13g2_nand2_1 _23261_ (.Y(_14143_),
    .A(net2851),
    .B(net8233));
 sg13g2_o21ai_1 _23262_ (.B1(_14143_),
    .Y(_00349_),
    .A1(net7568),
    .A2(net8233));
 sg13g2_nand2_1 _23263_ (.Y(_14144_),
    .A(net2750),
    .B(net8240));
 sg13g2_o21ai_1 _23264_ (.B1(_14144_),
    .Y(_00350_),
    .A1(net7543),
    .A2(net8240));
 sg13g2_nand2_1 _23265_ (.Y(_14145_),
    .A(net2811),
    .B(net8242));
 sg13g2_o21ai_1 _23266_ (.B1(_14145_),
    .Y(_00351_),
    .A1(net7552),
    .A2(net8242));
 sg13g2_nand2_1 _23267_ (.Y(_14146_),
    .A(net2701),
    .B(net8237));
 sg13g2_o21ai_1 _23268_ (.B1(_14146_),
    .Y(_00352_),
    .A1(net7585),
    .A2(net8237));
 sg13g2_nand2_1 _23269_ (.Y(_14147_),
    .A(net3469),
    .B(net8234));
 sg13g2_o21ai_1 _23270_ (.B1(_14147_),
    .Y(_00353_),
    .A1(net7564),
    .A2(net8234));
 sg13g2_nand2_1 _23271_ (.Y(_14148_),
    .A(net3056),
    .B(net8233));
 sg13g2_o21ai_1 _23272_ (.B1(_14148_),
    .Y(_00354_),
    .A1(net7525),
    .A2(net8233));
 sg13g2_nand2_1 _23273_ (.Y(_14149_),
    .A(net2933),
    .B(net8233));
 sg13g2_o21ai_1 _23274_ (.B1(_14149_),
    .Y(_00355_),
    .A1(net7534),
    .A2(net8233));
 sg13g2_nand2_1 _23275_ (.Y(_14150_),
    .A(net3377),
    .B(net8234));
 sg13g2_o21ai_1 _23276_ (.B1(_14150_),
    .Y(_00356_),
    .A1(net7528),
    .A2(net8234));
 sg13g2_nand2_1 _23277_ (.Y(_14151_),
    .A(net2988),
    .B(net8236));
 sg13g2_o21ai_1 _23278_ (.B1(_14151_),
    .Y(_00357_),
    .A1(net7518),
    .A2(net8236));
 sg13g2_nand2_1 _23279_ (.Y(_14152_),
    .A(net2695),
    .B(net8239));
 sg13g2_o21ai_1 _23280_ (.B1(_14152_),
    .Y(_00358_),
    .A1(net7505),
    .A2(net8239));
 sg13g2_nand2_1 _23281_ (.Y(_14153_),
    .A(net2689),
    .B(net8238));
 sg13g2_o21ai_1 _23282_ (.B1(_14153_),
    .Y(_00359_),
    .A1(net7513),
    .A2(net8238));
 sg13g2_nand2_1 _23283_ (.Y(_14154_),
    .A(net3289),
    .B(net8241));
 sg13g2_o21ai_1 _23284_ (.B1(_14154_),
    .Y(_00360_),
    .A1(net7496),
    .A2(net8241));
 sg13g2_nand2_1 _23285_ (.Y(_14155_),
    .A(net2723),
    .B(net8235));
 sg13g2_o21ai_1 _23286_ (.B1(_14155_),
    .Y(_00361_),
    .A1(net7502),
    .A2(net8235));
 sg13g2_nand2_1 _23287_ (.Y(_14156_),
    .A(net2737),
    .B(net8238));
 sg13g2_o21ai_1 _23288_ (.B1(_14156_),
    .Y(_00362_),
    .A1(net7644),
    .A2(net8238));
 sg13g2_nand2_1 _23289_ (.Y(_14157_),
    .A(net2763),
    .B(net8243));
 sg13g2_o21ai_1 _23290_ (.B1(_14157_),
    .Y(_00363_),
    .A1(net7650),
    .A2(net8243));
 sg13g2_nand2_1 _23291_ (.Y(_14158_),
    .A(net3293),
    .B(net8240));
 sg13g2_o21ai_1 _23292_ (.B1(_14158_),
    .Y(_00364_),
    .A1(net7654),
    .A2(net8240));
 sg13g2_nand2_1 _23293_ (.Y(_14159_),
    .A(net2801),
    .B(net8236));
 sg13g2_o21ai_1 _23294_ (.B1(_14159_),
    .Y(_00365_),
    .A1(net7658),
    .A2(net8236));
 sg13g2_nand2_1 _23295_ (.Y(_14160_),
    .A(net2793),
    .B(net8236));
 sg13g2_o21ai_1 _23296_ (.B1(_14160_),
    .Y(_00366_),
    .A1(net7636),
    .A2(net8236));
 sg13g2_nand2_1 _23297_ (.Y(_14161_),
    .A(net3060),
    .B(net8239));
 sg13g2_o21ai_1 _23298_ (.B1(_14161_),
    .Y(_00367_),
    .A1(net7625),
    .A2(net8239));
 sg13g2_nand2_1 _23299_ (.Y(_14162_),
    .A(net3379),
    .B(net8236));
 sg13g2_o21ai_1 _23300_ (.B1(_14162_),
    .Y(_00368_),
    .A1(net7621),
    .A2(net8236));
 sg13g2_nand2_1 _23301_ (.Y(_14163_),
    .A(net3063),
    .B(net8235));
 sg13g2_o21ai_1 _23302_ (.B1(_14163_),
    .Y(_00369_),
    .A1(net7631),
    .A2(net8235));
 sg13g2_nand2b_1 _23303_ (.Y(_14164_),
    .B(net9711),
    .A_N(\soc_I.kianv_I.Instr[9] ));
 sg13g2_nor2_2 _23304_ (.A(net9709),
    .B(_14164_),
    .Y(_14165_));
 sg13g2_nand3_1 _23305_ (.B(net8372),
    .C(_14165_),
    .A(_14126_),
    .Y(_14166_));
 sg13g2_nand2_1 _23306_ (.Y(_14167_),
    .A(net3333),
    .B(net8231));
 sg13g2_o21ai_1 _23307_ (.B1(_14167_),
    .Y(_00370_),
    .A1(net7489),
    .A2(net8231));
 sg13g2_nand2_1 _23308_ (.Y(_14168_),
    .A(net3303),
    .B(net8231));
 sg13g2_o21ai_1 _23309_ (.B1(_14168_),
    .Y(_00371_),
    .A1(net7663),
    .A2(net8231));
 sg13g2_nand2_1 _23310_ (.Y(_14169_),
    .A(net3240),
    .B(net8231));
 sg13g2_o21ai_1 _23311_ (.B1(_14169_),
    .Y(_00372_),
    .A1(net7612),
    .A2(net8231));
 sg13g2_nand2_1 _23312_ (.Y(_14170_),
    .A(net3345),
    .B(net8229));
 sg13g2_o21ai_1 _23313_ (.B1(_14170_),
    .Y(_00373_),
    .A1(net7610),
    .A2(net8229));
 sg13g2_nand2_1 _23314_ (.Y(_14171_),
    .A(net3298),
    .B(net8226));
 sg13g2_o21ai_1 _23315_ (.B1(_14171_),
    .Y(_00374_),
    .A1(net7588),
    .A2(net8226));
 sg13g2_nand2_1 _23316_ (.Y(_14172_),
    .A(net2758),
    .B(net8226));
 sg13g2_o21ai_1 _23317_ (.B1(_14172_),
    .Y(_00375_),
    .A1(net7597),
    .A2(net8226));
 sg13g2_nand2_1 _23318_ (.Y(_14173_),
    .A(net3109),
    .B(net8228));
 sg13g2_o21ai_1 _23319_ (.B1(_14173_),
    .Y(_00376_),
    .A1(net7595),
    .A2(net8228));
 sg13g2_nand2_1 _23320_ (.Y(_14174_),
    .A(net4111),
    .B(net8221));
 sg13g2_o21ai_1 _23321_ (.B1(_14174_),
    .Y(_00377_),
    .A1(net7603),
    .A2(net8221));
 sg13g2_nand2_1 _23322_ (.Y(_14175_),
    .A(net3264),
    .B(net8227));
 sg13g2_o21ai_1 _23323_ (.B1(_14175_),
    .Y(_00378_),
    .A1(net7557),
    .A2(net8227));
 sg13g2_nand2_1 _23324_ (.Y(_14176_),
    .A(net3163),
    .B(net8230));
 sg13g2_o21ai_1 _23325_ (.B1(_14176_),
    .Y(_00379_),
    .A1(net7575),
    .A2(net8230));
 sg13g2_nand2_1 _23326_ (.Y(_14177_),
    .A(net3005),
    .B(net8228));
 sg13g2_o21ai_1 _23327_ (.B1(_14177_),
    .Y(_00380_),
    .A1(net7548),
    .A2(net8228));
 sg13g2_nand2_1 _23328_ (.Y(_14178_),
    .A(net3462),
    .B(net8221));
 sg13g2_o21ai_1 _23329_ (.B1(_14178_),
    .Y(_00381_),
    .A1(net7570),
    .A2(net8221));
 sg13g2_nand2_1 _23330_ (.Y(_14179_),
    .A(net2939),
    .B(net8228));
 sg13g2_o21ai_1 _23331_ (.B1(_14179_),
    .Y(_00382_),
    .A1(net7544),
    .A2(net8228));
 sg13g2_nand2_1 _23332_ (.Y(_14180_),
    .A(net3208),
    .B(net8230));
 sg13g2_o21ai_1 _23333_ (.B1(_14180_),
    .Y(_00383_),
    .A1(net7553),
    .A2(net8230));
 sg13g2_nand2_1 _23334_ (.Y(_14181_),
    .A(net3435),
    .B(net8224));
 sg13g2_o21ai_1 _23335_ (.B1(_14181_),
    .Y(_00384_),
    .A1(net7583),
    .A2(net8224));
 sg13g2_nand2_1 _23336_ (.Y(_14182_),
    .A(net3319),
    .B(net8222));
 sg13g2_o21ai_1 _23337_ (.B1(_14182_),
    .Y(_00385_),
    .A1(net7564),
    .A2(net8222));
 sg13g2_nand2_1 _23338_ (.Y(_14183_),
    .A(net2989),
    .B(net8221));
 sg13g2_o21ai_1 _23339_ (.B1(_14183_),
    .Y(_00386_),
    .A1(net7523),
    .A2(net8221));
 sg13g2_nand2_1 _23340_ (.Y(_14184_),
    .A(net3015),
    .B(net8221));
 sg13g2_o21ai_1 _23341_ (.B1(_14184_),
    .Y(_00387_),
    .A1(net7536),
    .A2(net8221));
 sg13g2_nand2_1 _23342_ (.Y(_14185_),
    .A(net2796),
    .B(net8223));
 sg13g2_o21ai_1 _23343_ (.B1(_14185_),
    .Y(_00388_),
    .A1(net7529),
    .A2(net8223));
 sg13g2_nand2_1 _23344_ (.Y(_14186_),
    .A(net2766),
    .B(net8224));
 sg13g2_o21ai_1 _23345_ (.B1(_14186_),
    .Y(_00389_),
    .A1(net7520),
    .A2(net8224));
 sg13g2_nand2_1 _23346_ (.Y(_14187_),
    .A(net2627),
    .B(net8231));
 sg13g2_o21ai_1 _23347_ (.B1(_14187_),
    .Y(_00390_),
    .A1(net7507),
    .A2(net8231));
 sg13g2_nand2_1 _23348_ (.Y(_14188_),
    .A(net3118),
    .B(net8226));
 sg13g2_o21ai_1 _23349_ (.B1(_14188_),
    .Y(_00391_),
    .A1(net7514),
    .A2(net8226));
 sg13g2_nand2_1 _23350_ (.Y(_14189_),
    .A(net3082),
    .B(net8229));
 sg13g2_o21ai_1 _23351_ (.B1(_14189_),
    .Y(_00392_),
    .A1(net7495),
    .A2(net8229));
 sg13g2_nand2_1 _23352_ (.Y(_14190_),
    .A(net3684),
    .B(net8222));
 sg13g2_o21ai_1 _23353_ (.B1(_14190_),
    .Y(_00393_),
    .A1(net7499),
    .A2(net8222));
 sg13g2_nand2_1 _23354_ (.Y(_14191_),
    .A(net3341),
    .B(net8226));
 sg13g2_o21ai_1 _23355_ (.B1(_14191_),
    .Y(_00394_),
    .A1(net7645),
    .A2(net8226));
 sg13g2_nand2_1 _23356_ (.Y(_14192_),
    .A(net3575),
    .B(net8227));
 sg13g2_o21ai_1 _23357_ (.B1(_14192_),
    .Y(_00395_),
    .A1(net7648),
    .A2(net8227));
 sg13g2_nand2_1 _23358_ (.Y(_14193_),
    .A(net2938),
    .B(net8228));
 sg13g2_o21ai_1 _23359_ (.B1(_14193_),
    .Y(_00396_),
    .A1(net7654),
    .A2(net8228));
 sg13g2_nand2_1 _23360_ (.Y(_14194_),
    .A(net3447),
    .B(net8224));
 sg13g2_o21ai_1 _23361_ (.B1(_14194_),
    .Y(_00397_),
    .A1(net7658),
    .A2(net8224));
 sg13g2_nand2_1 _23362_ (.Y(_14195_),
    .A(net2792),
    .B(net8224));
 sg13g2_o21ai_1 _23363_ (.B1(_14195_),
    .Y(_00398_),
    .A1(net7639),
    .A2(net8224));
 sg13g2_nand2_1 _23364_ (.Y(_14196_),
    .A(net3499),
    .B(net8227));
 sg13g2_o21ai_1 _23365_ (.B1(_14196_),
    .Y(_00399_),
    .A1(net7628),
    .A2(net8227));
 sg13g2_nand2_1 _23366_ (.Y(_14197_),
    .A(net3088),
    .B(net8225));
 sg13g2_o21ai_1 _23367_ (.B1(_14197_),
    .Y(_00400_),
    .A1(net7623),
    .A2(net8225));
 sg13g2_nand2_1 _23368_ (.Y(_14198_),
    .A(net2817),
    .B(net8225));
 sg13g2_o21ai_1 _23369_ (.B1(_14198_),
    .Y(_00401_),
    .A1(net7630),
    .A2(net8225));
 sg13g2_nor2_2 _23370_ (.A(_10467_),
    .B(_10468_),
    .Y(_14199_));
 sg13g2_nand3_1 _23371_ (.B(_14165_),
    .C(_14199_),
    .A(net8371),
    .Y(_14200_));
 sg13g2_nand2_1 _23372_ (.Y(_14201_),
    .A(net3369),
    .B(net8219));
 sg13g2_o21ai_1 _23373_ (.B1(_14201_),
    .Y(_00402_),
    .A1(net7489),
    .A2(net8219));
 sg13g2_nand2_1 _23374_ (.Y(_14202_),
    .A(net3138),
    .B(net8219));
 sg13g2_o21ai_1 _23375_ (.B1(_14202_),
    .Y(_00403_),
    .A1(net7663),
    .A2(net8219));
 sg13g2_nand2_1 _23376_ (.Y(_14203_),
    .A(net3299),
    .B(net8219));
 sg13g2_o21ai_1 _23377_ (.B1(_14203_),
    .Y(_00404_),
    .A1(net7612),
    .A2(net8219));
 sg13g2_nand2_1 _23378_ (.Y(_14204_),
    .A(net3350),
    .B(net8217));
 sg13g2_o21ai_1 _23379_ (.B1(_14204_),
    .Y(_00405_),
    .A1(net7610),
    .A2(net8217));
 sg13g2_nand2_1 _23380_ (.Y(_14205_),
    .A(net3554),
    .B(net8214));
 sg13g2_o21ai_1 _23381_ (.B1(_14205_),
    .Y(_00406_),
    .A1(net7588),
    .A2(net8214));
 sg13g2_nand2_1 _23382_ (.Y(_14206_),
    .A(net3134),
    .B(net8214));
 sg13g2_o21ai_1 _23383_ (.B1(_14206_),
    .Y(_00407_),
    .A1(net7597),
    .A2(net8214));
 sg13g2_nand2_1 _23384_ (.Y(_14207_),
    .A(net3808),
    .B(net8216));
 sg13g2_o21ai_1 _23385_ (.B1(_14207_),
    .Y(_00408_),
    .A1(net7595),
    .A2(net8216));
 sg13g2_nand2_1 _23386_ (.Y(_14208_),
    .A(net3490),
    .B(net8209));
 sg13g2_o21ai_1 _23387_ (.B1(_14208_),
    .Y(_00409_),
    .A1(net7603),
    .A2(net8209));
 sg13g2_nand2_1 _23388_ (.Y(_14209_),
    .A(net3504),
    .B(net8215));
 sg13g2_o21ai_1 _23389_ (.B1(_14209_),
    .Y(_00410_),
    .A1(net7557),
    .A2(net8215));
 sg13g2_nand2_1 _23390_ (.Y(_14210_),
    .A(net3308),
    .B(net8218));
 sg13g2_o21ai_1 _23391_ (.B1(_14210_),
    .Y(_00411_),
    .A1(net7575),
    .A2(net8218));
 sg13g2_nand2_1 _23392_ (.Y(_14211_),
    .A(net3285),
    .B(net8216));
 sg13g2_o21ai_1 _23393_ (.B1(_14211_),
    .Y(_00412_),
    .A1(net7548),
    .A2(net8216));
 sg13g2_nand2_1 _23394_ (.Y(_14212_),
    .A(net3503),
    .B(net8209));
 sg13g2_o21ai_1 _23395_ (.B1(_14212_),
    .Y(_00413_),
    .A1(net7569),
    .A2(net8209));
 sg13g2_nand2_1 _23396_ (.Y(_14213_),
    .A(net3839),
    .B(net8216));
 sg13g2_o21ai_1 _23397_ (.B1(_14213_),
    .Y(_00414_),
    .A1(net7543),
    .A2(net8216));
 sg13g2_nand2_1 _23398_ (.Y(_14214_),
    .A(net3153),
    .B(net8218));
 sg13g2_o21ai_1 _23399_ (.B1(_14214_),
    .Y(_00415_),
    .A1(net7553),
    .A2(net8218));
 sg13g2_nand2_1 _23400_ (.Y(_14215_),
    .A(net3320),
    .B(net8212));
 sg13g2_o21ai_1 _23401_ (.B1(_14215_),
    .Y(_00416_),
    .A1(net7583),
    .A2(net8212));
 sg13g2_nand2_1 _23402_ (.Y(_14216_),
    .A(net3012),
    .B(net8211));
 sg13g2_o21ai_1 _23403_ (.B1(_14216_),
    .Y(_00417_),
    .A1(net7564),
    .A2(net8211));
 sg13g2_nand2_1 _23404_ (.Y(_14217_),
    .A(net3611),
    .B(net8209));
 sg13g2_o21ai_1 _23405_ (.B1(_14217_),
    .Y(_00418_),
    .A1(net7523),
    .A2(net8209));
 sg13g2_nand2_1 _23406_ (.Y(_14218_),
    .A(net3517),
    .B(net8209));
 sg13g2_o21ai_1 _23407_ (.B1(_14218_),
    .Y(_00419_),
    .A1(net7536),
    .A2(net8209));
 sg13g2_nand2_1 _23408_ (.Y(_14219_),
    .A(net4051),
    .B(net8210));
 sg13g2_o21ai_1 _23409_ (.B1(_14219_),
    .Y(_00420_),
    .A1(net7529),
    .A2(net8210));
 sg13g2_nand2_1 _23410_ (.Y(_14220_),
    .A(net3465),
    .B(net8212));
 sg13g2_o21ai_1 _23411_ (.B1(_14220_),
    .Y(_00421_),
    .A1(net7520),
    .A2(net8212));
 sg13g2_nand2_1 _23412_ (.Y(_14221_),
    .A(net3645),
    .B(net8219));
 sg13g2_o21ai_1 _23413_ (.B1(_14221_),
    .Y(_00422_),
    .A1(net7507),
    .A2(net8219));
 sg13g2_nand2_1 _23414_ (.Y(_14222_),
    .A(net3592),
    .B(net8214));
 sg13g2_o21ai_1 _23415_ (.B1(_14222_),
    .Y(_00423_),
    .A1(net7513),
    .A2(net8214));
 sg13g2_nand2_1 _23416_ (.Y(_14223_),
    .A(net3228),
    .B(net8217));
 sg13g2_o21ai_1 _23417_ (.B1(_14223_),
    .Y(_00424_),
    .A1(net7495),
    .A2(net8217));
 sg13g2_nand2_1 _23418_ (.Y(_14224_),
    .A(net3596),
    .B(net8210));
 sg13g2_o21ai_1 _23419_ (.B1(_14224_),
    .Y(_00425_),
    .A1(net7499),
    .A2(net8210));
 sg13g2_nand2_1 _23420_ (.Y(_14225_),
    .A(net3992),
    .B(net8214));
 sg13g2_o21ai_1 _23421_ (.B1(_14225_),
    .Y(_00426_),
    .A1(net7644),
    .A2(net8214));
 sg13g2_nand2_1 _23422_ (.Y(_14226_),
    .A(net3463),
    .B(net8215));
 sg13g2_o21ai_1 _23423_ (.B1(_14226_),
    .Y(_00427_),
    .A1(net7648),
    .A2(net8215));
 sg13g2_nand2_1 _23424_ (.Y(_14227_),
    .A(net3591),
    .B(net8216));
 sg13g2_o21ai_1 _23425_ (.B1(_14227_),
    .Y(_00428_),
    .A1(net7655),
    .A2(net8216));
 sg13g2_nand2_1 _23426_ (.Y(_14228_),
    .A(net3960),
    .B(net8212));
 sg13g2_o21ai_1 _23427_ (.B1(_14228_),
    .Y(_00429_),
    .A1(net7658),
    .A2(net8212));
 sg13g2_nand2_1 _23428_ (.Y(_14229_),
    .A(net3656),
    .B(net8212));
 sg13g2_o21ai_1 _23429_ (.B1(_14229_),
    .Y(_00430_),
    .A1(net7638),
    .A2(net8212));
 sg13g2_nand2_1 _23430_ (.Y(_14230_),
    .A(net3359),
    .B(net8215));
 sg13g2_o21ai_1 _23431_ (.B1(_14230_),
    .Y(_00431_),
    .A1(net7628),
    .A2(net8215));
 sg13g2_nand2_1 _23432_ (.Y(_14231_),
    .A(net3466),
    .B(net8213));
 sg13g2_o21ai_1 _23433_ (.B1(_14231_),
    .Y(_00432_),
    .A1(net7622),
    .A2(net8213));
 sg13g2_nand2_1 _23434_ (.Y(_14232_),
    .A(net3662),
    .B(net8211));
 sg13g2_o21ai_1 _23435_ (.B1(_14232_),
    .Y(_00433_),
    .A1(net7633),
    .A2(net8211));
 sg13g2_nand4_1 _23436_ (.B(net8961),
    .C(_14127_),
    .A(net9710),
    .Y(_14233_),
    .D(net8371));
 sg13g2_nand2_1 _23437_ (.Y(_14234_),
    .A(net3473),
    .B(net8203));
 sg13g2_o21ai_1 _23438_ (.B1(_14234_),
    .Y(_00434_),
    .A1(net7488),
    .A2(net8203));
 sg13g2_nand2_1 _23439_ (.Y(_14235_),
    .A(net2968),
    .B(net8207));
 sg13g2_o21ai_1 _23440_ (.B1(_14235_),
    .Y(_00435_),
    .A1(net7664),
    .A2(net8207));
 sg13g2_nand2_1 _23441_ (.Y(_14236_),
    .A(net3006),
    .B(net8203));
 sg13g2_o21ai_1 _23442_ (.B1(_14236_),
    .Y(_00436_),
    .A1(net7614),
    .A2(net8203));
 sg13g2_nand2_1 _23443_ (.Y(_14237_),
    .A(net3185),
    .B(net8205));
 sg13g2_o21ai_1 _23444_ (.B1(_14237_),
    .Y(_00437_),
    .A1(net7610),
    .A2(net8205));
 sg13g2_nand2_1 _23445_ (.Y(_14238_),
    .A(net4005),
    .B(net8203));
 sg13g2_o21ai_1 _23446_ (.B1(_14238_),
    .Y(_00438_),
    .A1(net7589),
    .A2(net8203));
 sg13g2_nand2_1 _23447_ (.Y(_14239_),
    .A(net3703),
    .B(net8201));
 sg13g2_o21ai_1 _23448_ (.B1(_14239_),
    .Y(_00439_),
    .A1(net7597),
    .A2(net8201));
 sg13g2_nand2_1 _23449_ (.Y(_14240_),
    .A(net3068),
    .B(net8204));
 sg13g2_o21ai_1 _23450_ (.B1(_14240_),
    .Y(_00440_),
    .A1(net7595),
    .A2(net8204));
 sg13g2_nand2_1 _23451_ (.Y(_14241_),
    .A(net2928),
    .B(net8197));
 sg13g2_o21ai_1 _23452_ (.B1(_14241_),
    .Y(_00441_),
    .A1(net7602),
    .A2(net8197));
 sg13g2_nand2_1 _23453_ (.Y(_14242_),
    .A(net3043),
    .B(net8202));
 sg13g2_o21ai_1 _23454_ (.B1(_14242_),
    .Y(_00442_),
    .A1(net7560),
    .A2(net8202));
 sg13g2_nand2_1 _23455_ (.Y(_14243_),
    .A(net3049),
    .B(net8206));
 sg13g2_o21ai_1 _23456_ (.B1(_14243_),
    .Y(_00443_),
    .A1(net7575),
    .A2(net8206));
 sg13g2_nand2_1 _23457_ (.Y(_14244_),
    .A(net3167),
    .B(net8205));
 sg13g2_o21ai_1 _23458_ (.B1(_14244_),
    .Y(_00444_),
    .A1(net7548),
    .A2(net8205));
 sg13g2_nand2_1 _23459_ (.Y(_14245_),
    .A(net3262),
    .B(net8197));
 sg13g2_o21ai_1 _23460_ (.B1(_14245_),
    .Y(_00445_),
    .A1(net7569),
    .A2(net8197));
 sg13g2_nand2_1 _23461_ (.Y(_14246_),
    .A(net2879),
    .B(net8204));
 sg13g2_o21ai_1 _23462_ (.B1(_14246_),
    .Y(_00446_),
    .A1(net7543),
    .A2(net8204));
 sg13g2_nand2_1 _23463_ (.Y(_14247_),
    .A(net3371),
    .B(net8206));
 sg13g2_o21ai_1 _23464_ (.B1(_14247_),
    .Y(_00447_),
    .A1(net7553),
    .A2(net8206));
 sg13g2_nand2_1 _23465_ (.Y(_14248_),
    .A(net3456),
    .B(net8199));
 sg13g2_o21ai_1 _23466_ (.B1(_14248_),
    .Y(_00448_),
    .A1(net7585),
    .A2(net8199));
 sg13g2_nand2_1 _23467_ (.Y(_14249_),
    .A(net3270),
    .B(net8198));
 sg13g2_o21ai_1 _23468_ (.B1(_14249_),
    .Y(_00449_),
    .A1(net7563),
    .A2(net8198));
 sg13g2_nand2_1 _23469_ (.Y(_14250_),
    .A(net4073),
    .B(net8197));
 sg13g2_o21ai_1 _23470_ (.B1(_14250_),
    .Y(_00450_),
    .A1(net7524),
    .A2(net8197));
 sg13g2_nand2_1 _23471_ (.Y(_14251_),
    .A(net2951),
    .B(net8197));
 sg13g2_o21ai_1 _23472_ (.B1(_14251_),
    .Y(_00451_),
    .A1(net7536),
    .A2(net8197));
 sg13g2_nand2_1 _23473_ (.Y(_14252_),
    .A(net3430),
    .B(net8198));
 sg13g2_o21ai_1 _23474_ (.B1(_14252_),
    .Y(_00452_),
    .A1(net7528),
    .A2(net8198));
 sg13g2_nand2_1 _23475_ (.Y(_14253_),
    .A(net3124),
    .B(net8199));
 sg13g2_o21ai_1 _23476_ (.B1(_14253_),
    .Y(_00453_),
    .A1(net7520),
    .A2(net8199));
 sg13g2_nand2_1 _23477_ (.Y(_14254_),
    .A(net3363),
    .B(net8203));
 sg13g2_o21ai_1 _23478_ (.B1(_14254_),
    .Y(_00454_),
    .A1(net7506),
    .A2(net8203));
 sg13g2_nand2_1 _23479_ (.Y(_14255_),
    .A(net2908),
    .B(net8201));
 sg13g2_o21ai_1 _23480_ (.B1(_14255_),
    .Y(_00455_),
    .A1(net7514),
    .A2(net8201));
 sg13g2_nand2_1 _23481_ (.Y(_14256_),
    .A(net3556),
    .B(net8204));
 sg13g2_o21ai_1 _23482_ (.B1(_14256_),
    .Y(_00456_),
    .A1(net7495),
    .A2(net8204));
 sg13g2_nand2_1 _23483_ (.Y(_14257_),
    .A(net3372),
    .B(net8198));
 sg13g2_o21ai_1 _23484_ (.B1(_14257_),
    .Y(_00457_),
    .A1(net7501),
    .A2(net8198));
 sg13g2_nand2_1 _23485_ (.Y(_14258_),
    .A(net3995),
    .B(net8201));
 sg13g2_o21ai_1 _23486_ (.B1(_14258_),
    .Y(_00458_),
    .A1(net7644),
    .A2(net8201));
 sg13g2_nand2_1 _23487_ (.Y(_14259_),
    .A(net3560),
    .B(net8201));
 sg13g2_o21ai_1 _23488_ (.B1(_14259_),
    .Y(_00459_),
    .A1(net7649),
    .A2(net8201));
 sg13g2_nand2_1 _23489_ (.Y(_14260_),
    .A(net3261),
    .B(net8204));
 sg13g2_o21ai_1 _23490_ (.B1(_14260_),
    .Y(_00460_),
    .A1(net7654),
    .A2(net8204));
 sg13g2_nand2_1 _23491_ (.Y(_14261_),
    .A(net3322),
    .B(net8200));
 sg13g2_o21ai_1 _23492_ (.B1(_14261_),
    .Y(_00461_),
    .A1(net7660),
    .A2(net8200));
 sg13g2_nand2_1 _23493_ (.Y(_14262_),
    .A(net3179),
    .B(net8199));
 sg13g2_o21ai_1 _23494_ (.B1(_14262_),
    .Y(_00462_),
    .A1(net7641),
    .A2(net8199));
 sg13g2_nand2_1 _23495_ (.Y(_14263_),
    .A(net3231),
    .B(net8202));
 sg13g2_o21ai_1 _23496_ (.B1(_14263_),
    .Y(_00463_),
    .A1(net7627),
    .A2(net8202));
 sg13g2_nand2_1 _23497_ (.Y(_14264_),
    .A(net3126),
    .B(net8199));
 sg13g2_o21ai_1 _23498_ (.B1(_14264_),
    .Y(_00464_),
    .A1(net7619),
    .A2(net8199));
 sg13g2_nand2_1 _23499_ (.Y(_14265_),
    .A(net3216),
    .B(net8200));
 sg13g2_o21ai_1 _23500_ (.B1(_14265_),
    .Y(_00465_),
    .A1(net7633),
    .A2(net8200));
 sg13g2_o21ai_1 _23501_ (.B1(_10571_),
    .Y(_14266_),
    .A1(net9265),
    .A2(_11847_));
 sg13g2_nor3_1 _23502_ (.A(net9265),
    .B(\soc_I.qqspi_I.xfer_cycles[1] ),
    .C(\soc_I.qqspi_I.xfer_cycles[0] ),
    .Y(_14267_));
 sg13g2_o21ai_1 _23503_ (.B1(_14266_),
    .Y(_14268_),
    .A1(_10571_),
    .A2(_14267_));
 sg13g2_a21oi_1 _23504_ (.A1(net9265),
    .A2(_10694_),
    .Y(_14269_),
    .B1(net8683));
 sg13g2_nor3_1 _23505_ (.A(_00243_),
    .B(net8681),
    .C(_12557_),
    .Y(_14270_));
 sg13g2_nor2_1 _23506_ (.A(_10377_),
    .B(net8684),
    .Y(_14271_));
 sg13g2_nor2_1 _23507_ (.A(\soc_I.qqspi_I.state[1] ),
    .B(\soc_I.qqspi_I.state[0] ),
    .Y(_14272_));
 sg13g2_nor2_1 _23508_ (.A(\soc_I.qqspi_I.state[5] ),
    .B(net8682),
    .Y(_14273_));
 sg13g2_inv_1 _23509_ (.Y(_14274_),
    .A(net8603));
 sg13g2_nand3b_1 _23510_ (.B(_00242_),
    .C(_14273_),
    .Y(_14275_),
    .A_N(\soc_I.qqspi_I.state[2] ));
 sg13g2_nor3_1 _23511_ (.A(\soc_I.qqspi_I.state[1] ),
    .B(\soc_I.qqspi_I.state[0] ),
    .C(_14275_),
    .Y(_14276_));
 sg13g2_nor3_2 _23512_ (.A(_14270_),
    .B(_14271_),
    .C(_14276_),
    .Y(_14277_));
 sg13g2_nand2_1 _23513_ (.Y(_14278_),
    .A(\soc_I.qqspi_I.state[1] ),
    .B(net8684));
 sg13g2_a22oi_1 _23514_ (.Y(_14279_),
    .B1(_14268_),
    .B2(_14269_),
    .A2(net8683),
    .A1(\soc_I.qqspi_I.state[1] ));
 sg13g2_o21ai_1 _23515_ (.B1(net9344),
    .Y(_14280_),
    .A1(net4856),
    .A2(net7389));
 sg13g2_a21oi_1 _23516_ (.A1(net7389),
    .A2(_14279_),
    .Y(_00466_),
    .B1(_14280_));
 sg13g2_nor2_1 _23517_ (.A(\soc_I.qqspi_I.xfer_cycles[3] ),
    .B(_14266_),
    .Y(_14281_));
 sg13g2_xnor2_1 _23518_ (.Y(_14282_),
    .A(net5182),
    .B(_14266_));
 sg13g2_nor2_1 _23519_ (.A(\soc_I.qqspi_I.state[2] ),
    .B(\soc_I.qqspi_I.state[6] ),
    .Y(_14283_));
 sg13g2_nor2_1 _23520_ (.A(\soc_I.qqspi_I.state[1] ),
    .B(net9195),
    .Y(_14284_));
 sg13g2_a21oi_2 _23521_ (.B1(net8681),
    .Y(_14285_),
    .A2(_14284_),
    .A1(_14283_));
 sg13g2_nand3_1 _23522_ (.B(net8665),
    .C(net8958),
    .A(net9195),
    .Y(_14286_));
 sg13g2_nand2_1 _23523_ (.Y(_14287_),
    .A(_14283_),
    .B(_14286_));
 sg13g2_a22oi_1 _23524_ (.Y(_14288_),
    .B1(_14285_),
    .B2(_14287_),
    .A2(_14282_),
    .A1(net8681));
 sg13g2_o21ai_1 _23525_ (.B1(net9343),
    .Y(_14289_),
    .A1(net5182),
    .A2(net7389));
 sg13g2_a21oi_1 _23526_ (.A1(net7389),
    .A2(_14288_),
    .Y(_00467_),
    .B1(_14289_));
 sg13g2_nand3_1 _23527_ (.B(net8666),
    .C(net8962),
    .A(net9195),
    .Y(_14290_));
 sg13g2_nand2_1 _23528_ (.Y(_14291_),
    .A(_00242_),
    .B(_14290_));
 sg13g2_xor2_1 _23529_ (.B(_14281_),
    .A(net5050),
    .X(_14292_));
 sg13g2_a22oi_1 _23530_ (.Y(_14293_),
    .B1(_14292_),
    .B2(net8681),
    .A2(_14291_),
    .A1(_14285_));
 sg13g2_o21ai_1 _23531_ (.B1(net9343),
    .Y(_14294_),
    .A1(net5050),
    .A2(_14277_));
 sg13g2_a21oi_1 _23532_ (.A1(net7389),
    .A2(_14293_),
    .Y(_00468_),
    .B1(_14294_));
 sg13g2_nand2_1 _23533_ (.Y(_14295_),
    .A(net9265),
    .B(_11848_));
 sg13g2_xnor2_1 _23534_ (.Y(_14296_),
    .A(net5104),
    .B(_14295_));
 sg13g2_nand2b_2 _23535_ (.Y(_14297_),
    .B(net8666),
    .A_N(net9700));
 sg13g2_nor2b_1 _23536_ (.A(_00291_),
    .B_N(_14285_),
    .Y(_14298_));
 sg13g2_a22oi_1 _23537_ (.Y(_14299_),
    .B1(_14297_),
    .B2(_14298_),
    .A2(_14296_),
    .A1(_11849_));
 sg13g2_o21ai_1 _23538_ (.B1(net9343),
    .Y(_14300_),
    .A1(net5104),
    .A2(net7389));
 sg13g2_a21oi_1 _23539_ (.A1(net7389),
    .A2(_14299_),
    .Y(_00469_),
    .B1(_14300_));
 sg13g2_nor2_2 _23540_ (.A(\soc_I.kianv_I.Instr[8] ),
    .B(_10468_),
    .Y(_14301_));
 sg13g2_nor2b_2 _23541_ (.A(_14128_),
    .B_N(_14301_),
    .Y(_14302_));
 sg13g2_and3_1 _23542_ (.X(_14303_),
    .A(net9710),
    .B(_14127_),
    .C(_14302_));
 sg13g2_nor2_1 _23543_ (.A(net3991),
    .B(net8191),
    .Y(_14304_));
 sg13g2_a21oi_1 _23544_ (.A1(net7488),
    .A2(net8191),
    .Y(_00470_),
    .B1(_14304_));
 sg13g2_nor2_1 _23545_ (.A(net3634),
    .B(net8195),
    .Y(_14305_));
 sg13g2_a21oi_1 _23546_ (.A1(net7664),
    .A2(net8195),
    .Y(_00471_),
    .B1(_14305_));
 sg13g2_nor2_1 _23547_ (.A(net3980),
    .B(net8191),
    .Y(_14306_));
 sg13g2_a21oi_1 _23548_ (.A1(net7614),
    .A2(net8191),
    .Y(_00472_),
    .B1(_14306_));
 sg13g2_nor2_1 _23549_ (.A(net3523),
    .B(net8193),
    .Y(_14307_));
 sg13g2_a21oi_1 _23550_ (.A1(net7610),
    .A2(net8193),
    .Y(_00473_),
    .B1(_14307_));
 sg13g2_nor2_1 _23551_ (.A(net4066),
    .B(net8191),
    .Y(_14308_));
 sg13g2_a21oi_1 _23552_ (.A1(net7589),
    .A2(net8191),
    .Y(_00474_),
    .B1(_14308_));
 sg13g2_nor2_1 _23553_ (.A(net4018),
    .B(net8189),
    .Y(_14309_));
 sg13g2_a21oi_1 _23554_ (.A1(net7601),
    .A2(net8189),
    .Y(_00475_),
    .B1(_14309_));
 sg13g2_nor2_1 _23555_ (.A(net3599),
    .B(net8192),
    .Y(_14310_));
 sg13g2_a21oi_1 _23556_ (.A1(net7594),
    .A2(net8192),
    .Y(_00476_),
    .B1(_14310_));
 sg13g2_nor2_1 _23557_ (.A(net4587),
    .B(net8185),
    .Y(_14311_));
 sg13g2_a21oi_1 _23558_ (.A1(_12918_),
    .A2(net8185),
    .Y(_00477_),
    .B1(_14311_));
 sg13g2_nor2_1 _23559_ (.A(net4206),
    .B(net8190),
    .Y(_14312_));
 sg13g2_a21oi_1 _23560_ (.A1(net7560),
    .A2(net8190),
    .Y(_00478_),
    .B1(_14312_));
 sg13g2_nor2_1 _23561_ (.A(net3804),
    .B(net8194),
    .Y(_14313_));
 sg13g2_a21oi_1 _23562_ (.A1(net7575),
    .A2(net8194),
    .Y(_00479_),
    .B1(_14313_));
 sg13g2_nor2_1 _23563_ (.A(net3900),
    .B(net8193),
    .Y(_14314_));
 sg13g2_a21oi_1 _23564_ (.A1(net7548),
    .A2(net8193),
    .Y(_00480_),
    .B1(_14314_));
 sg13g2_nor2_1 _23565_ (.A(net3521),
    .B(net8184),
    .Y(_14315_));
 sg13g2_a21oi_1 _23566_ (.A1(net7569),
    .A2(net8184),
    .Y(_00481_),
    .B1(_14315_));
 sg13g2_nor2_1 _23567_ (.A(net3603),
    .B(net8192),
    .Y(_14316_));
 sg13g2_a21oi_1 _23568_ (.A1(net7543),
    .A2(net8192),
    .Y(_00482_),
    .B1(_14316_));
 sg13g2_nor2_1 _23569_ (.A(net3914),
    .B(net8194),
    .Y(_14317_));
 sg13g2_a21oi_1 _23570_ (.A1(net7555),
    .A2(net8194),
    .Y(_00483_),
    .B1(_14317_));
 sg13g2_nor2_1 _23571_ (.A(net3730),
    .B(net8187),
    .Y(_14318_));
 sg13g2_a21oi_1 _23572_ (.A1(net7584),
    .A2(net8187),
    .Y(_00484_),
    .B1(_14318_));
 sg13g2_nor2_1 _23573_ (.A(net3889),
    .B(net8185),
    .Y(_14319_));
 sg13g2_a21oi_1 _23574_ (.A1(net7563),
    .A2(net8185),
    .Y(_00485_),
    .B1(_14319_));
 sg13g2_nor2_1 _23575_ (.A(net3331),
    .B(net8184),
    .Y(_14320_));
 sg13g2_a21oi_1 _23576_ (.A1(net7523),
    .A2(net8184),
    .Y(_00486_),
    .B1(_14320_));
 sg13g2_nor2_1 _23577_ (.A(net3834),
    .B(net8184),
    .Y(_14321_));
 sg13g2_a21oi_1 _23578_ (.A1(net7536),
    .A2(net8184),
    .Y(_00487_),
    .B1(_14321_));
 sg13g2_nor2_1 _23579_ (.A(net3840),
    .B(net8184),
    .Y(_14322_));
 sg13g2_a21oi_1 _23580_ (.A1(net7528),
    .A2(net8184),
    .Y(_00488_),
    .B1(_14322_));
 sg13g2_nor2_1 _23581_ (.A(net3571),
    .B(net8187),
    .Y(_14323_));
 sg13g2_a21oi_1 _23582_ (.A1(net7520),
    .A2(net8187),
    .Y(_00489_),
    .B1(_14323_));
 sg13g2_nor2_1 _23583_ (.A(net3569),
    .B(net8191),
    .Y(_14324_));
 sg13g2_a21oi_1 _23584_ (.A1(net7506),
    .A2(net8191),
    .Y(_00490_),
    .B1(_14324_));
 sg13g2_nor2_1 _23585_ (.A(net4122),
    .B(net8189),
    .Y(_14325_));
 sg13g2_a21oi_1 _23586_ (.A1(net7514),
    .A2(net8189),
    .Y(_00491_),
    .B1(_14325_));
 sg13g2_nor2_1 _23587_ (.A(net3740),
    .B(net8192),
    .Y(_14326_));
 sg13g2_a21oi_1 _23588_ (.A1(net7495),
    .A2(net8192),
    .Y(_00492_),
    .B1(_14326_));
 sg13g2_nor2_1 _23589_ (.A(net3623),
    .B(net8185),
    .Y(_14327_));
 sg13g2_a21oi_1 _23590_ (.A1(net7501),
    .A2(net8185),
    .Y(_00493_),
    .B1(_14327_));
 sg13g2_nor2_1 _23591_ (.A(net3782),
    .B(net8189),
    .Y(_14328_));
 sg13g2_a21oi_1 _23592_ (.A1(net7643),
    .A2(net8189),
    .Y(_00494_),
    .B1(_14328_));
 sg13g2_nor2_1 _23593_ (.A(net3932),
    .B(net8189),
    .Y(_14329_));
 sg13g2_a21oi_1 _23594_ (.A1(net7648),
    .A2(net8189),
    .Y(_00495_),
    .B1(_14329_));
 sg13g2_nor2_1 _23595_ (.A(net3568),
    .B(net8192),
    .Y(_14330_));
 sg13g2_a21oi_1 _23596_ (.A1(net7654),
    .A2(net8192),
    .Y(_00496_),
    .B1(_14330_));
 sg13g2_nor2_1 _23597_ (.A(net3990),
    .B(net8188),
    .Y(_14331_));
 sg13g2_a21oi_1 _23598_ (.A1(net7661),
    .A2(net8188),
    .Y(_00497_),
    .B1(_14331_));
 sg13g2_nor2_1 _23599_ (.A(net3529),
    .B(net8187),
    .Y(_14332_));
 sg13g2_a21oi_1 _23600_ (.A1(net7640),
    .A2(net8187),
    .Y(_00498_),
    .B1(_14332_));
 sg13g2_nor2_1 _23601_ (.A(net3677),
    .B(net8190),
    .Y(_14333_));
 sg13g2_a21oi_1 _23602_ (.A1(net7627),
    .A2(net8190),
    .Y(_00499_),
    .B1(_14333_));
 sg13g2_nor2_1 _23603_ (.A(net3917),
    .B(net8187),
    .Y(_14334_));
 sg13g2_a21oi_1 _23604_ (.A1(net7621),
    .A2(net8187),
    .Y(_00500_),
    .B1(_14334_));
 sg13g2_nor2_1 _23605_ (.A(net3843),
    .B(net8186),
    .Y(_14335_));
 sg13g2_a21oi_1 _23606_ (.A1(net7633),
    .A2(net8186),
    .Y(_00501_),
    .B1(_14335_));
 sg13g2_nand4_1 _23607_ (.B(_14126_),
    .C(_14127_),
    .A(net9710),
    .Y(_14336_),
    .D(net8371));
 sg13g2_nand2_1 _23608_ (.Y(_14337_),
    .A(net3045),
    .B(net8178));
 sg13g2_o21ai_1 _23609_ (.B1(_14337_),
    .Y(_00502_),
    .A1(net7488),
    .A2(net8178));
 sg13g2_nand2_1 _23610_ (.Y(_14338_),
    .A(net2686),
    .B(net8182));
 sg13g2_o21ai_1 _23611_ (.B1(_14338_),
    .Y(_00503_),
    .A1(net7664),
    .A2(net8182));
 sg13g2_nand2_1 _23612_ (.Y(_14339_),
    .A(net3022),
    .B(net8178));
 sg13g2_o21ai_1 _23613_ (.B1(_14339_),
    .Y(_00504_),
    .A1(net7612),
    .A2(net8178));
 sg13g2_nand2_1 _23614_ (.Y(_14340_),
    .A(net3271),
    .B(net8180));
 sg13g2_o21ai_1 _23615_ (.B1(_14340_),
    .Y(_00505_),
    .A1(net7610),
    .A2(net8180));
 sg13g2_nand2_1 _23616_ (.Y(_14341_),
    .A(net3905),
    .B(net8178));
 sg13g2_o21ai_1 _23617_ (.B1(_14341_),
    .Y(_00506_),
    .A1(net7589),
    .A2(net8178));
 sg13g2_nand2_1 _23618_ (.Y(_14342_),
    .A(net2919),
    .B(net8176));
 sg13g2_o21ai_1 _23619_ (.B1(_14342_),
    .Y(_00507_),
    .A1(net7600),
    .A2(net8176));
 sg13g2_nand2_1 _23620_ (.Y(_14343_),
    .A(net3150),
    .B(net8179));
 sg13g2_o21ai_1 _23621_ (.B1(_14343_),
    .Y(_00508_),
    .A1(net7594),
    .A2(net8179));
 sg13g2_nand2_1 _23622_ (.Y(_14344_),
    .A(net3637),
    .B(net8171));
 sg13g2_o21ai_1 _23623_ (.B1(_14344_),
    .Y(_00509_),
    .A1(net7602),
    .A2(net8171));
 sg13g2_nand2_1 _23624_ (.Y(_14345_),
    .A(net3272),
    .B(net8177));
 sg13g2_o21ai_1 _23625_ (.B1(_14345_),
    .Y(_00510_),
    .A1(net7560),
    .A2(net8177));
 sg13g2_nand2_1 _23626_ (.Y(_14346_),
    .A(net2981),
    .B(net8181));
 sg13g2_o21ai_1 _23627_ (.B1(_14346_),
    .Y(_00511_),
    .A1(net7574),
    .A2(net8181));
 sg13g2_nand2_1 _23628_ (.Y(_14347_),
    .A(net3391),
    .B(net8180));
 sg13g2_o21ai_1 _23629_ (.B1(_14347_),
    .Y(_00512_),
    .A1(net7549),
    .A2(net8180));
 sg13g2_nand2_1 _23630_ (.Y(_14348_),
    .A(net2738),
    .B(net8172));
 sg13g2_o21ai_1 _23631_ (.B1(_14348_),
    .Y(_00513_),
    .A1(net7570),
    .A2(net8172));
 sg13g2_nand2_1 _23632_ (.Y(_14349_),
    .A(net2842),
    .B(net8179));
 sg13g2_o21ai_1 _23633_ (.B1(_14349_),
    .Y(_00514_),
    .A1(net7544),
    .A2(net8179));
 sg13g2_nand2_1 _23634_ (.Y(_14350_),
    .A(net2657),
    .B(net8181));
 sg13g2_o21ai_1 _23635_ (.B1(_14350_),
    .Y(_00515_),
    .A1(net7555),
    .A2(net8181));
 sg13g2_nand2_1 _23636_ (.Y(_14351_),
    .A(net2626),
    .B(net8174));
 sg13g2_o21ai_1 _23637_ (.B1(_14351_),
    .Y(_00516_),
    .A1(net7584),
    .A2(net8174));
 sg13g2_nand2_1 _23638_ (.Y(_14352_),
    .A(net2992),
    .B(net8172));
 sg13g2_o21ai_1 _23639_ (.B1(_14352_),
    .Y(_00517_),
    .A1(net7563),
    .A2(net8172));
 sg13g2_nand2_1 _23640_ (.Y(_14353_),
    .A(net3112),
    .B(net8171));
 sg13g2_o21ai_1 _23641_ (.B1(_14353_),
    .Y(_00518_),
    .A1(net7522),
    .A2(net8171));
 sg13g2_nand2_1 _23642_ (.Y(_14354_),
    .A(net2632),
    .B(net8171));
 sg13g2_o21ai_1 _23643_ (.B1(_14354_),
    .Y(_00519_),
    .A1(net7535),
    .A2(net8171));
 sg13g2_nand2_1 _23644_ (.Y(_14355_),
    .A(net2953),
    .B(net8171));
 sg13g2_o21ai_1 _23645_ (.B1(_14355_),
    .Y(_00520_),
    .A1(net7528),
    .A2(net8171));
 sg13g2_nand2_1 _23646_ (.Y(_14356_),
    .A(net2676),
    .B(net8174));
 sg13g2_o21ai_1 _23647_ (.B1(_14356_),
    .Y(_00521_),
    .A1(net7520),
    .A2(net8174));
 sg13g2_nand2_1 _23648_ (.Y(_14357_),
    .A(net2699),
    .B(net8178));
 sg13g2_o21ai_1 _23649_ (.B1(_14357_),
    .Y(_00522_),
    .A1(net7507),
    .A2(net8178));
 sg13g2_nand2_1 _23650_ (.Y(_14358_),
    .A(net2844),
    .B(net8176));
 sg13g2_o21ai_1 _23651_ (.B1(_14358_),
    .Y(_00523_),
    .A1(net7514),
    .A2(net8176));
 sg13g2_nand2_1 _23652_ (.Y(_14359_),
    .A(net2900),
    .B(net8179));
 sg13g2_o21ai_1 _23653_ (.B1(_14359_),
    .Y(_00524_),
    .A1(net7495),
    .A2(net8179));
 sg13g2_nand2_1 _23654_ (.Y(_14360_),
    .A(net2625),
    .B(net8172));
 sg13g2_o21ai_1 _23655_ (.B1(_14360_),
    .Y(_00525_),
    .A1(net7500),
    .A2(net8172));
 sg13g2_nand2_1 _23656_ (.Y(_14361_),
    .A(net2671),
    .B(net8176));
 sg13g2_o21ai_1 _23657_ (.B1(_14361_),
    .Y(_00526_),
    .A1(net7643),
    .A2(net8176));
 sg13g2_nand2_1 _23658_ (.Y(_14362_),
    .A(net3642),
    .B(net8176));
 sg13g2_o21ai_1 _23659_ (.B1(_14362_),
    .Y(_00527_),
    .A1(net7648),
    .A2(net8176));
 sg13g2_nand2_1 _23660_ (.Y(_14363_),
    .A(net3058),
    .B(net8179));
 sg13g2_o21ai_1 _23661_ (.B1(_14363_),
    .Y(_00528_),
    .A1(net7654),
    .A2(net8179));
 sg13g2_nand2_1 _23662_ (.Y(_14364_),
    .A(net2748),
    .B(net8174));
 sg13g2_o21ai_1 _23663_ (.B1(_14364_),
    .Y(_00529_),
    .A1(net7661),
    .A2(net8174));
 sg13g2_nand2_1 _23664_ (.Y(_14365_),
    .A(net2713),
    .B(net8174));
 sg13g2_o21ai_1 _23665_ (.B1(_14365_),
    .Y(_00530_),
    .A1(net7640),
    .A2(net8174));
 sg13g2_nand2_1 _23666_ (.Y(_14366_),
    .A(net3174),
    .B(net8177));
 sg13g2_o21ai_1 _23667_ (.B1(_14366_),
    .Y(_00531_),
    .A1(net7628),
    .A2(net8177));
 sg13g2_nand2_1 _23668_ (.Y(_14367_),
    .A(net2789),
    .B(net8175));
 sg13g2_o21ai_1 _23669_ (.B1(_14367_),
    .Y(_00532_),
    .A1(net7622),
    .A2(net8175));
 sg13g2_nand2_1 _23670_ (.Y(_14368_),
    .A(net3467),
    .B(net8173));
 sg13g2_o21ai_1 _23671_ (.B1(_14368_),
    .Y(_00533_),
    .A1(net7634),
    .A2(net8173));
 sg13g2_nand2_1 _23672_ (.Y(_14369_),
    .A(net9709),
    .B(net8372));
 sg13g2_nor2_2 _23673_ (.A(_14164_),
    .B(_14369_),
    .Y(_14370_));
 sg13g2_nand2_1 _23674_ (.Y(_14371_),
    .A(net8961),
    .B(_14370_));
 sg13g2_nand2_1 _23675_ (.Y(_14372_),
    .A(net2962),
    .B(net7901));
 sg13g2_o21ai_1 _23676_ (.B1(_14372_),
    .Y(_00534_),
    .A1(net7486),
    .A2(net7901));
 sg13g2_nand2_1 _23677_ (.Y(_14373_),
    .A(net2906),
    .B(net7898));
 sg13g2_o21ai_1 _23678_ (.B1(_14373_),
    .Y(_00535_),
    .A1(net7664),
    .A2(net7898));
 sg13g2_nand2_1 _23679_ (.Y(_14374_),
    .A(net2955),
    .B(net7900));
 sg13g2_o21ai_1 _23680_ (.B1(_14374_),
    .Y(_00536_),
    .A1(net7614),
    .A2(net7898));
 sg13g2_nand2_1 _23681_ (.Y(_14375_),
    .A(net3200),
    .B(net7900));
 sg13g2_o21ai_1 _23682_ (.B1(_14375_),
    .Y(_00537_),
    .A1(net7607),
    .A2(net7899));
 sg13g2_nand2_1 _23683_ (.Y(_14376_),
    .A(net3128),
    .B(net7901));
 sg13g2_o21ai_1 _23684_ (.B1(_14376_),
    .Y(_00538_),
    .A1(net7589),
    .A2(net7901));
 sg13g2_nand2_1 _23685_ (.Y(_14377_),
    .A(net3111),
    .B(net7902));
 sg13g2_o21ai_1 _23686_ (.B1(_14377_),
    .Y(_00539_),
    .A1(net7600),
    .A2(net7902));
 sg13g2_nand2_1 _23687_ (.Y(_14378_),
    .A(net2917),
    .B(net7899));
 sg13g2_o21ai_1 _23688_ (.B1(_14378_),
    .Y(_00540_),
    .A1(net7592),
    .A2(net7899));
 sg13g2_nand2_1 _23689_ (.Y(_14379_),
    .A(net3039),
    .B(net7895));
 sg13g2_o21ai_1 _23690_ (.B1(_14379_),
    .Y(_00541_),
    .A1(net7604),
    .A2(net7895));
 sg13g2_nand2_1 _23691_ (.Y(_14380_),
    .A(net3464),
    .B(net7902));
 sg13g2_o21ai_1 _23692_ (.B1(_14380_),
    .Y(_00542_),
    .A1(net7558),
    .A2(net7902));
 sg13g2_nand2_1 _23693_ (.Y(_14381_),
    .A(net3120),
    .B(net7899));
 sg13g2_o21ai_1 _23694_ (.B1(_14381_),
    .Y(_00543_),
    .A1(net7574),
    .A2(net7898));
 sg13g2_nand2_1 _23695_ (.Y(_14382_),
    .A(net3297),
    .B(net7900));
 sg13g2_o21ai_1 _23696_ (.B1(_14382_),
    .Y(_00544_),
    .A1(net7546),
    .A2(net7900));
 sg13g2_nand2_1 _23697_ (.Y(_14383_),
    .A(net3492),
    .B(net7893));
 sg13g2_o21ai_1 _23698_ (.B1(_14383_),
    .Y(_00545_),
    .A1(net7571),
    .A2(net7893));
 sg13g2_nand2_1 _23699_ (.Y(_14384_),
    .A(net3300),
    .B(net7898));
 sg13g2_o21ai_1 _23700_ (.B1(_14384_),
    .Y(_00546_),
    .A1(net7542),
    .A2(net7898));
 sg13g2_nand2_1 _23701_ (.Y(_14385_),
    .A(net3165),
    .B(net7898));
 sg13g2_o21ai_1 _23702_ (.B1(_14385_),
    .Y(_00547_),
    .A1(net7551),
    .A2(net7898));
 sg13g2_nand2_1 _23703_ (.Y(_14386_),
    .A(net3170),
    .B(net7896));
 sg13g2_o21ai_1 _23704_ (.B1(_14386_),
    .Y(_00548_),
    .A1(net7581),
    .A2(net7896));
 sg13g2_nand2_1 _23705_ (.Y(_14387_),
    .A(net3347),
    .B(net7893));
 sg13g2_o21ai_1 _23706_ (.B1(_14387_),
    .Y(_00549_),
    .A1(net7565),
    .A2(net7893));
 sg13g2_nand2_1 _23707_ (.Y(_14388_),
    .A(net3196),
    .B(net7893));
 sg13g2_o21ai_1 _23708_ (.B1(_14388_),
    .Y(_00550_),
    .A1(net7524),
    .A2(net7893));
 sg13g2_nand2_1 _23709_ (.Y(_14389_),
    .A(net2885),
    .B(net7893));
 sg13g2_o21ai_1 _23710_ (.B1(_14389_),
    .Y(_00551_),
    .A1(net7538),
    .A2(net7893));
 sg13g2_nand2_1 _23711_ (.Y(_14390_),
    .A(net3963),
    .B(net7895));
 sg13g2_o21ai_1 _23712_ (.B1(_14390_),
    .Y(_00552_),
    .A1(net7530),
    .A2(net7895));
 sg13g2_nand2_1 _23713_ (.Y(_14391_),
    .A(net3602),
    .B(net7896));
 sg13g2_o21ai_1 _23714_ (.B1(_14391_),
    .Y(_00553_),
    .A1(net7521),
    .A2(net7896));
 sg13g2_nand2_1 _23715_ (.Y(_14392_),
    .A(net3047),
    .B(net7901));
 sg13g2_o21ai_1 _23716_ (.B1(_14392_),
    .Y(_00554_),
    .A1(net7508),
    .A2(net7901));
 sg13g2_nand2_1 _23717_ (.Y(_14393_),
    .A(net3180),
    .B(net7897));
 sg13g2_o21ai_1 _23718_ (.B1(_14393_),
    .Y(_00555_),
    .A1(net7511),
    .A2(net7897));
 sg13g2_nand2_1 _23719_ (.Y(_14394_),
    .A(net2935),
    .B(net7899));
 sg13g2_o21ai_1 _23720_ (.B1(_14394_),
    .Y(_00556_),
    .A1(net7498),
    .A2(net7899));
 sg13g2_nand2_1 _23721_ (.Y(_14395_),
    .A(net3865),
    .B(net7894));
 sg13g2_o21ai_1 _23722_ (.B1(_14395_),
    .Y(_00557_),
    .A1(net7500),
    .A2(net7894));
 sg13g2_nand2_1 _23723_ (.Y(_14396_),
    .A(net3516),
    .B(net7902));
 sg13g2_o21ai_1 _23724_ (.B1(_14396_),
    .Y(_00558_),
    .A1(net7642),
    .A2(net7902));
 sg13g2_nand2_1 _23725_ (.Y(_14397_),
    .A(net3488),
    .B(net7901));
 sg13g2_o21ai_1 _23726_ (.B1(_14397_),
    .Y(_00559_),
    .A1(net7651),
    .A2(net7901));
 sg13g2_nand2_1 _23727_ (.Y(_14398_),
    .A(net2837),
    .B(net7899));
 sg13g2_o21ai_1 _23728_ (.B1(_14398_),
    .Y(_00560_),
    .A1(net7653),
    .A2(net7899));
 sg13g2_nand2_1 _23729_ (.Y(_14399_),
    .A(net3344),
    .B(net7897));
 sg13g2_o21ai_1 _23730_ (.B1(_14399_),
    .Y(_00561_),
    .A1(net7660),
    .A2(net7897));
 sg13g2_nand2_1 _23731_ (.Y(_14400_),
    .A(net2918),
    .B(net7897));
 sg13g2_o21ai_1 _23732_ (.B1(_14400_),
    .Y(_00562_),
    .A1(net7636),
    .A2(net7897));
 sg13g2_nand2_1 _23733_ (.Y(_14401_),
    .A(net3354),
    .B(net7902));
 sg13g2_o21ai_1 _23734_ (.B1(_14401_),
    .Y(_00563_),
    .A1(net7626),
    .A2(net7902));
 sg13g2_nand2_1 _23735_ (.Y(_14402_),
    .A(net3534),
    .B(net7897));
 sg13g2_o21ai_1 _23736_ (.B1(_14402_),
    .Y(_00564_),
    .A1(net7619),
    .A2(net7903));
 sg13g2_nand2_1 _23737_ (.Y(_14403_),
    .A(net2846),
    .B(net7894));
 sg13g2_o21ai_1 _23738_ (.B1(_14403_),
    .Y(_00565_),
    .A1(net7632),
    .A2(net7894));
 sg13g2_nand3_1 _23739_ (.B(_14130_),
    .C(_14199_),
    .A(net8371),
    .Y(_14404_));
 sg13g2_nand2_1 _23740_ (.Y(_14405_),
    .A(net3835),
    .B(net8169));
 sg13g2_o21ai_1 _23741_ (.B1(_14405_),
    .Y(_00566_),
    .A1(net7488),
    .A2(net8169));
 sg13g2_nand2_1 _23742_ (.Y(_14406_),
    .A(net3729),
    .B(net8169));
 sg13g2_o21ai_1 _23743_ (.B1(_14406_),
    .Y(_00567_),
    .A1(net7663),
    .A2(net8169));
 sg13g2_nand2_1 _23744_ (.Y(_14407_),
    .A(net3567),
    .B(net8169));
 sg13g2_o21ai_1 _23745_ (.B1(_14407_),
    .Y(_00568_),
    .A1(net7612),
    .A2(net8169));
 sg13g2_nand2_1 _23746_ (.Y(_14408_),
    .A(net3882),
    .B(net8167));
 sg13g2_o21ai_1 _23747_ (.B1(_14408_),
    .Y(_00569_),
    .A1(net7609),
    .A2(net8167));
 sg13g2_nand2_1 _23748_ (.Y(_14409_),
    .A(net3798),
    .B(net8164));
 sg13g2_o21ai_1 _23749_ (.B1(_14409_),
    .Y(_00570_),
    .A1(net7586),
    .A2(net8164));
 sg13g2_nand2_1 _23750_ (.Y(_14410_),
    .A(net3238),
    .B(net8164));
 sg13g2_o21ai_1 _23751_ (.B1(_14410_),
    .Y(_00571_),
    .A1(net7598),
    .A2(net8164));
 sg13g2_nand2_1 _23752_ (.Y(_14411_),
    .A(net3498),
    .B(net8166));
 sg13g2_o21ai_1 _23753_ (.B1(_14411_),
    .Y(_00572_),
    .A1(net7594),
    .A2(net8166));
 sg13g2_nand2_1 _23754_ (.Y(_14412_),
    .A(net3902),
    .B(net8160));
 sg13g2_o21ai_1 _23755_ (.B1(_14412_),
    .Y(_00573_),
    .A1(net7602),
    .A2(net8160));
 sg13g2_nand2_1 _23756_ (.Y(_14413_),
    .A(net3433),
    .B(net8165));
 sg13g2_o21ai_1 _23757_ (.B1(_14413_),
    .Y(_00574_),
    .A1(net7557),
    .A2(net8165));
 sg13g2_nand2_1 _23758_ (.Y(_14414_),
    .A(net3437),
    .B(net8168));
 sg13g2_o21ai_1 _23759_ (.B1(_14414_),
    .Y(_00575_),
    .A1(net7576),
    .A2(net8168));
 sg13g2_nand2_1 _23760_ (.Y(_14415_),
    .A(net3046),
    .B(net8166));
 sg13g2_o21ai_1 _23761_ (.B1(_14415_),
    .Y(_00576_),
    .A1(net7550),
    .A2(net8166));
 sg13g2_nand2_1 _23762_ (.Y(_14416_),
    .A(net4044),
    .B(net8160));
 sg13g2_o21ai_1 _23763_ (.B1(_14416_),
    .Y(_00577_),
    .A1(net7568),
    .A2(net8160));
 sg13g2_nand2_1 _23764_ (.Y(_14417_),
    .A(net4022),
    .B(net8166));
 sg13g2_o21ai_1 _23765_ (.B1(_14417_),
    .Y(_00578_),
    .A1(net7543),
    .A2(net8166));
 sg13g2_nand2_1 _23766_ (.Y(_14418_),
    .A(net3011),
    .B(net8168));
 sg13g2_o21ai_1 _23767_ (.B1(_14418_),
    .Y(_00579_),
    .A1(net7552),
    .A2(net8168));
 sg13g2_nand2_1 _23768_ (.Y(_14419_),
    .A(net3443),
    .B(net8163));
 sg13g2_o21ai_1 _23769_ (.B1(_14419_),
    .Y(_00580_),
    .A1(net7585),
    .A2(net8163));
 sg13g2_nand2_1 _23770_ (.Y(_14420_),
    .A(net3273),
    .B(net8161));
 sg13g2_o21ai_1 _23771_ (.B1(_14420_),
    .Y(_00581_),
    .A1(net7564),
    .A2(net8161));
 sg13g2_nand2_1 _23772_ (.Y(_14421_),
    .A(net3855),
    .B(net8160));
 sg13g2_o21ai_1 _23773_ (.B1(_14421_),
    .Y(_00582_),
    .A1(net7522),
    .A2(net8160));
 sg13g2_nand2_1 _23774_ (.Y(_14422_),
    .A(net3763),
    .B(net8160));
 sg13g2_o21ai_1 _23775_ (.B1(_14422_),
    .Y(_00583_),
    .A1(net7535),
    .A2(net8160));
 sg13g2_nand2_1 _23776_ (.Y(_14423_),
    .A(net3987),
    .B(net8161));
 sg13g2_o21ai_1 _23777_ (.B1(_14423_),
    .Y(_00584_),
    .A1(net7528),
    .A2(net8161));
 sg13g2_nand2_1 _23778_ (.Y(_14424_),
    .A(net3751),
    .B(net8162));
 sg13g2_o21ai_1 _23779_ (.B1(_14424_),
    .Y(_00585_),
    .A1(net7518),
    .A2(net8162));
 sg13g2_nand2_1 _23780_ (.Y(_14425_),
    .A(net3296),
    .B(net8165));
 sg13g2_o21ai_1 _23781_ (.B1(_14425_),
    .Y(_00586_),
    .A1(net7505),
    .A2(net8165));
 sg13g2_nand2_1 _23782_ (.Y(_14426_),
    .A(net3723),
    .B(net8164));
 sg13g2_o21ai_1 _23783_ (.B1(_14426_),
    .Y(_00587_),
    .A1(net7513),
    .A2(net8164));
 sg13g2_nand2_1 _23784_ (.Y(_14427_),
    .A(net3316),
    .B(net8166));
 sg13g2_o21ai_1 _23785_ (.B1(_14427_),
    .Y(_00588_),
    .A1(net7496),
    .A2(net8166));
 sg13g2_nand2_1 _23786_ (.Y(_14428_),
    .A(net3945),
    .B(net8161));
 sg13g2_o21ai_1 _23787_ (.B1(_14428_),
    .Y(_00589_),
    .A1(net7500),
    .A2(net8161));
 sg13g2_nand2_1 _23788_ (.Y(_14429_),
    .A(net3735),
    .B(net8164));
 sg13g2_o21ai_1 _23789_ (.B1(_14429_),
    .Y(_00590_),
    .A1(net7643),
    .A2(net8164));
 sg13g2_nand2_1 _23790_ (.Y(_14430_),
    .A(net3288),
    .B(net8169));
 sg13g2_o21ai_1 _23791_ (.B1(_14430_),
    .Y(_00591_),
    .A1(net7650),
    .A2(net8169));
 sg13g2_nand2_1 _23792_ (.Y(_14431_),
    .A(net3678),
    .B(net8167));
 sg13g2_o21ai_1 _23793_ (.B1(_14431_),
    .Y(_00592_),
    .A1(net7655),
    .A2(net8167));
 sg13g2_nand2_1 _23794_ (.Y(_14432_),
    .A(net3657),
    .B(net8162));
 sg13g2_o21ai_1 _23795_ (.B1(_14432_),
    .Y(_00593_),
    .A1(net7659),
    .A2(net8162));
 sg13g2_nand2_1 _23796_ (.Y(_14433_),
    .A(net3660),
    .B(net8162));
 sg13g2_o21ai_1 _23797_ (.B1(_14433_),
    .Y(_00594_),
    .A1(net7636),
    .A2(net8162));
 sg13g2_nand2_1 _23798_ (.Y(_14434_),
    .A(net2925),
    .B(net8165));
 sg13g2_o21ai_1 _23799_ (.B1(_14434_),
    .Y(_00595_),
    .A1(net7625),
    .A2(net8165));
 sg13g2_nand2_1 _23800_ (.Y(_14435_),
    .A(net3809),
    .B(net8162));
 sg13g2_o21ai_1 _23801_ (.B1(_14435_),
    .Y(_00596_),
    .A1(net7621),
    .A2(net8162));
 sg13g2_nand2_1 _23802_ (.Y(_14436_),
    .A(net3600),
    .B(net8163));
 sg13g2_o21ai_1 _23803_ (.B1(_14436_),
    .Y(_00597_),
    .A1(net7631),
    .A2(net8163));
 sg13g2_a21oi_2 _23804_ (.B1(_13972_),
    .Y(_14437_),
    .A2(net8958),
    .A1(\soc_I.clint_I.addr[0] ));
 sg13g2_a21o_2 _23805_ (.A2(net8958),
    .A1(\soc_I.clint_I.addr[0] ),
    .B1(_13972_),
    .X(_14438_));
 sg13g2_nor2_2 _23806_ (.A(net7424),
    .B(_14438_),
    .Y(_14439_));
 sg13g2_nor3_1 _23807_ (.A(_12955_),
    .B(net7466),
    .C(_14438_),
    .Y(_14440_));
 sg13g2_o21ai_1 _23808_ (.B1(net9321),
    .Y(_14441_),
    .A1(net4592),
    .A2(net7436));
 sg13g2_a21oi_1 _23809_ (.A1(_13978_),
    .A2(net7436),
    .Y(_00598_),
    .B1(_14441_));
 sg13g2_o21ai_1 _23810_ (.B1(net9321),
    .Y(_14442_),
    .A1(net4945),
    .A2(net7436));
 sg13g2_a21oi_1 _23811_ (.A1(net8612),
    .A2(_14439_),
    .Y(_00599_),
    .B1(_14442_));
 sg13g2_o21ai_1 _23812_ (.B1(net9321),
    .Y(_14443_),
    .A1(net5005),
    .A2(net7436));
 sg13g2_a21oi_1 _23813_ (.A1(net8610),
    .A2(_14439_),
    .Y(_00600_),
    .B1(_14443_));
 sg13g2_o21ai_1 _23814_ (.B1(net9310),
    .Y(_14444_),
    .A1(net4662),
    .A2(net7435));
 sg13g2_a21oi_1 _23815_ (.A1(net8549),
    .A2(net7435),
    .Y(_00601_),
    .B1(_14444_));
 sg13g2_o21ai_1 _23816_ (.B1(net9310),
    .Y(_14445_),
    .A1(net4751),
    .A2(net7435));
 sg13g2_a21oi_1 _23817_ (.A1(net8608),
    .A2(_14439_),
    .Y(_00602_),
    .B1(_14445_));
 sg13g2_o21ai_1 _23818_ (.B1(net9310),
    .Y(_14446_),
    .A1(net4687),
    .A2(net7435));
 sg13g2_a21oi_1 _23819_ (.A1(net8606),
    .A2(_14439_),
    .Y(_00603_),
    .B1(_14446_));
 sg13g2_o21ai_1 _23820_ (.B1(net9309),
    .Y(_14447_),
    .A1(net4775),
    .A2(net7435));
 sg13g2_a21oi_1 _23821_ (.A1(net8604),
    .A2(net7435),
    .Y(_00604_),
    .B1(_14447_));
 sg13g2_o21ai_1 _23822_ (.B1(net9308),
    .Y(_14448_),
    .A1(net4754),
    .A2(net7435));
 sg13g2_a21oi_1 _23823_ (.A1(_14024_),
    .A2(net7435),
    .Y(_00605_),
    .B1(_14448_));
 sg13g2_nor3_2 _23824_ (.A(net7479),
    .B(net7425),
    .C(_13973_),
    .Y(_14449_));
 sg13g2_nand2_1 _23825_ (.Y(_14450_),
    .A(net7480),
    .B(net7452));
 sg13g2_nor2_2 _23826_ (.A(_13973_),
    .B(_14450_),
    .Y(_14451_));
 sg13g2_o21ai_1 _23827_ (.B1(net9308),
    .Y(_14452_),
    .A1(net4855),
    .A2(_14451_));
 sg13g2_a21oi_1 _23828_ (.A1(_13979_),
    .A2(_14449_),
    .Y(_00606_),
    .B1(_14452_));
 sg13g2_o21ai_1 _23829_ (.B1(net9308),
    .Y(_14453_),
    .A1(net4924),
    .A2(_14451_));
 sg13g2_a21oi_1 _23830_ (.A1(_13988_),
    .A2(_14449_),
    .Y(_00607_),
    .B1(_14453_));
 sg13g2_o21ai_1 _23831_ (.B1(net9300),
    .Y(_14454_),
    .A1(net4860),
    .A2(_14451_));
 sg13g2_a21oi_1 _23832_ (.A1(_13995_),
    .A2(_14449_),
    .Y(_00608_),
    .B1(_14454_));
 sg13g2_o21ai_1 _23833_ (.B1(net9311),
    .Y(_14455_),
    .A1(net4870),
    .A2(_14451_));
 sg13g2_a21oi_1 _23834_ (.A1(_14001_),
    .A2(_14449_),
    .Y(_00609_),
    .B1(_14455_));
 sg13g2_o21ai_1 _23835_ (.B1(net9300),
    .Y(_14456_),
    .A1(net4273),
    .A2(_14451_));
 sg13g2_a21oi_1 _23836_ (.A1(_14007_),
    .A2(_14449_),
    .Y(_00610_),
    .B1(_14456_));
 sg13g2_o21ai_1 _23837_ (.B1(net9315),
    .Y(_14457_),
    .A1(net4955),
    .A2(_14451_));
 sg13g2_a21oi_1 _23838_ (.A1(_14014_),
    .A2(_14449_),
    .Y(_00611_),
    .B1(_14457_));
 sg13g2_o21ai_1 _23839_ (.B1(net9316),
    .Y(_14458_),
    .A1(net4804),
    .A2(_14451_));
 sg13g2_a21oi_1 _23840_ (.A1(_14020_),
    .A2(_14449_),
    .Y(_00612_),
    .B1(_14458_));
 sg13g2_o21ai_1 _23841_ (.B1(net9315),
    .Y(_14459_),
    .A1(net4908),
    .A2(_14451_));
 sg13g2_a21oi_1 _23842_ (.A1(_14029_),
    .A2(_14449_),
    .Y(_00613_),
    .B1(_14459_));
 sg13g2_nor4_1 _23843_ (.A(net7479),
    .B(_12955_),
    .C(net7466),
    .D(_14033_),
    .Y(_14460_));
 sg13g2_nor2_1 _23844_ (.A(_14033_),
    .B(_14450_),
    .Y(_14461_));
 sg13g2_o21ai_1 _23845_ (.B1(net9315),
    .Y(_14462_),
    .A1(net4938),
    .A2(net7421));
 sg13g2_a21oi_1 _23846_ (.A1(_14037_),
    .A2(net7397),
    .Y(_00614_),
    .B1(_14462_));
 sg13g2_nand2_1 _23847_ (.Y(_14463_),
    .A(_14041_),
    .B(net7397));
 sg13g2_o21ai_1 _23848_ (.B1(_14463_),
    .Y(_14464_),
    .A1(net4837),
    .A2(net7421));
 sg13g2_nor2_1 _23849_ (.A(net9008),
    .B(_14464_),
    .Y(_00615_));
 sg13g2_nand2_1 _23850_ (.Y(_14465_),
    .A(_14046_),
    .B(net7397));
 sg13g2_o21ai_1 _23851_ (.B1(_14465_),
    .Y(_14466_),
    .A1(net4865),
    .A2(net7421));
 sg13g2_nor2_1 _23852_ (.A(net9008),
    .B(_14466_),
    .Y(_00616_));
 sg13g2_nor2_1 _23853_ (.A(net4225),
    .B(net7421),
    .Y(_14467_));
 sg13g2_a21oi_1 _23854_ (.A1(_14051_),
    .A2(net7421),
    .Y(_14468_),
    .B1(net9009));
 sg13g2_nor2b_1 _23855_ (.A(_14467_),
    .B_N(_14468_),
    .Y(_00617_));
 sg13g2_nand2_1 _23856_ (.Y(_14469_),
    .A(_14056_),
    .B(net7397));
 sg13g2_o21ai_1 _23857_ (.B1(_14469_),
    .Y(_14470_),
    .A1(net4956),
    .A2(net7423));
 sg13g2_nor2_1 _23858_ (.A(net9008),
    .B(_14470_),
    .Y(_00618_));
 sg13g2_nand2_1 _23859_ (.Y(_14471_),
    .A(_14060_),
    .B(net7398));
 sg13g2_o21ai_1 _23860_ (.B1(_14471_),
    .Y(_02781_),
    .A1(net4842),
    .A2(net7422));
 sg13g2_nor2_1 _23861_ (.A(net9010),
    .B(_02781_),
    .Y(_00619_));
 sg13g2_nand2_1 _23862_ (.Y(_02782_),
    .A(_14065_),
    .B(net7398));
 sg13g2_o21ai_1 _23863_ (.B1(_02782_),
    .Y(_02783_),
    .A1(net5085),
    .A2(net7422));
 sg13g2_nor2_1 _23864_ (.A(net9010),
    .B(_02783_),
    .Y(_00620_));
 sg13g2_mux2_1 _23865_ (.A0(_10561_),
    .A1(_14070_),
    .S(net7397),
    .X(_02784_));
 sg13g2_nor2_1 _23866_ (.A(net9021),
    .B(_02784_),
    .Y(_00621_));
 sg13g2_nand2_1 _23867_ (.Y(_02785_),
    .A(_14076_),
    .B(net7398));
 sg13g2_o21ai_1 _23868_ (.B1(_02785_),
    .Y(_02786_),
    .A1(net5078),
    .A2(net7422));
 sg13g2_nor2_1 _23869_ (.A(net9011),
    .B(_02786_),
    .Y(_00622_));
 sg13g2_o21ai_1 _23870_ (.B1(net9319),
    .Y(_02787_),
    .A1(net5095),
    .A2(net7423));
 sg13g2_a21oi_1 _23871_ (.A1(_14082_),
    .A2(net7423),
    .Y(_00623_),
    .B1(_02787_));
 sg13g2_nand2_1 _23872_ (.Y(_02788_),
    .A(_14088_),
    .B(net7398));
 sg13g2_o21ai_1 _23873_ (.B1(_02788_),
    .Y(_02789_),
    .A1(net5136),
    .A2(net7422));
 sg13g2_nor2_1 _23874_ (.A(net9011),
    .B(_02789_),
    .Y(_00624_));
 sg13g2_o21ai_1 _23875_ (.B1(net9328),
    .Y(_02790_),
    .A1(net4737),
    .A2(net7422));
 sg13g2_a21oi_1 _23876_ (.A1(_14092_),
    .A2(net7422),
    .Y(_00625_),
    .B1(_02790_));
 sg13g2_nand2_1 _23877_ (.Y(_02791_),
    .A(_14099_),
    .B(net7397));
 sg13g2_o21ai_1 _23878_ (.B1(_02791_),
    .Y(_02792_),
    .A1(net4832),
    .A2(net7421));
 sg13g2_nor2_1 _23879_ (.A(net9008),
    .B(_02792_),
    .Y(_00626_));
 sg13g2_nand2_1 _23880_ (.Y(_02793_),
    .A(_14104_),
    .B(net7397));
 sg13g2_o21ai_1 _23881_ (.B1(_02793_),
    .Y(_02794_),
    .A1(net4830),
    .A2(net7421));
 sg13g2_nor2_1 _23882_ (.A(net9009),
    .B(_02794_),
    .Y(_00627_));
 sg13g2_o21ai_1 _23883_ (.B1(net9327),
    .Y(_02795_),
    .A1(net4895),
    .A2(net7422));
 sg13g2_a21oi_1 _23884_ (.A1(_14111_),
    .A2(net7422),
    .Y(_00628_),
    .B1(_02795_));
 sg13g2_nand2_1 _23885_ (.Y(_02796_),
    .A(_14116_),
    .B(net7397));
 sg13g2_o21ai_1 _23886_ (.B1(_02796_),
    .Y(_02797_),
    .A1(net4979),
    .A2(net7421));
 sg13g2_nor2_1 _23887_ (.A(net9013),
    .B(_02797_),
    .Y(_00629_));
 sg13g2_nor2_2 _23888_ (.A(\soc_I.rx_uart_i.fifo_i.wr_ptr[3] ),
    .B(net9273),
    .Y(_02798_));
 sg13g2_nand2_1 _23889_ (.Y(_02799_),
    .A(_14122_),
    .B(_02798_));
 sg13g2_nand2_1 _23890_ (.Y(_02800_),
    .A(net2658),
    .B(net8547));
 sg13g2_o21ai_1 _23891_ (.B1(_02800_),
    .Y(_00630_),
    .A1(net9170),
    .A2(net8547));
 sg13g2_mux2_1 _23892_ (.A0(\soc_I.rx_uart_i.fifo_i.din[1] ),
    .A1(net4328),
    .S(net8547),
    .X(_00631_));
 sg13g2_mux2_1 _23893_ (.A0(net3981),
    .A1(\soc_I.rx_uart_i.fifo_i.ram[0][2] ),
    .S(_02799_),
    .X(_00632_));
 sg13g2_mux2_1 _23894_ (.A0(\soc_I.rx_uart_i.fifo_i.din[3] ),
    .A1(net4142),
    .S(net8547),
    .X(_00633_));
 sg13g2_mux2_1 _23895_ (.A0(net9283),
    .A1(net4214),
    .S(net8547),
    .X(_00634_));
 sg13g2_mux2_1 _23896_ (.A0(net9279),
    .A1(net4024),
    .S(net8547),
    .X(_00635_));
 sg13g2_mux2_1 _23897_ (.A0(net9278),
    .A1(net4127),
    .S(net8547),
    .X(_00636_));
 sg13g2_mux2_1 _23898_ (.A0(net9275),
    .A1(net4047),
    .S(net8547),
    .X(_00637_));
 sg13g2_nor3_2 _23899_ (.A(_10391_),
    .B(\soc_I.rx_uart_i.fifo_i.wr_ptr[0] ),
    .C(_14121_),
    .Y(_02801_));
 sg13g2_nor2b_2 _23900_ (.A(\soc_I.rx_uart_i.fifo_i.wr_ptr[2] ),
    .B_N(\soc_I.rx_uart_i.fifo_i.wr_ptr[3] ),
    .Y(_02802_));
 sg13g2_nand2_1 _23901_ (.Y(_02803_),
    .A(_02801_),
    .B(_02802_));
 sg13g2_nand2_1 _23902_ (.Y(_02804_),
    .A(net2744),
    .B(_02803_));
 sg13g2_o21ai_1 _23903_ (.B1(_02804_),
    .Y(_00638_),
    .A1(net9171),
    .A2(net8546));
 sg13g2_mux2_1 _23904_ (.A0(net9289),
    .A1(net3639),
    .S(net8546),
    .X(_00639_));
 sg13g2_mux2_1 _23905_ (.A0(net9286),
    .A1(net3540),
    .S(net8546),
    .X(_00640_));
 sg13g2_mux2_1 _23906_ (.A0(net9285),
    .A1(net4161),
    .S(net8546),
    .X(_00641_));
 sg13g2_mux2_1 _23907_ (.A0(net9282),
    .A1(net3752),
    .S(net8546),
    .X(_00642_));
 sg13g2_mux2_1 _23908_ (.A0(net9280),
    .A1(net3609),
    .S(net8546),
    .X(_00643_));
 sg13g2_mux2_1 _23909_ (.A0(\soc_I.rx_uart_i.fifo_i.din[6] ),
    .A1(net4104),
    .S(net8546),
    .X(_00644_));
 sg13g2_mux2_1 _23910_ (.A0(net9276),
    .A1(net4077),
    .S(net8546),
    .X(_00645_));
 sg13g2_and3_2 _23911_ (.X(_02805_),
    .A(\soc_I.rx_uart_i.fifo_i.wr_ptr[1] ),
    .B(\soc_I.rx_uart_i.fifo_i.wr_ptr[0] ),
    .C(_14120_));
 sg13g2_nand2_1 _23912_ (.Y(_02806_),
    .A(_02802_),
    .B(_02805_));
 sg13g2_nand2_1 _23913_ (.Y(_02807_),
    .A(net2709),
    .B(_02806_));
 sg13g2_o21ai_1 _23914_ (.B1(net2710),
    .Y(_00646_),
    .A1(net9171),
    .A2(net8600));
 sg13g2_mux2_1 _23915_ (.A0(net9289),
    .A1(net4212),
    .S(net8600),
    .X(_00647_));
 sg13g2_mux2_1 _23916_ (.A0(net9286),
    .A1(net4050),
    .S(net8600),
    .X(_00648_));
 sg13g2_mux2_1 _23917_ (.A0(net9285),
    .A1(net3912),
    .S(net8600),
    .X(_00649_));
 sg13g2_mux2_1 _23918_ (.A0(net9282),
    .A1(net4219),
    .S(net8600),
    .X(_00650_));
 sg13g2_mux2_1 _23919_ (.A0(net9280),
    .A1(net4099),
    .S(net8600),
    .X(_00651_));
 sg13g2_mux2_1 _23920_ (.A0(\soc_I.rx_uart_i.fifo_i.din[6] ),
    .A1(net4237),
    .S(net8600),
    .X(_00652_));
 sg13g2_mux2_1 _23921_ (.A0(net9276),
    .A1(net3965),
    .S(net8600),
    .X(_00653_));
 sg13g2_nand3_1 _23922_ (.B(net9273),
    .C(_14122_),
    .A(\soc_I.rx_uart_i.fifo_i.wr_ptr[3] ),
    .Y(_02808_));
 sg13g2_nand2_1 _23923_ (.Y(_02809_),
    .A(net2647),
    .B(_02808_));
 sg13g2_o21ai_1 _23924_ (.B1(net2648),
    .Y(_00654_),
    .A1(net9171),
    .A2(net8545));
 sg13g2_mux2_1 _23925_ (.A0(net9288),
    .A1(net4049),
    .S(net8545),
    .X(_00655_));
 sg13g2_mux2_1 _23926_ (.A0(net9286),
    .A1(net3832),
    .S(net8545),
    .X(_00656_));
 sg13g2_mux2_1 _23927_ (.A0(net9285),
    .A1(net4192),
    .S(net8545),
    .X(_00657_));
 sg13g2_mux2_1 _23928_ (.A0(net9282),
    .A1(net4109),
    .S(net8545),
    .X(_00658_));
 sg13g2_mux2_1 _23929_ (.A0(net9279),
    .A1(net3812),
    .S(net8545),
    .X(_00659_));
 sg13g2_mux2_1 _23930_ (.A0(net9277),
    .A1(net4240),
    .S(net8545),
    .X(_00660_));
 sg13g2_mux2_1 _23931_ (.A0(net9275),
    .A1(net4154),
    .S(net8545),
    .X(_00661_));
 sg13g2_and3_2 _23932_ (.X(_02810_),
    .A(_10391_),
    .B(\soc_I.rx_uart_i.fifo_i.wr_ptr[0] ),
    .C(net8819));
 sg13g2_and3_1 _23933_ (.X(_02811_),
    .A(\soc_I.rx_uart_i.fifo_i.wr_ptr[3] ),
    .B(net9273),
    .C(_02810_));
 sg13g2_nor2_1 _23934_ (.A(net3384),
    .B(net8599),
    .Y(_02812_));
 sg13g2_a21oi_1 _23935_ (.A1(net9171),
    .A2(_02811_),
    .Y(_00662_),
    .B1(_02812_));
 sg13g2_mux2_1 _23936_ (.A0(net3353),
    .A1(net9288),
    .S(net8599),
    .X(_00663_));
 sg13g2_mux2_1 _23937_ (.A0(net3195),
    .A1(net9286),
    .S(net8599),
    .X(_00664_));
 sg13g2_mux2_1 _23938_ (.A0(net3431),
    .A1(net9285),
    .S(net8599),
    .X(_00665_));
 sg13g2_mux2_1 _23939_ (.A0(net3130),
    .A1(net9282),
    .S(net8599),
    .X(_00666_));
 sg13g2_mux2_1 _23940_ (.A0(net3438),
    .A1(net9279),
    .S(net8599),
    .X(_00667_));
 sg13g2_mux2_1 _23941_ (.A0(net3362),
    .A1(net9277),
    .S(net8599),
    .X(_00668_));
 sg13g2_mux2_1 _23942_ (.A0(net3168),
    .A1(net9275),
    .S(net8599),
    .X(_00669_));
 sg13g2_and3_1 _23943_ (.X(_02813_),
    .A(\soc_I.rx_uart_i.fifo_i.wr_ptr[3] ),
    .B(net9273),
    .C(_02801_));
 sg13g2_nor2_1 _23944_ (.A(net3984),
    .B(_02813_),
    .Y(_02814_));
 sg13g2_a21oi_1 _23945_ (.A1(_10396_),
    .A2(net8544),
    .Y(_00670_),
    .B1(net3985));
 sg13g2_mux2_1 _23946_ (.A0(net3619),
    .A1(net9288),
    .S(net8544),
    .X(_00671_));
 sg13g2_mux2_1 _23947_ (.A0(net2731),
    .A1(net9287),
    .S(net8544),
    .X(_00672_));
 sg13g2_mux2_1 _23948_ (.A0(net3259),
    .A1(net9285),
    .S(net8544),
    .X(_00673_));
 sg13g2_mux2_1 _23949_ (.A0(net3393),
    .A1(net9282),
    .S(net8544),
    .X(_00674_));
 sg13g2_mux2_1 _23950_ (.A0(net2771),
    .A1(net9279),
    .S(net8544),
    .X(_00675_));
 sg13g2_mux2_1 _23951_ (.A0(net3304),
    .A1(net9277),
    .S(net8544),
    .X(_00676_));
 sg13g2_mux2_1 _23952_ (.A0(net3551),
    .A1(net9275),
    .S(net8544),
    .X(_00677_));
 sg13g2_nand3_1 _23953_ (.B(net8372),
    .C(_14165_),
    .A(net8961),
    .Y(_02815_));
 sg13g2_nand2_1 _23954_ (.Y(_02816_),
    .A(net2847),
    .B(net8158));
 sg13g2_o21ai_1 _23955_ (.B1(_02816_),
    .Y(_00678_),
    .A1(net7489),
    .A2(net8158));
 sg13g2_nand2_1 _23956_ (.Y(_02817_),
    .A(net4030),
    .B(net8154));
 sg13g2_o21ai_1 _23957_ (.B1(_02817_),
    .Y(_00679_),
    .A1(net7663),
    .A2(net8154));
 sg13g2_nand2_1 _23958_ (.Y(_02818_),
    .A(net4270),
    .B(net8154));
 sg13g2_o21ai_1 _23959_ (.B1(_02818_),
    .Y(_00680_),
    .A1(net7617),
    .A2(net8154));
 sg13g2_nand2_1 _23960_ (.Y(_02819_),
    .A(net3279),
    .B(net8156));
 sg13g2_o21ai_1 _23961_ (.B1(_02819_),
    .Y(_00681_),
    .A1(net7610),
    .A2(net8156));
 sg13g2_nand2_1 _23962_ (.Y(_02820_),
    .A(net3266),
    .B(net8154));
 sg13g2_o21ai_1 _23963_ (.B1(_02820_),
    .Y(_00682_),
    .A1(net7588),
    .A2(net8154));
 sg13g2_nand2_1 _23964_ (.Y(_02821_),
    .A(net3355),
    .B(net8152));
 sg13g2_o21ai_1 _23965_ (.B1(_02821_),
    .Y(_00683_),
    .A1(net7597),
    .A2(net8152));
 sg13g2_nand2_1 _23966_ (.Y(_02822_),
    .A(net3280),
    .B(net8155));
 sg13g2_o21ai_1 _23967_ (.B1(_02822_),
    .Y(_00684_),
    .A1(net7595),
    .A2(net8155));
 sg13g2_nand2_1 _23968_ (.Y(_02823_),
    .A(net3584),
    .B(net8148));
 sg13g2_o21ai_1 _23969_ (.B1(_02823_),
    .Y(_00685_),
    .A1(net7602),
    .A2(net8148));
 sg13g2_nand2_1 _23970_ (.Y(_02824_),
    .A(net3287),
    .B(net8153));
 sg13g2_o21ai_1 _23971_ (.B1(_02824_),
    .Y(_00686_),
    .A1(net7557),
    .A2(net8153));
 sg13g2_nand2_1 _23972_ (.Y(_02825_),
    .A(net3004),
    .B(net8157));
 sg13g2_o21ai_1 _23973_ (.B1(_02825_),
    .Y(_00687_),
    .A1(net7574),
    .A2(net8157));
 sg13g2_nand2_1 _23974_ (.Y(_02826_),
    .A(net3624),
    .B(net8155));
 sg13g2_o21ai_1 _23975_ (.B1(_02826_),
    .Y(_00688_),
    .A1(net7549),
    .A2(net8155));
 sg13g2_nand2_1 _23976_ (.Y(_02827_),
    .A(net3650),
    .B(net8148));
 sg13g2_o21ai_1 _23977_ (.B1(_02827_),
    .Y(_00689_),
    .A1(net7569),
    .A2(net8148));
 sg13g2_nand2_1 _23978_ (.Y(_02828_),
    .A(net2888),
    .B(net8155));
 sg13g2_o21ai_1 _23979_ (.B1(_02828_),
    .Y(_00690_),
    .A1(net7544),
    .A2(net8155));
 sg13g2_nand2_1 _23980_ (.Y(_02829_),
    .A(net3020),
    .B(net8157));
 sg13g2_o21ai_1 _23981_ (.B1(_02829_),
    .Y(_00691_),
    .A1(net7553),
    .A2(net8157));
 sg13g2_nand2_1 _23982_ (.Y(_02830_),
    .A(net3897),
    .B(net8151));
 sg13g2_o21ai_1 _23983_ (.B1(_02830_),
    .Y(_00692_),
    .A1(net7583),
    .A2(net8151));
 sg13g2_nand2_1 _23984_ (.Y(_02831_),
    .A(net3176),
    .B(net8149));
 sg13g2_o21ai_1 _23985_ (.B1(_02831_),
    .Y(_00693_),
    .A1(net7563),
    .A2(net8149));
 sg13g2_nand2_1 _23986_ (.Y(_02832_),
    .A(net3368),
    .B(net8148));
 sg13g2_o21ai_1 _23987_ (.B1(_02832_),
    .Y(_00694_),
    .A1(net7522),
    .A2(net8148));
 sg13g2_nand2_1 _23988_ (.Y(_02833_),
    .A(net3286),
    .B(net8148));
 sg13g2_o21ai_1 _23989_ (.B1(_02833_),
    .Y(_00695_),
    .A1(net7534),
    .A2(net8148));
 sg13g2_nand2_1 _23990_ (.Y(_02834_),
    .A(net2909),
    .B(net8149));
 sg13g2_o21ai_1 _23991_ (.B1(_02834_),
    .Y(_00696_),
    .A1(net7529),
    .A2(net8149));
 sg13g2_nand2_1 _23992_ (.Y(_02835_),
    .A(net3034),
    .B(net8159));
 sg13g2_o21ai_1 _23993_ (.B1(_02835_),
    .Y(_00697_),
    .A1(net7520),
    .A2(net8151));
 sg13g2_nand2_1 _23994_ (.Y(_02836_),
    .A(net2896),
    .B(net8154));
 sg13g2_o21ai_1 _23995_ (.B1(_02836_),
    .Y(_00698_),
    .A1(net7507),
    .A2(net8154));
 sg13g2_nand2_1 _23996_ (.Y(_02837_),
    .A(net3961),
    .B(net8152));
 sg13g2_o21ai_1 _23997_ (.B1(_02837_),
    .Y(_00699_),
    .A1(net7513),
    .A2(net8152));
 sg13g2_nand2_1 _23998_ (.Y(_02838_),
    .A(net3268),
    .B(net8156));
 sg13g2_o21ai_1 _23999_ (.B1(_02838_),
    .Y(_00700_),
    .A1(net7495),
    .A2(net8156));
 sg13g2_nand2_1 _24000_ (.Y(_02839_),
    .A(net3769),
    .B(net8149));
 sg13g2_o21ai_1 _24001_ (.B1(_02839_),
    .Y(_00701_),
    .A1(net7499),
    .A2(net8149));
 sg13g2_nand2_1 _24002_ (.Y(_02840_),
    .A(net3785),
    .B(net8152));
 sg13g2_o21ai_1 _24003_ (.B1(_02840_),
    .Y(_00702_),
    .A1(net7644),
    .A2(net8152));
 sg13g2_nand2_1 _24004_ (.Y(_02841_),
    .A(net3136),
    .B(net8153));
 sg13g2_o21ai_1 _24005_ (.B1(_02841_),
    .Y(_00703_),
    .A1(net7648),
    .A2(net8153));
 sg13g2_nand2_1 _24006_ (.Y(_02842_),
    .A(net3307),
    .B(net8155));
 sg13g2_o21ai_1 _24007_ (.B1(_02842_),
    .Y(_00704_),
    .A1(net7654),
    .A2(net8155));
 sg13g2_nand2_1 _24008_ (.Y(_02843_),
    .A(net3035),
    .B(net8151));
 sg13g2_o21ai_1 _24009_ (.B1(_02843_),
    .Y(_00705_),
    .A1(net7658),
    .A2(net8151));
 sg13g2_nand2_1 _24010_ (.Y(_02844_),
    .A(net3929),
    .B(net8152));
 sg13g2_o21ai_1 _24011_ (.B1(_02844_),
    .Y(_00706_),
    .A1(net7640),
    .A2(net8152));
 sg13g2_nand2_1 _24012_ (.Y(_02845_),
    .A(net3029),
    .B(net8153));
 sg13g2_o21ai_1 _24013_ (.B1(_02845_),
    .Y(_00707_),
    .A1(net7625),
    .A2(net8153));
 sg13g2_nand2_1 _24014_ (.Y(_02846_),
    .A(net2877),
    .B(net8151));
 sg13g2_o21ai_1 _24015_ (.B1(_02846_),
    .Y(_00708_),
    .A1(net7622),
    .A2(net8151));
 sg13g2_nand2_1 _24016_ (.Y(_02847_),
    .A(net3836),
    .B(net8150));
 sg13g2_o21ai_1 _24017_ (.B1(_02847_),
    .Y(_00709_),
    .A1(net7631),
    .A2(net8150));
 sg13g2_nor2_1 _24018_ (.A(_10466_),
    .B(_00185_),
    .Y(_02848_));
 sg13g2_nand3_1 _24019_ (.B(_14302_),
    .C(_02848_),
    .A(net9710),
    .Y(_02849_));
 sg13g2_nand2_1 _24020_ (.Y(_02850_),
    .A(net3212),
    .B(net8145));
 sg13g2_o21ai_1 _24021_ (.B1(_02850_),
    .Y(_00710_),
    .A1(net7485),
    .A2(net8145));
 sg13g2_nand2_1 _24022_ (.Y(_02851_),
    .A(net2915),
    .B(net8144));
 sg13g2_o21ai_1 _24023_ (.B1(_02851_),
    .Y(_00711_),
    .A1(net7666),
    .A2(net8144));
 sg13g2_nand2_1 _24024_ (.Y(_02852_),
    .A(net3476),
    .B(net8144));
 sg13g2_o21ai_1 _24025_ (.B1(_02852_),
    .Y(_00712_),
    .A1(net7615),
    .A2(net8144));
 sg13g2_nand2_1 _24026_ (.Y(_02853_),
    .A(net3530),
    .B(net8143));
 sg13g2_o21ai_1 _24027_ (.B1(_02853_),
    .Y(_00713_),
    .A1(net7608),
    .A2(net8143));
 sg13g2_nand2_1 _24028_ (.Y(_02854_),
    .A(net2959),
    .B(net8142));
 sg13g2_o21ai_1 _24029_ (.B1(_02854_),
    .Y(_00714_),
    .A1(net7590),
    .A2(net8142));
 sg13g2_nand2_1 _24030_ (.Y(_02855_),
    .A(net3065),
    .B(net8142));
 sg13g2_o21ai_1 _24031_ (.B1(_02855_),
    .Y(_00715_),
    .A1(net7599),
    .A2(net8142));
 sg13g2_nand2_1 _24032_ (.Y(_02856_),
    .A(net3312),
    .B(net8143));
 sg13g2_o21ai_1 _24033_ (.B1(_02856_),
    .Y(_00716_),
    .A1(net7592),
    .A2(net8143));
 sg13g2_nand2_1 _24034_ (.Y(_02857_),
    .A(net3644),
    .B(net8139));
 sg13g2_o21ai_1 _24035_ (.B1(_02857_),
    .Y(_00717_),
    .A1(net7604),
    .A2(net8139));
 sg13g2_nand2_1 _24036_ (.Y(_02858_),
    .A(net3543),
    .B(net8147));
 sg13g2_o21ai_1 _24037_ (.B1(_02858_),
    .Y(_00718_),
    .A1(net7560),
    .A2(net8147));
 sg13g2_nand2_1 _24038_ (.Y(_02859_),
    .A(net3282),
    .B(net8144));
 sg13g2_o21ai_1 _24039_ (.B1(_02859_),
    .Y(_00719_),
    .A1(net7578),
    .A2(net8144));
 sg13g2_nand2_1 _24040_ (.Y(_02860_),
    .A(net3542),
    .B(net8146));
 sg13g2_o21ai_1 _24041_ (.B1(_02860_),
    .Y(_00720_),
    .A1(net7549),
    .A2(net8146));
 sg13g2_nand2_1 _24042_ (.Y(_02861_),
    .A(net3001),
    .B(net8137));
 sg13g2_o21ai_1 _24043_ (.B1(_02861_),
    .Y(_00721_),
    .A1(net7573),
    .A2(net8137));
 sg13g2_nand2_1 _24044_ (.Y(_02862_),
    .A(net3638),
    .B(net8145));
 sg13g2_o21ai_1 _24045_ (.B1(_02862_),
    .Y(_00722_),
    .A1(net7540),
    .A2(net8145));
 sg13g2_nand2_1 _24046_ (.Y(_02863_),
    .A(net2843),
    .B(net8144));
 sg13g2_o21ai_1 _24047_ (.B1(_02863_),
    .Y(_00723_),
    .A1(net7554),
    .A2(net8144));
 sg13g2_nand2_1 _24048_ (.Y(_02864_),
    .A(net4048),
    .B(net8140));
 sg13g2_o21ai_1 _24049_ (.B1(_02864_),
    .Y(_00724_),
    .A1(net7581),
    .A2(net8140));
 sg13g2_nand2_1 _24050_ (.Y(_02865_),
    .A(net3903),
    .B(net8138));
 sg13g2_o21ai_1 _24051_ (.B1(_02865_),
    .Y(_00725_),
    .A1(net7567),
    .A2(net8138));
 sg13g2_nand2_1 _24052_ (.Y(_02866_),
    .A(net3496),
    .B(net8137));
 sg13g2_o21ai_1 _24053_ (.B1(_02866_),
    .Y(_00726_),
    .A1(net7526),
    .A2(net8137));
 sg13g2_nand2_1 _24054_ (.Y(_02867_),
    .A(net2826),
    .B(net8137));
 sg13g2_o21ai_1 _24055_ (.B1(_02867_),
    .Y(_00727_),
    .A1(net7539),
    .A2(net8137));
 sg13g2_nand2_1 _24056_ (.Y(_02868_),
    .A(net4852),
    .B(net8137));
 sg13g2_o21ai_1 _24057_ (.B1(_02868_),
    .Y(_00728_),
    .A1(net7530),
    .A2(net8137));
 sg13g2_nand2_1 _24058_ (.Y(_02869_),
    .A(net3415),
    .B(net8140));
 sg13g2_o21ai_1 _24059_ (.B1(_02869_),
    .Y(_00729_),
    .A1(net7516),
    .A2(net8139));
 sg13g2_nand2_1 _24060_ (.Y(_02870_),
    .A(net2875),
    .B(net8145));
 sg13g2_o21ai_1 _24061_ (.B1(_02870_),
    .Y(_00730_),
    .A1(net7508),
    .A2(net8145));
 sg13g2_nand2_1 _24062_ (.Y(_02871_),
    .A(net3547),
    .B(net8141));
 sg13g2_o21ai_1 _24063_ (.B1(_02871_),
    .Y(_00731_),
    .A1(net7511),
    .A2(net8141));
 sg13g2_nand2_1 _24064_ (.Y(_02872_),
    .A(net3113),
    .B(net8143));
 sg13g2_o21ai_1 _24065_ (.B1(_02872_),
    .Y(_00732_),
    .A1(net7497),
    .A2(net8143));
 sg13g2_nand2_1 _24066_ (.Y(_02873_),
    .A(net3864),
    .B(net8138));
 sg13g2_o21ai_1 _24067_ (.B1(_02873_),
    .Y(_00733_),
    .A1(net7501),
    .A2(net8138));
 sg13g2_nand2_1 _24068_ (.Y(_02874_),
    .A(net3846),
    .B(net8142));
 sg13g2_o21ai_1 _24069_ (.B1(_02874_),
    .Y(_00734_),
    .A1(net7642),
    .A2(net8142));
 sg13g2_nand2_1 _24070_ (.Y(_02875_),
    .A(net2848),
    .B(net8145));
 sg13g2_o21ai_1 _24071_ (.B1(_02875_),
    .Y(_00735_),
    .A1(net7651),
    .A2(net8145));
 sg13g2_nand2_1 _24072_ (.Y(_02876_),
    .A(net2892),
    .B(net8143));
 sg13g2_o21ai_1 _24073_ (.B1(_02876_),
    .Y(_00736_),
    .A1(net7653),
    .A2(net8143));
 sg13g2_nand2_1 _24074_ (.Y(_02877_),
    .A(net3526),
    .B(net8141));
 sg13g2_o21ai_1 _24075_ (.B1(_02877_),
    .Y(_00737_),
    .A1(net7659),
    .A2(net8141));
 sg13g2_nand2_1 _24076_ (.Y(_02878_),
    .A(net3574),
    .B(net8141));
 sg13g2_o21ai_1 _24077_ (.B1(_02878_),
    .Y(_00738_),
    .A1(net7637),
    .A2(net8141));
 sg13g2_nand2_1 _24078_ (.Y(_02879_),
    .A(net3330),
    .B(net8142));
 sg13g2_o21ai_1 _24079_ (.B1(_02879_),
    .Y(_00739_),
    .A1(net7627),
    .A2(net8142));
 sg13g2_nand2_1 _24080_ (.Y(_02880_),
    .A(net3994),
    .B(net8141));
 sg13g2_o21ai_1 _24081_ (.B1(_02880_),
    .Y(_00740_),
    .A1(net7619),
    .A2(net8140));
 sg13g2_nand2_1 _24082_ (.Y(_02881_),
    .A(net3916),
    .B(net8139));
 sg13g2_o21ai_1 _24083_ (.B1(_02881_),
    .Y(_00741_),
    .A1(net7635),
    .A2(net8139));
 sg13g2_mux4_1 _24084_ (.S0(net9679),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][0] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][0] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][0] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][0] ),
    .S1(net9624),
    .X(_02882_));
 sg13g2_nor2_1 _24085_ (.A(net9576),
    .B(_02882_),
    .Y(_02883_));
 sg13g2_mux4_1 _24086_ (.S0(net9679),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][0] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][0] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][0] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][0] ),
    .S1(net9624),
    .X(_02884_));
 sg13g2_o21ai_1 _24087_ (.B1(net9562),
    .Y(_02885_),
    .A1(net9109),
    .A2(_02884_));
 sg13g2_nor2_1 _24088_ (.A(_02883_),
    .B(_02885_),
    .Y(_02886_));
 sg13g2_nor2b_1 _24089_ (.A(net9677),
    .B_N(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][0] ),
    .Y(_02887_));
 sg13g2_a21oi_1 _24090_ (.A1(net9676),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][0] ),
    .Y(_02888_),
    .B1(_02887_));
 sg13g2_nor2_1 _24091_ (.A(net9557),
    .B(net9108),
    .Y(_02889_));
 sg13g2_mux2_1 _24092_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][0] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][0] ),
    .S(net9678),
    .X(_02890_));
 sg13g2_o21ai_1 _24093_ (.B1(net8814),
    .Y(_02891_),
    .A1(net9621),
    .A2(_02890_));
 sg13g2_a21oi_1 _24094_ (.A1(net9621),
    .A2(_02888_),
    .Y(_02892_),
    .B1(_02891_));
 sg13g2_nor2_2 _24095_ (.A(net9559),
    .B(net9575),
    .Y(_02893_));
 sg13g2_nand2_2 _24096_ (.Y(_02894_),
    .A(_10462_),
    .B(net9108));
 sg13g2_nor2_2 _24097_ (.A(net9613),
    .B(_02894_),
    .Y(_02895_));
 sg13g2_nand2_1 _24098_ (.Y(_02896_),
    .A(net9099),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][0] ));
 sg13g2_nor2b_1 _24099_ (.A(net9679),
    .B_N(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][0] ),
    .Y(_02897_));
 sg13g2_a21oi_1 _24100_ (.A1(net9679),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][0] ),
    .Y(_02898_),
    .B1(_02897_));
 sg13g2_and2_2 _24101_ (.A(net9599),
    .B(net8948),
    .X(_02899_));
 sg13g2_a21oi_1 _24102_ (.A1(net9679),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][0] ),
    .Y(_02900_),
    .B1(net9620));
 sg13g2_a221oi_1 _24103_ (.B2(_02896_),
    .C1(_02894_),
    .B1(_02900_),
    .A1(net9620),
    .Y(_02901_),
    .A2(_02898_));
 sg13g2_nor4_2 _24104_ (.A(net9551),
    .B(_02886_),
    .C(_02892_),
    .Y(_02902_),
    .D(_02901_));
 sg13g2_nor2_2 _24105_ (.A(net9548),
    .B(net9665),
    .Y(_02903_));
 sg13g2_and2_2 _24106_ (.A(_02895_),
    .B(_02903_),
    .X(_02904_));
 sg13g2_nand2_1 _24107_ (.Y(_02905_),
    .A(_02895_),
    .B(_02903_));
 sg13g2_mux4_1 _24108_ (.S0(net9676),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][0] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][0] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][0] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][0] ),
    .S1(net9620),
    .X(_02906_));
 sg13g2_nor2_1 _24109_ (.A(net9575),
    .B(_02906_),
    .Y(_02907_));
 sg13g2_mux4_1 _24110_ (.S0(net9676),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][0] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][0] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][0] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][0] ),
    .S1(net9620),
    .X(_02908_));
 sg13g2_o21ai_1 _24111_ (.B1(net9559),
    .Y(_02909_),
    .A1(net9109),
    .A2(_02908_));
 sg13g2_nor2_1 _24112_ (.A(_02907_),
    .B(_02909_),
    .Y(_02910_));
 sg13g2_nor2_1 _24113_ (.A(net9096),
    .B(_10697_),
    .Y(_02911_));
 sg13g2_a21oi_1 _24114_ (.A1(net9096),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][0] ),
    .Y(_02912_),
    .B1(_02911_));
 sg13g2_mux2_1 _24115_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][0] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][0] ),
    .S(net9676),
    .X(_02913_));
 sg13g2_o21ai_1 _24116_ (.B1(net8814),
    .Y(_02914_),
    .A1(net9620),
    .A2(_02913_));
 sg13g2_a21oi_1 _24117_ (.A1(net9620),
    .A2(_02912_),
    .Y(_02915_),
    .B1(_02914_));
 sg13g2_nand2_1 _24118_ (.Y(_02916_),
    .A(net9099),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][0] ));
 sg13g2_nor2b_1 _24119_ (.A(net9676),
    .B_N(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][0] ),
    .Y(_02917_));
 sg13g2_a21oi_1 _24120_ (.A1(net9676),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][0] ),
    .Y(_02918_),
    .B1(_02917_));
 sg13g2_a21oi_1 _24121_ (.A1(net9676),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][0] ),
    .Y(_02919_),
    .B1(net9620));
 sg13g2_a221oi_1 _24122_ (.B2(_02916_),
    .C1(_02894_),
    .B1(_02919_),
    .A1(net9620),
    .Y(_02920_),
    .A2(_02918_));
 sg13g2_nor3_2 _24123_ (.A(_02910_),
    .B(_02915_),
    .C(_02920_),
    .Y(_02921_));
 sg13g2_a221oi_1 _24124_ (.B2(net9548),
    .C1(_02902_),
    .B1(_02921_),
    .A1(_02895_),
    .Y(_00742_),
    .A2(_02903_));
 sg13g2_nor2_1 _24125_ (.A(net9099),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][1] ),
    .Y(_02922_));
 sg13g2_nor2_1 _24126_ (.A(net9682),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][1] ),
    .Y(_02923_));
 sg13g2_nor3_1 _24127_ (.A(net9626),
    .B(_02922_),
    .C(_02923_),
    .Y(_02924_));
 sg13g2_nor2_1 _24128_ (.A(net9682),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][1] ),
    .Y(_02925_));
 sg13g2_o21ai_1 _24129_ (.B1(net9626),
    .Y(_02926_),
    .A1(net9099),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][1] ));
 sg13g2_o21ai_1 _24130_ (.B1(net9576),
    .Y(_02927_),
    .A1(_02925_),
    .A2(_02926_));
 sg13g2_mux4_1 _24131_ (.S0(net9682),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][1] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][1] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][1] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][1] ),
    .S1(net9627),
    .X(_02928_));
 sg13g2_nor2_1 _24132_ (.A(net9575),
    .B(_02928_),
    .Y(_02929_));
 sg13g2_o21ai_1 _24133_ (.B1(net9559),
    .Y(_02930_),
    .A1(_02924_),
    .A2(_02927_));
 sg13g2_mux4_1 _24134_ (.S0(net9681),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][1] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][1] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][1] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][1] ),
    .S1(net9625),
    .X(_02931_));
 sg13g2_mux4_1 _24135_ (.S0(net9681),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][1] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][1] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][1] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][1] ),
    .S1(net9625),
    .X(_02932_));
 sg13g2_a221oi_1 _24136_ (.B2(net8814),
    .C1(net9551),
    .B1(_02932_),
    .A1(net8954),
    .Y(_02933_),
    .A2(_02931_));
 sg13g2_o21ai_1 _24137_ (.B1(_02933_),
    .Y(_02934_),
    .A1(_02929_),
    .A2(_02930_));
 sg13g2_a21oi_1 _24138_ (.A1(net9106),
    .A2(_10701_),
    .Y(_02935_),
    .B1(net9626));
 sg13g2_o21ai_1 _24139_ (.B1(_02935_),
    .Y(_02936_),
    .A1(net9102),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][1] ));
 sg13g2_nor2_1 _24140_ (.A(net9106),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][1] ),
    .Y(_02937_));
 sg13g2_a21oi_1 _24141_ (.A1(net9102),
    .A2(_10702_),
    .Y(_02938_),
    .B1(_02937_));
 sg13g2_a21oi_1 _24142_ (.A1(net9626),
    .A2(_02938_),
    .Y(_02939_),
    .B1(net9109));
 sg13g2_mux4_1 _24143_ (.S0(net9682),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][1] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][1] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][1] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][1] ),
    .S1(net9627),
    .X(_02940_));
 sg13g2_o21ai_1 _24144_ (.B1(net9561),
    .Y(_02941_),
    .A1(net9581),
    .A2(_02940_));
 sg13g2_a21o_1 _24145_ (.A2(_02939_),
    .A1(_02936_),
    .B1(_02941_),
    .X(_02942_));
 sg13g2_mux4_1 _24146_ (.S0(net9682),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][1] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][1] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][1] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][1] ),
    .S1(net9626),
    .X(_02943_));
 sg13g2_mux4_1 _24147_ (.S0(net9686),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][1] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][1] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][1] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][1] ),
    .S1(net9631),
    .X(_02944_));
 sg13g2_a221oi_1 _24148_ (.B2(net8814),
    .C1(net9113),
    .B1(_02944_),
    .A1(net8954),
    .Y(_02945_),
    .A2(_02943_));
 sg13g2_nand2_1 _24149_ (.Y(_02946_),
    .A(net8596),
    .B(_02934_));
 sg13g2_a21oi_2 _24150_ (.B1(_02946_),
    .Y(_00743_),
    .A2(_02945_),
    .A1(_02942_));
 sg13g2_nor2_1 _24151_ (.A(net9100),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][2] ),
    .Y(_02947_));
 sg13g2_nor2_1 _24152_ (.A(net9681),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][2] ),
    .Y(_02948_));
 sg13g2_nor3_1 _24153_ (.A(net9625),
    .B(_02947_),
    .C(_02948_),
    .Y(_02949_));
 sg13g2_nor2_1 _24154_ (.A(net9679),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][2] ),
    .Y(_02950_));
 sg13g2_o21ai_1 _24155_ (.B1(net9624),
    .Y(_02951_),
    .A1(net9100),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][2] ));
 sg13g2_o21ai_1 _24156_ (.B1(net9576),
    .Y(_02952_),
    .A1(_02950_),
    .A2(_02951_));
 sg13g2_mux4_1 _24157_ (.S0(net9681),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][2] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][2] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][2] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][2] ),
    .S1(net9625),
    .X(_02953_));
 sg13g2_nor2_1 _24158_ (.A(net9576),
    .B(_02953_),
    .Y(_02954_));
 sg13g2_o21ai_1 _24159_ (.B1(net9559),
    .Y(_02955_),
    .A1(_02949_),
    .A2(_02952_));
 sg13g2_mux4_1 _24160_ (.S0(net9681),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][2] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][2] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][2] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][2] ),
    .S1(net9625),
    .X(_02956_));
 sg13g2_mux4_1 _24161_ (.S0(net9681),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][2] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][2] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][2] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][2] ),
    .S1(net9625),
    .X(_02957_));
 sg13g2_a221oi_1 _24162_ (.B2(net8814),
    .C1(net9551),
    .B1(_02957_),
    .A1(net8954),
    .Y(_02958_),
    .A2(_02956_));
 sg13g2_o21ai_1 _24163_ (.B1(_02958_),
    .Y(_02959_),
    .A1(_02954_),
    .A2(_02955_));
 sg13g2_a21oi_1 _24164_ (.A1(net9100),
    .A2(_10705_),
    .Y(_02960_),
    .B1(net9626));
 sg13g2_o21ai_1 _24165_ (.B1(_02960_),
    .Y(_02961_),
    .A1(net9100),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][2] ));
 sg13g2_nor2_1 _24166_ (.A(net9100),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][2] ),
    .Y(_02962_));
 sg13g2_a21oi_1 _24167_ (.A1(net9100),
    .A2(_10706_),
    .Y(_02963_),
    .B1(_02962_));
 sg13g2_a21oi_1 _24168_ (.A1(net9626),
    .A2(_02963_),
    .Y(_02964_),
    .B1(net9108));
 sg13g2_mux4_1 _24169_ (.S0(net9682),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][2] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][2] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][2] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][2] ),
    .S1(net9626),
    .X(_02965_));
 sg13g2_o21ai_1 _24170_ (.B1(net9559),
    .Y(_02966_),
    .A1(net9576),
    .A2(_02965_));
 sg13g2_a21o_1 _24171_ (.A2(_02964_),
    .A1(_02961_),
    .B1(_02966_),
    .X(_02967_));
 sg13g2_mux4_1 _24172_ (.S0(net9681),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][2] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][2] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][2] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][2] ),
    .S1(net9625),
    .X(_02968_));
 sg13g2_mux4_1 _24173_ (.S0(net9681),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][2] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][2] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][2] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][2] ),
    .S1(net9625),
    .X(_02969_));
 sg13g2_a221oi_1 _24174_ (.B2(net8814),
    .C1(net9113),
    .B1(_02969_),
    .A1(net8954),
    .Y(_02970_),
    .A2(_02968_));
 sg13g2_nand2_1 _24175_ (.Y(_02971_),
    .A(net8596),
    .B(_02959_));
 sg13g2_a21oi_2 _24176_ (.B1(_02971_),
    .Y(_00744_),
    .A2(_02970_),
    .A1(_02967_));
 sg13g2_nor2_1 _24177_ (.A(net9104),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][3] ),
    .Y(_02972_));
 sg13g2_nor2_1 _24178_ (.A(net9691),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][3] ),
    .Y(_02973_));
 sg13g2_nor3_1 _24179_ (.A(net9638),
    .B(_02972_),
    .C(_02973_),
    .Y(_02974_));
 sg13g2_nor2_1 _24180_ (.A(net9691),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][3] ),
    .Y(_02975_));
 sg13g2_o21ai_1 _24181_ (.B1(net9638),
    .Y(_02976_),
    .A1(net9103),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][3] ));
 sg13g2_o21ai_1 _24182_ (.B1(net9579),
    .Y(_02977_),
    .A1(_02975_),
    .A2(_02976_));
 sg13g2_mux4_1 _24183_ (.S0(net9691),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][3] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][3] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][3] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][3] ),
    .S1(net9638),
    .X(_02978_));
 sg13g2_nor2_1 _24184_ (.A(net9579),
    .B(_02978_),
    .Y(_02979_));
 sg13g2_o21ai_1 _24185_ (.B1(net9560),
    .Y(_02980_),
    .A1(_02974_),
    .A2(_02977_));
 sg13g2_mux4_1 _24186_ (.S0(net9693),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][3] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][3] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][3] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][3] ),
    .S1(net9637),
    .X(_02981_));
 sg13g2_mux4_1 _24187_ (.S0(net9693),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][3] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][3] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][3] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][3] ),
    .S1(net9637),
    .X(_02982_));
 sg13g2_a221oi_1 _24188_ (.B2(net8815),
    .C1(net9550),
    .B1(_02982_),
    .A1(net8953),
    .Y(_02983_),
    .A2(_02981_));
 sg13g2_o21ai_1 _24189_ (.B1(_02983_),
    .Y(_02984_),
    .A1(_02979_),
    .A2(_02980_));
 sg13g2_nor2_1 _24190_ (.A(net9102),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][3] ),
    .Y(_02985_));
 sg13g2_nor2_1 _24191_ (.A(net9687),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][3] ),
    .Y(_02986_));
 sg13g2_nor3_1 _24192_ (.A(net9632),
    .B(_02985_),
    .C(_02986_),
    .Y(_02987_));
 sg13g2_nor2_1 _24193_ (.A(net9686),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][3] ),
    .Y(_02988_));
 sg13g2_o21ai_1 _24194_ (.B1(net9631),
    .Y(_02989_),
    .A1(net9102),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][3] ));
 sg13g2_o21ai_1 _24195_ (.B1(net9577),
    .Y(_02990_),
    .A1(_02988_),
    .A2(_02989_));
 sg13g2_mux4_1 _24196_ (.S0(net9686),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][3] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][3] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][3] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][3] ),
    .S1(net9631),
    .X(_02991_));
 sg13g2_nor2_1 _24197_ (.A(net9581),
    .B(_02991_),
    .Y(_02992_));
 sg13g2_o21ai_1 _24198_ (.B1(net9561),
    .Y(_02993_),
    .A1(_02987_),
    .A2(_02990_));
 sg13g2_mux4_1 _24199_ (.S0(net9686),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][3] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][3] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][3] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][3] ),
    .S1(net9630),
    .X(_02994_));
 sg13g2_mux4_1 _24200_ (.S0(net9687),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][3] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][3] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][3] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][3] ),
    .S1(net9630),
    .X(_02995_));
 sg13g2_a22oi_1 _24201_ (.Y(_02996_),
    .B1(_02995_),
    .B2(net8953),
    .A2(_02994_),
    .A1(net8815));
 sg13g2_o21ai_1 _24202_ (.B1(_02996_),
    .Y(_02997_),
    .A1(_02992_),
    .A2(_02993_));
 sg13g2_o21ai_1 _24203_ (.B1(_02984_),
    .Y(_02998_),
    .A1(net9113),
    .A2(_02997_));
 sg13g2_nor2_1 _24204_ (.A(net8598),
    .B(_02998_),
    .Y(_00745_));
 sg13g2_nor2_1 _24205_ (.A(net9096),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][4] ),
    .Y(_02999_));
 sg13g2_nor2_1 _24206_ (.A(net9674),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][4] ),
    .Y(_03000_));
 sg13g2_nor3_1 _24207_ (.A(net9616),
    .B(_02999_),
    .C(_03000_),
    .Y(_03001_));
 sg13g2_nor2_1 _24208_ (.A(net9674),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][4] ),
    .Y(_03002_));
 sg13g2_o21ai_1 _24209_ (.B1(net9617),
    .Y(_03003_),
    .A1(net9096),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][4] ));
 sg13g2_o21ai_1 _24210_ (.B1(net9573),
    .Y(_03004_),
    .A1(_03002_),
    .A2(_03003_));
 sg13g2_mux4_1 _24211_ (.S0(net9674),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][4] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][4] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][4] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][4] ),
    .S1(net9617),
    .X(_03005_));
 sg13g2_nor2_1 _24212_ (.A(net9573),
    .B(_03005_),
    .Y(_03006_));
 sg13g2_o21ai_1 _24213_ (.B1(net9557),
    .Y(_03007_),
    .A1(_03001_),
    .A2(_03004_));
 sg13g2_mux4_1 _24214_ (.S0(net9673),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][4] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][4] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][4] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][4] ),
    .S1(net9616),
    .X(_03008_));
 sg13g2_mux4_1 _24215_ (.S0(net9673),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][4] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][4] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][4] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][4] ),
    .S1(net9616),
    .X(_03009_));
 sg13g2_a221oi_1 _24216_ (.B2(net8950),
    .C1(net9549),
    .B1(_03009_),
    .A1(net8813),
    .Y(_03010_),
    .A2(_03008_));
 sg13g2_o21ai_1 _24217_ (.B1(_03010_),
    .Y(_03011_),
    .A1(_03006_),
    .A2(_03007_));
 sg13g2_mux4_1 _24218_ (.S0(net9677),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][4] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][4] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][4] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][4] ),
    .S1(net9619),
    .X(_03012_));
 sg13g2_nor2_1 _24219_ (.A(net9573),
    .B(_03012_),
    .Y(_03013_));
 sg13g2_nor2_1 _24220_ (.A(net9094),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][4] ),
    .Y(_03014_));
 sg13g2_nor2_1 _24221_ (.A(net9674),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][4] ),
    .Y(_03015_));
 sg13g2_nor3_1 _24222_ (.A(net9617),
    .B(_03014_),
    .C(_03015_),
    .Y(_03016_));
 sg13g2_nor2_1 _24223_ (.A(net9674),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][4] ),
    .Y(_03017_));
 sg13g2_o21ai_1 _24224_ (.B1(net9617),
    .Y(_03018_),
    .A1(net9094),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][4] ));
 sg13g2_o21ai_1 _24225_ (.B1(net9573),
    .Y(_03019_),
    .A1(_03017_),
    .A2(_03018_));
 sg13g2_o21ai_1 _24226_ (.B1(net9557),
    .Y(_03020_),
    .A1(_03016_),
    .A2(_03019_));
 sg13g2_mux4_1 _24227_ (.S0(net9673),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][4] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][4] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][4] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][4] ),
    .S1(net9616),
    .X(_03021_));
 sg13g2_mux4_1 _24228_ (.S0(net9673),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][4] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][4] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][4] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][4] ),
    .S1(net9616),
    .X(_03022_));
 sg13g2_a221oi_1 _24229_ (.B2(net8951),
    .C1(net9115),
    .B1(_03022_),
    .A1(net8813),
    .Y(_03023_),
    .A2(_03021_));
 sg13g2_o21ai_1 _24230_ (.B1(_03023_),
    .Y(_03024_),
    .A1(_03013_),
    .A2(_03020_));
 sg13g2_and3_2 _24231_ (.X(_00746_),
    .A(net8595),
    .B(_03011_),
    .C(_03024_));
 sg13g2_mux4_1 _24232_ (.S0(net9667),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][5] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][5] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][5] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][5] ),
    .S1(net9610),
    .X(_03025_));
 sg13g2_nor2_1 _24233_ (.A(net9571),
    .B(_03025_),
    .Y(_03026_));
 sg13g2_nor2_1 _24234_ (.A(net9092),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][5] ),
    .Y(_03027_));
 sg13g2_nor2_1 _24235_ (.A(net9668),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][5] ),
    .Y(_03028_));
 sg13g2_nor3_1 _24236_ (.A(net9608),
    .B(_03027_),
    .C(_03028_),
    .Y(_03029_));
 sg13g2_nor2_1 _24237_ (.A(net9668),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][5] ),
    .Y(_03030_));
 sg13g2_o21ai_1 _24238_ (.B1(net9611),
    .Y(_03031_),
    .A1(net9095),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][5] ));
 sg13g2_o21ai_1 _24239_ (.B1(net9571),
    .Y(_03032_),
    .A1(_03030_),
    .A2(_03031_));
 sg13g2_o21ai_1 _24240_ (.B1(net9557),
    .Y(_03033_),
    .A1(_03029_),
    .A2(_03032_));
 sg13g2_mux4_1 _24241_ (.S0(net9669),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][5] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][5] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][5] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][5] ),
    .S1(net9612),
    .X(_03034_));
 sg13g2_mux4_1 _24242_ (.S0(net9669),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][5] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][5] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][5] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][5] ),
    .S1(net9612),
    .X(_03035_));
 sg13g2_a221oi_1 _24243_ (.B2(net8950),
    .C1(net9548),
    .B1(_03035_),
    .A1(net8812),
    .Y(_03036_),
    .A2(_03034_));
 sg13g2_o21ai_1 _24244_ (.B1(_03036_),
    .Y(_03037_),
    .A1(_03026_),
    .A2(_03033_));
 sg13g2_nor2_1 _24245_ (.A(net9095),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][5] ),
    .Y(_03038_));
 sg13g2_nor2_1 _24246_ (.A(net9668),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][5] ),
    .Y(_03039_));
 sg13g2_nor3_1 _24247_ (.A(net9610),
    .B(_03038_),
    .C(_03039_),
    .Y(_03040_));
 sg13g2_nor2_1 _24248_ (.A(net9668),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][5] ),
    .Y(_03041_));
 sg13g2_o21ai_1 _24249_ (.B1(net9610),
    .Y(_03042_),
    .A1(net9092),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][5] ));
 sg13g2_o21ai_1 _24250_ (.B1(net9574),
    .Y(_03043_),
    .A1(_03041_),
    .A2(_03042_));
 sg13g2_mux4_1 _24251_ (.S0(net9668),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][5] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][5] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][5] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][5] ),
    .S1(net9611),
    .X(_03044_));
 sg13g2_nor2_1 _24252_ (.A(net9571),
    .B(_03044_),
    .Y(_03045_));
 sg13g2_o21ai_1 _24253_ (.B1(net9557),
    .Y(_03046_),
    .A1(_03040_),
    .A2(_03043_));
 sg13g2_a22oi_1 _24254_ (.Y(_03047_),
    .B1(_02899_),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][5] ),
    .A2(net8674),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][5] ));
 sg13g2_o21ai_1 _24255_ (.B1(net9548),
    .Y(_03048_),
    .A1(net9667),
    .A2(_03047_));
 sg13g2_mux4_1 _24256_ (.S0(net9667),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][5] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][5] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][5] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][5] ),
    .S1(net9610),
    .X(_03049_));
 sg13g2_a22oi_1 _24257_ (.Y(_03050_),
    .B1(_02899_),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][5] ),
    .A2(net8674),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][5] ));
 sg13g2_inv_1 _24258_ (.Y(_03051_),
    .A(_03050_));
 sg13g2_a221oi_1 _24259_ (.B2(net9667),
    .C1(_03048_),
    .B1(_03051_),
    .A1(net8812),
    .Y(_03052_),
    .A2(_03049_));
 sg13g2_o21ai_1 _24260_ (.B1(_03052_),
    .Y(_03053_),
    .A1(_03045_),
    .A2(_03046_));
 sg13g2_and3_1 _24261_ (.X(_00747_),
    .A(net8595),
    .B(_03037_),
    .C(_03053_));
 sg13g2_nor2_1 _24262_ (.A(net9105),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][6] ),
    .Y(_03054_));
 sg13g2_nor2_1 _24263_ (.A(net9688),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][6] ),
    .Y(_03055_));
 sg13g2_nor3_1 _24264_ (.A(net9634),
    .B(_03054_),
    .C(_03055_),
    .Y(_03056_));
 sg13g2_nor2_1 _24265_ (.A(net9688),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][6] ),
    .Y(_03057_));
 sg13g2_o21ai_1 _24266_ (.B1(net9634),
    .Y(_03058_),
    .A1(net9105),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][6] ));
 sg13g2_o21ai_1 _24267_ (.B1(net9580),
    .Y(_03059_),
    .A1(_03057_),
    .A2(_03058_));
 sg13g2_mux4_1 _24268_ (.S0(net9690),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][6] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][6] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][6] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][6] ),
    .S1(net9633),
    .X(_03060_));
 sg13g2_nor2_1 _24269_ (.A(net9580),
    .B(_03060_),
    .Y(_03061_));
 sg13g2_o21ai_1 _24270_ (.B1(net9560),
    .Y(_03062_),
    .A1(_03056_),
    .A2(_03059_));
 sg13g2_mux4_1 _24271_ (.S0(net9688),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][6] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][6] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][6] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][6] ),
    .S1(net9634),
    .X(_03063_));
 sg13g2_mux4_1 _24272_ (.S0(net9688),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][6] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][6] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][6] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][6] ),
    .S1(net9634),
    .X(_03064_));
 sg13g2_a221oi_1 _24273_ (.B2(net8952),
    .C1(net9551),
    .B1(_03064_),
    .A1(net8816),
    .Y(_03065_),
    .A2(_03063_));
 sg13g2_o21ai_1 _24274_ (.B1(_03065_),
    .Y(_03066_),
    .A1(_03061_),
    .A2(_03062_));
 sg13g2_nor2_1 _24275_ (.A(net9105),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][6] ),
    .Y(_03067_));
 sg13g2_nor2_1 _24276_ (.A(net9690),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][6] ),
    .Y(_03068_));
 sg13g2_nor3_1 _24277_ (.A(net9633),
    .B(_03067_),
    .C(_03068_),
    .Y(_03069_));
 sg13g2_nor2_1 _24278_ (.A(net9690),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][6] ),
    .Y(_03070_));
 sg13g2_o21ai_1 _24279_ (.B1(net9633),
    .Y(_03071_),
    .A1(net9105),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][6] ));
 sg13g2_o21ai_1 _24280_ (.B1(net9580),
    .Y(_03072_),
    .A1(_03070_),
    .A2(_03071_));
 sg13g2_mux4_1 _24281_ (.S0(net9684),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][6] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][6] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][6] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][6] ),
    .S1(net9628),
    .X(_03073_));
 sg13g2_nor2_1 _24282_ (.A(net9580),
    .B(_03073_),
    .Y(_03074_));
 sg13g2_o21ai_1 _24283_ (.B1(net9560),
    .Y(_03075_),
    .A1(_03069_),
    .A2(_03072_));
 sg13g2_mux4_1 _24284_ (.S0(net9684),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][6] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][6] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][6] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][6] ),
    .S1(net9629),
    .X(_03076_));
 sg13g2_mux4_1 _24285_ (.S0(net9690),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][6] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][6] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][6] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][6] ),
    .S1(net9633),
    .X(_03077_));
 sg13g2_a22oi_1 _24286_ (.Y(_03078_),
    .B1(_03077_),
    .B2(net8952),
    .A2(_03076_),
    .A1(net8816));
 sg13g2_o21ai_1 _24287_ (.B1(_03078_),
    .Y(_03079_),
    .A1(_03074_),
    .A2(_03075_));
 sg13g2_o21ai_1 _24288_ (.B1(_03066_),
    .Y(_03080_),
    .A1(net9113),
    .A2(_03079_));
 sg13g2_nor2_1 _24289_ (.A(net8598),
    .B(_03080_),
    .Y(_00748_));
 sg13g2_nor2_1 _24290_ (.A(net9079),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][7] ),
    .Y(_03081_));
 sg13g2_nor2_1 _24291_ (.A(net9644),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][7] ),
    .Y(_03082_));
 sg13g2_nor3_1 _24292_ (.A(net9585),
    .B(_03081_),
    .C(_03082_),
    .Y(_03083_));
 sg13g2_nor2_1 _24293_ (.A(net9644),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][7] ),
    .Y(_03084_));
 sg13g2_o21ai_1 _24294_ (.B1(net9585),
    .Y(_03085_),
    .A1(net9079),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][7] ));
 sg13g2_o21ai_1 _24295_ (.B1(net9564),
    .Y(_03086_),
    .A1(_03084_),
    .A2(_03085_));
 sg13g2_mux4_1 _24296_ (.S0(net9642),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][7] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][7] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][7] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][7] ),
    .S1(net9583),
    .X(_03087_));
 sg13g2_nor2_1 _24297_ (.A(net9564),
    .B(_03087_),
    .Y(_03088_));
 sg13g2_o21ai_1 _24298_ (.B1(net9553),
    .Y(_03089_),
    .A1(_03083_),
    .A2(_03086_));
 sg13g2_mux4_1 _24299_ (.S0(net9642),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][7] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][7] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][7] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][7] ),
    .S1(net9583),
    .X(_03090_));
 sg13g2_mux4_1 _24300_ (.S0(net9642),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][7] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][7] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][7] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][7] ),
    .S1(net9583),
    .X(_03091_));
 sg13g2_a221oi_1 _24301_ (.B2(net8808),
    .C1(net9546),
    .B1(_03091_),
    .A1(net8946),
    .Y(_03092_),
    .A2(_03090_));
 sg13g2_o21ai_1 _24302_ (.B1(_03092_),
    .Y(_03093_),
    .A1(_03088_),
    .A2(_03089_));
 sg13g2_a21oi_1 _24303_ (.A1(net9082),
    .A2(_10720_),
    .Y(_03094_),
    .B1(net9594));
 sg13g2_o21ai_1 _24304_ (.B1(_03094_),
    .Y(_03095_),
    .A1(net9082),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][7] ));
 sg13g2_o21ai_1 _24305_ (.B1(net9595),
    .Y(_03096_),
    .A1(net9653),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][7] ));
 sg13g2_a21oi_1 _24306_ (.A1(net9653),
    .A2(_10721_),
    .Y(_03097_),
    .B1(_03096_));
 sg13g2_nor2_1 _24307_ (.A(net9110),
    .B(_03097_),
    .Y(_03098_));
 sg13g2_mux4_1 _24308_ (.S0(net9654),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][7] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][7] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][7] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][7] ),
    .S1(net9594),
    .X(_03099_));
 sg13g2_o21ai_1 _24309_ (.B1(net9556),
    .Y(_03100_),
    .A1(net9567),
    .A2(_03099_));
 sg13g2_a21o_1 _24310_ (.A2(_03098_),
    .A1(_03095_),
    .B1(_03100_),
    .X(_03101_));
 sg13g2_mux4_1 _24311_ (.S0(net9651),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][7] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][7] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][7] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][7] ),
    .S1(net9592),
    .X(_03102_));
 sg13g2_mux4_1 _24312_ (.S0(net9651),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][7] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][7] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][7] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][7] ),
    .S1(net9592),
    .X(_03103_));
 sg13g2_a221oi_1 _24313_ (.B2(net8809),
    .C1(net9111),
    .B1(_03103_),
    .A1(net8946),
    .Y(_03104_),
    .A2(_03102_));
 sg13g2_nand2_1 _24314_ (.Y(_03105_),
    .A(net8594),
    .B(_03093_));
 sg13g2_a21oi_2 _24315_ (.B1(_03105_),
    .Y(_00749_),
    .A2(_03104_),
    .A1(_03101_));
 sg13g2_a21oi_1 _24316_ (.A1(net9093),
    .A2(_10723_),
    .Y(_03106_),
    .B1(net9614));
 sg13g2_o21ai_1 _24317_ (.B1(_03106_),
    .Y(_03107_),
    .A1(net9093),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][8] ));
 sg13g2_o21ai_1 _24318_ (.B1(net9614),
    .Y(_03108_),
    .A1(net9671),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][8] ));
 sg13g2_a21oi_1 _24319_ (.A1(net9671),
    .A2(_10724_),
    .Y(_03109_),
    .B1(_03108_));
 sg13g2_nor2_1 _24320_ (.A(net9108),
    .B(_03109_),
    .Y(_03110_));
 sg13g2_mux4_1 _24321_ (.S0(net9670),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][8] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][8] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][8] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][8] ),
    .S1(net9613),
    .X(_03111_));
 sg13g2_o21ai_1 _24322_ (.B1(net9558),
    .Y(_03112_),
    .A1(net9572),
    .A2(_03111_));
 sg13g2_a21o_1 _24323_ (.A2(_03110_),
    .A1(_03107_),
    .B1(_03112_),
    .X(_03113_));
 sg13g2_mux4_1 _24324_ (.S0(net9670),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][8] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][8] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][8] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][8] ),
    .S1(net9613),
    .X(_03114_));
 sg13g2_mux4_1 _24325_ (.S0(net9670),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][8] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][8] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][8] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][8] ),
    .S1(net9613),
    .X(_03115_));
 sg13g2_a221oi_1 _24326_ (.B2(net8812),
    .C1(net9548),
    .B1(_03115_),
    .A1(net8950),
    .Y(_03116_),
    .A2(_03114_));
 sg13g2_a21oi_1 _24327_ (.A1(net9093),
    .A2(_10726_),
    .Y(_03117_),
    .B1(net9614));
 sg13g2_o21ai_1 _24328_ (.B1(_03117_),
    .Y(_03118_),
    .A1(net9093),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][8] ));
 sg13g2_o21ai_1 _24329_ (.B1(net9614),
    .Y(_03119_),
    .A1(net9671),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][8] ));
 sg13g2_a21oi_1 _24330_ (.A1(net9671),
    .A2(_10727_),
    .Y(_03120_),
    .B1(_03119_));
 sg13g2_nor2_1 _24331_ (.A(net9108),
    .B(_03120_),
    .Y(_03121_));
 sg13g2_mux4_1 _24332_ (.S0(net9671),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][8] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][8] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][8] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][8] ),
    .S1(net9614),
    .X(_03122_));
 sg13g2_o21ai_1 _24333_ (.B1(net9558),
    .Y(_03123_),
    .A1(net9572),
    .A2(_03122_));
 sg13g2_a21oi_1 _24334_ (.A1(_03118_),
    .A2(_03121_),
    .Y(_03124_),
    .B1(_03123_));
 sg13g2_mux4_1 _24335_ (.S0(net9670),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][8] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][8] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][8] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][8] ),
    .S1(net9613),
    .X(_03125_));
 sg13g2_mux4_1 _24336_ (.S0(net9671),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][8] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][8] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][8] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][8] ),
    .S1(net9614),
    .X(_03126_));
 sg13g2_a221oi_1 _24337_ (.B2(net8813),
    .C1(_03124_),
    .B1(_03126_),
    .A1(net8951),
    .Y(_03127_),
    .A2(_03125_));
 sg13g2_a221oi_1 _24338_ (.B2(net9549),
    .C1(net8598),
    .B1(_03127_),
    .A1(_03113_),
    .Y(_00750_),
    .A2(_03116_));
 sg13g2_mux4_1 _24339_ (.S0(net9685),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][9] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][9] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][9] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][9] ),
    .S1(net9628),
    .X(_03128_));
 sg13g2_nor2_1 _24340_ (.A(net9577),
    .B(_03128_),
    .Y(_03129_));
 sg13g2_nor2_1 _24341_ (.A(net9101),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][9] ),
    .Y(_03130_));
 sg13g2_nor2_1 _24342_ (.A(net9685),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][9] ),
    .Y(_03131_));
 sg13g2_nor3_1 _24343_ (.A(net9628),
    .B(_03130_),
    .C(_03131_),
    .Y(_03132_));
 sg13g2_nor2_1 _24344_ (.A(net9685),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][9] ),
    .Y(_03133_));
 sg13g2_o21ai_1 _24345_ (.B1(net9628),
    .Y(_03134_),
    .A1(net9102),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][9] ));
 sg13g2_o21ai_1 _24346_ (.B1(net9577),
    .Y(_03135_),
    .A1(_03133_),
    .A2(_03134_));
 sg13g2_o21ai_1 _24347_ (.B1(net9561),
    .Y(_03136_),
    .A1(_03132_),
    .A2(_03135_));
 sg13g2_mux4_1 _24348_ (.S0(net9686),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][9] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][9] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][9] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][9] ),
    .S1(net9631),
    .X(_03137_));
 sg13g2_mux4_1 _24349_ (.S0(net9687),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][9] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][9] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][9] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][9] ),
    .S1(net9630),
    .X(_03138_));
 sg13g2_a221oi_1 _24350_ (.B2(net8953),
    .C1(net9550),
    .B1(_03138_),
    .A1(net8815),
    .Y(_03139_),
    .A2(_03137_));
 sg13g2_o21ai_1 _24351_ (.B1(_03139_),
    .Y(_03140_),
    .A1(_03129_),
    .A2(_03136_));
 sg13g2_nand2b_1 _24352_ (.Y(_03141_),
    .B(net9685),
    .A_N(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][9] ));
 sg13g2_a21oi_1 _24353_ (.A1(net9101),
    .A2(_10730_),
    .Y(_03142_),
    .B1(net9628));
 sg13g2_mux2_1 _24354_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][9] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][9] ),
    .S(net9685),
    .X(_03143_));
 sg13g2_a221oi_1 _24355_ (.B2(net9623),
    .C1(net9577),
    .B1(_03143_),
    .A1(_03141_),
    .Y(_03144_),
    .A2(_03142_));
 sg13g2_nor2_1 _24356_ (.A(net9101),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][9] ),
    .Y(_03145_));
 sg13g2_nor2_1 _24357_ (.A(net9680),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][9] ),
    .Y(_03146_));
 sg13g2_nor3_1 _24358_ (.A(net9624),
    .B(_03145_),
    .C(_03146_),
    .Y(_03147_));
 sg13g2_nor2_1 _24359_ (.A(net9679),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][9] ),
    .Y(_03148_));
 sg13g2_o21ai_1 _24360_ (.B1(net9623),
    .Y(_03149_),
    .A1(net9101),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][9] ));
 sg13g2_o21ai_1 _24361_ (.B1(net9577),
    .Y(_03150_),
    .A1(_03148_),
    .A2(_03149_));
 sg13g2_o21ai_1 _24362_ (.B1(net9561),
    .Y(_03151_),
    .A1(_03147_),
    .A2(_03150_));
 sg13g2_mux4_1 _24363_ (.S0(net9686),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][9] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][9] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][9] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][9] ),
    .S1(net9631),
    .X(_03152_));
 sg13g2_mux4_1 _24364_ (.S0(net9686),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][9] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][9] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][9] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][9] ),
    .S1(net9631),
    .X(_03153_));
 sg13g2_a221oi_1 _24365_ (.B2(net8954),
    .C1(net9113),
    .B1(_03153_),
    .A1(net8814),
    .Y(_03154_),
    .A2(_03152_));
 sg13g2_o21ai_1 _24366_ (.B1(_03154_),
    .Y(_03155_),
    .A1(_03144_),
    .A2(_03151_));
 sg13g2_and3_2 _24367_ (.X(_00751_),
    .A(net8596),
    .B(_03140_),
    .C(_03155_));
 sg13g2_mux4_1 _24368_ (.S0(net9688),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][10] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][10] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][10] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][10] ),
    .S1(net9634),
    .X(_03156_));
 sg13g2_nor2_1 _24369_ (.A(net9580),
    .B(_03156_),
    .Y(_03157_));
 sg13g2_nor2_1 _24370_ (.A(net9103),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][10] ),
    .Y(_03158_));
 sg13g2_nor2_1 _24371_ (.A(net9689),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][10] ),
    .Y(_03159_));
 sg13g2_nor3_1 _24372_ (.A(net9636),
    .B(_03158_),
    .C(_03159_),
    .Y(_03160_));
 sg13g2_nor2_1 _24373_ (.A(net9689),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][10] ),
    .Y(_03161_));
 sg13g2_o21ai_1 _24374_ (.B1(net9634),
    .Y(_03162_),
    .A1(net9103),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][10] ));
 sg13g2_o21ai_1 _24375_ (.B1(net9579),
    .Y(_03163_),
    .A1(_03161_),
    .A2(_03162_));
 sg13g2_o21ai_1 _24376_ (.B1(net9560),
    .Y(_03164_),
    .A1(_03160_),
    .A2(_03163_));
 sg13g2_mux4_1 _24377_ (.S0(net9688),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][10] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][10] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][10] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][10] ),
    .S1(net9634),
    .X(_03165_));
 sg13g2_mux4_1 _24378_ (.S0(net9692),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][10] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][10] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][10] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][10] ),
    .S1(net9636),
    .X(_03166_));
 sg13g2_a221oi_1 _24379_ (.B2(net8816),
    .C1(net9550),
    .B1(_03166_),
    .A1(net8952),
    .Y(_03167_),
    .A2(_03165_));
 sg13g2_o21ai_1 _24380_ (.B1(_03167_),
    .Y(_03168_),
    .A1(_03157_),
    .A2(_03164_));
 sg13g2_mux4_1 _24381_ (.S0(net9691),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][10] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][10] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][10] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][10] ),
    .S1(net9638),
    .X(_03169_));
 sg13g2_nor2_1 _24382_ (.A(net9578),
    .B(_03169_),
    .Y(_03170_));
 sg13g2_nor2_1 _24383_ (.A(net9103),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][10] ),
    .Y(_03171_));
 sg13g2_nor2_1 _24384_ (.A(net9690),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][10] ),
    .Y(_03172_));
 sg13g2_nor3_1 _24385_ (.A(net9635),
    .B(_03171_),
    .C(_03172_),
    .Y(_03173_));
 sg13g2_nor2_1 _24386_ (.A(net9690),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][10] ),
    .Y(_03174_));
 sg13g2_o21ai_1 _24387_ (.B1(net9633),
    .Y(_03175_),
    .A1(net9104),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][10] ));
 sg13g2_o21ai_1 _24388_ (.B1(net9578),
    .Y(_03176_),
    .A1(_03174_),
    .A2(_03175_));
 sg13g2_o21ai_1 _24389_ (.B1(net9560),
    .Y(_03177_),
    .A1(_03173_),
    .A2(_03176_));
 sg13g2_mux4_1 _24390_ (.S0(net9690),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][10] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][10] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][10] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][10] ),
    .S1(net9633),
    .X(_03178_));
 sg13g2_mux4_1 _24391_ (.S0(net9685),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][10] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][10] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][10] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][10] ),
    .S1(net9629),
    .X(_03179_));
 sg13g2_a22oi_1 _24392_ (.Y(_03180_),
    .B1(_03179_),
    .B2(net8816),
    .A2(_03178_),
    .A1(net8952));
 sg13g2_o21ai_1 _24393_ (.B1(_03180_),
    .Y(_03181_),
    .A1(_03170_),
    .A2(_03177_));
 sg13g2_o21ai_1 _24394_ (.B1(_03168_),
    .Y(_03182_),
    .A1(net9113),
    .A2(_03181_));
 sg13g2_nor2_2 _24395_ (.A(net8597),
    .B(_03182_),
    .Y(_00752_));
 sg13g2_nor2_1 _24396_ (.A(net9079),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][11] ),
    .Y(_03183_));
 sg13g2_nor2_1 _24397_ (.A(net9644),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][11] ),
    .Y(_03184_));
 sg13g2_nor3_1 _24398_ (.A(net9585),
    .B(_03183_),
    .C(_03184_),
    .Y(_03185_));
 sg13g2_nor2_1 _24399_ (.A(net9644),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][11] ),
    .Y(_03186_));
 sg13g2_o21ai_1 _24400_ (.B1(net9585),
    .Y(_03187_),
    .A1(net9079),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][11] ));
 sg13g2_o21ai_1 _24401_ (.B1(net9564),
    .Y(_03188_),
    .A1(_03186_),
    .A2(_03187_));
 sg13g2_mux4_1 _24402_ (.S0(net9642),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][11] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][11] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][11] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][11] ),
    .S1(net9583),
    .X(_03189_));
 sg13g2_nor2_1 _24403_ (.A(net9564),
    .B(_03189_),
    .Y(_03190_));
 sg13g2_o21ai_1 _24404_ (.B1(net9553),
    .Y(_03191_),
    .A1(_03185_),
    .A2(_03188_));
 sg13g2_mux4_1 _24405_ (.S0(net9642),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][11] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][11] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][11] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][11] ),
    .S1(net9583),
    .X(_03192_));
 sg13g2_mux4_1 _24406_ (.S0(net9642),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][11] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][11] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][11] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][11] ),
    .S1(net9583),
    .X(_03193_));
 sg13g2_a221oi_1 _24407_ (.B2(net8808),
    .C1(net9546),
    .B1(_03193_),
    .A1(net8946),
    .Y(_03194_),
    .A2(_03192_));
 sg13g2_o21ai_1 _24408_ (.B1(_03194_),
    .Y(_03195_),
    .A1(_03190_),
    .A2(_03191_));
 sg13g2_mux4_1 _24409_ (.S0(net9648),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][11] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][11] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][11] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][11] ),
    .S1(net9589),
    .X(_03196_));
 sg13g2_nor2_1 _24410_ (.A(net9081),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][11] ),
    .Y(_03197_));
 sg13g2_nor2_1 _24411_ (.A(net9650),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][11] ),
    .Y(_03198_));
 sg13g2_nor3_1 _24412_ (.A(net9591),
    .B(_03197_),
    .C(_03198_),
    .Y(_03199_));
 sg13g2_nor2_1 _24413_ (.A(net9650),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][11] ),
    .Y(_03200_));
 sg13g2_o21ai_1 _24414_ (.B1(net9591),
    .Y(_03201_),
    .A1(net9081),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][11] ));
 sg13g2_o21ai_1 _24415_ (.B1(net9565),
    .Y(_03202_),
    .A1(_03200_),
    .A2(_03201_));
 sg13g2_o21ai_1 _24416_ (.B1(net9554),
    .Y(_03203_),
    .A1(_03199_),
    .A2(_03202_));
 sg13g2_inv_1 _24417_ (.Y(_03204_),
    .A(_03203_));
 sg13g2_o21ai_1 _24418_ (.B1(_03204_),
    .Y(_03205_),
    .A1(net9565),
    .A2(_03196_));
 sg13g2_mux4_1 _24419_ (.S0(net9648),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][11] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][11] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][11] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][11] ),
    .S1(net9589),
    .X(_03206_));
 sg13g2_mux4_1 _24420_ (.S0(net9647),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][11] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][11] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][11] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][11] ),
    .S1(net9588),
    .X(_03207_));
 sg13g2_a221oi_1 _24421_ (.B2(net8809),
    .C1(net9111),
    .B1(_03207_),
    .A1(net8947),
    .Y(_03208_),
    .A2(_03206_));
 sg13g2_nand2_1 _24422_ (.Y(_03209_),
    .A(net8594),
    .B(_03195_));
 sg13g2_a21oi_2 _24423_ (.B1(_03209_),
    .Y(_00753_),
    .A2(_03208_),
    .A1(_03205_));
 sg13g2_nor2_1 _24424_ (.A(net9105),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][12] ),
    .Y(_03210_));
 sg13g2_nor2_1 _24425_ (.A(net9688),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][12] ),
    .Y(_03211_));
 sg13g2_nor3_1 _24426_ (.A(net9634),
    .B(_03210_),
    .C(_03211_),
    .Y(_03212_));
 sg13g2_nor2_1 _24427_ (.A(net9688),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][12] ),
    .Y(_03213_));
 sg13g2_o21ai_1 _24428_ (.B1(net9633),
    .Y(_03214_),
    .A1(net9105),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][12] ));
 sg13g2_o21ai_1 _24429_ (.B1(net9580),
    .Y(_03215_),
    .A1(_03213_),
    .A2(_03214_));
 sg13g2_mux4_1 _24430_ (.S0(net9690),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][12] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][12] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][12] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][12] ),
    .S1(net9633),
    .X(_03216_));
 sg13g2_nor2_1 _24431_ (.A(net9580),
    .B(_03216_),
    .Y(_03217_));
 sg13g2_o21ai_1 _24432_ (.B1(net9560),
    .Y(_03218_),
    .A1(_03212_),
    .A2(_03215_));
 sg13g2_mux4_1 _24433_ (.S0(net9689),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][12] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][12] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][12] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][12] ),
    .S1(net9635),
    .X(_03219_));
 sg13g2_mux4_1 _24434_ (.S0(net9689),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][12] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][12] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][12] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][12] ),
    .S1(net9635),
    .X(_03220_));
 sg13g2_a221oi_1 _24435_ (.B2(net8816),
    .C1(net9550),
    .B1(_03220_),
    .A1(net8952),
    .Y(_03221_),
    .A2(_03219_));
 sg13g2_o21ai_1 _24436_ (.B1(_03221_),
    .Y(_03222_),
    .A1(_03217_),
    .A2(_03218_));
 sg13g2_a21oi_1 _24437_ (.A1(net9099),
    .A2(_10742_),
    .Y(_03223_),
    .B1(net9623));
 sg13g2_o21ai_1 _24438_ (.B1(_03223_),
    .Y(_03224_),
    .A1(net9099),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][12] ));
 sg13g2_nor2_1 _24439_ (.A(net9099),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][12] ),
    .Y(_03225_));
 sg13g2_a21oi_1 _24440_ (.A1(net9099),
    .A2(_10743_),
    .Y(_03226_),
    .B1(_03225_));
 sg13g2_a21oi_1 _24441_ (.A1(net9623),
    .A2(_03226_),
    .Y(_03227_),
    .B1(net9108));
 sg13g2_mux4_1 _24442_ (.S0(net9679),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][12] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][12] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][12] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][12] ),
    .S1(net9624),
    .X(_03228_));
 sg13g2_o21ai_1 _24443_ (.B1(net9562),
    .Y(_03229_),
    .A1(net9576),
    .A2(_03228_));
 sg13g2_a21o_1 _24444_ (.A2(_03227_),
    .A1(_03224_),
    .B1(_03229_),
    .X(_03230_));
 sg13g2_mux4_1 _24445_ (.S0(net9680),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][12] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][12] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][12] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][12] ),
    .S1(net9623),
    .X(_03231_));
 sg13g2_mux4_1 _24446_ (.S0(net9680),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][12] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][12] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][12] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][12] ),
    .S1(net9623),
    .X(_03232_));
 sg13g2_a221oi_1 _24447_ (.B2(net8817),
    .C1(net9113),
    .B1(_03232_),
    .A1(net8954),
    .Y(_03233_),
    .A2(_03231_));
 sg13g2_nand2_2 _24448_ (.Y(_03234_),
    .A(net8595),
    .B(_03222_));
 sg13g2_a21oi_2 _24449_ (.B1(_03234_),
    .Y(_00754_),
    .A2(_03233_),
    .A1(_03230_));
 sg13g2_nor2_1 _24450_ (.A(net9102),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][13] ),
    .Y(_03235_));
 sg13g2_nor2_1 _24451_ (.A(net9684),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][13] ),
    .Y(_03236_));
 sg13g2_nor3_1 _24452_ (.A(net9629),
    .B(_03235_),
    .C(_03236_),
    .Y(_03237_));
 sg13g2_nor2_1 _24453_ (.A(net9684),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][13] ),
    .Y(_03238_));
 sg13g2_o21ai_1 _24454_ (.B1(net9629),
    .Y(_03239_),
    .A1(net9102),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][13] ));
 sg13g2_o21ai_1 _24455_ (.B1(net9577),
    .Y(_03240_),
    .A1(_03238_),
    .A2(_03239_));
 sg13g2_mux4_1 _24456_ (.S0(net9684),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][13] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][13] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][13] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][13] ),
    .S1(net9629),
    .X(_03241_));
 sg13g2_nor2_1 _24457_ (.A(net9577),
    .B(_03241_),
    .Y(_03242_));
 sg13g2_o21ai_1 _24458_ (.B1(net9561),
    .Y(_03243_),
    .A1(_03237_),
    .A2(_03240_));
 sg13g2_mux4_1 _24459_ (.S0(net9684),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][13] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][13] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][13] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][13] ),
    .S1(net9629),
    .X(_03244_));
 sg13g2_mux4_1 _24460_ (.S0(net9684),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][13] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][13] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][13] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][13] ),
    .S1(net9629),
    .X(_03245_));
 sg13g2_a221oi_1 _24461_ (.B2(net8815),
    .C1(net9550),
    .B1(_03245_),
    .A1(net8953),
    .Y(_03246_),
    .A2(_03244_));
 sg13g2_o21ai_1 _24462_ (.B1(_03246_),
    .Y(_03247_),
    .A1(_03242_),
    .A2(_03243_));
 sg13g2_a21oi_1 _24463_ (.A1(net9101),
    .A2(_10746_),
    .Y(_03248_),
    .B1(net9628));
 sg13g2_o21ai_1 _24464_ (.B1(_03248_),
    .Y(_03249_),
    .A1(net9101),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][13] ));
 sg13g2_nor2_1 _24465_ (.A(net9101),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][13] ),
    .Y(_03250_));
 sg13g2_a21oi_1 _24466_ (.A1(net9101),
    .A2(_10747_),
    .Y(_03251_),
    .B1(_03250_));
 sg13g2_a21oi_1 _24467_ (.A1(net9628),
    .A2(_03251_),
    .Y(_03252_),
    .B1(net9109));
 sg13g2_mux4_1 _24468_ (.S0(net9680),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][13] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][13] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][13] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][13] ),
    .S1(net9623),
    .X(_03253_));
 sg13g2_o21ai_1 _24469_ (.B1(net9561),
    .Y(_03254_),
    .A1(net9577),
    .A2(_03253_));
 sg13g2_a21o_1 _24470_ (.A2(_03252_),
    .A1(_03249_),
    .B1(_03254_),
    .X(_03255_));
 sg13g2_mux4_1 _24471_ (.S0(net9685),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][13] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][13] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][13] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][13] ),
    .S1(net9628),
    .X(_03256_));
 sg13g2_mux4_1 _24472_ (.S0(net9680),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][13] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][13] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][13] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][13] ),
    .S1(net9623),
    .X(_03257_));
 sg13g2_a221oi_1 _24473_ (.B2(net8817),
    .C1(net9113),
    .B1(_03257_),
    .A1(net8954),
    .Y(_03258_),
    .A2(_03256_));
 sg13g2_nand2_1 _24474_ (.Y(_03259_),
    .A(net8595),
    .B(_03247_));
 sg13g2_a21oi_2 _24475_ (.B1(_03259_),
    .Y(_00755_),
    .A2(_03258_),
    .A1(_03255_));
 sg13g2_a21oi_1 _24476_ (.A1(net9086),
    .A2(_10749_),
    .Y(_03260_),
    .B1(net9598));
 sg13g2_o21ai_1 _24477_ (.B1(_03260_),
    .Y(_03261_),
    .A1(net9086),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][14] ));
 sg13g2_mux2_1 _24478_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][14] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][14] ),
    .S(net9657),
    .X(_03262_));
 sg13g2_a21oi_1 _24479_ (.A1(net9599),
    .A2(_03262_),
    .Y(_03263_),
    .B1(net9110));
 sg13g2_mux4_1 _24480_ (.S0(net9657),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][14] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][14] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][14] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][14] ),
    .S1(net9599),
    .X(_03264_));
 sg13g2_o21ai_1 _24481_ (.B1(net9555),
    .Y(_03265_),
    .A1(net9569),
    .A2(_03264_));
 sg13g2_a21o_1 _24482_ (.A2(_03263_),
    .A1(_03261_),
    .B1(_03265_),
    .X(_03266_));
 sg13g2_mux4_1 _24483_ (.S0(net9660),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][14] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][14] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][14] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][14] ),
    .S1(net9602),
    .X(_03267_));
 sg13g2_mux4_1 _24484_ (.S0(net9660),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][14] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][14] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][14] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][14] ),
    .S1(net9602),
    .X(_03268_));
 sg13g2_a221oi_1 _24485_ (.B2(net8811),
    .C1(net9552),
    .B1(_03268_),
    .A1(net8948),
    .Y(_03269_),
    .A2(_03267_));
 sg13g2_a21oi_1 _24486_ (.A1(net9087),
    .A2(_10751_),
    .Y(_03270_),
    .B1(net9598));
 sg13g2_o21ai_1 _24487_ (.B1(_03270_),
    .Y(_03271_),
    .A1(net9086),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][14] ));
 sg13g2_o21ai_1 _24488_ (.B1(net9599),
    .Y(_03272_),
    .A1(net9657),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][14] ));
 sg13g2_a21oi_1 _24489_ (.A1(net9657),
    .A2(_10752_),
    .Y(_03273_),
    .B1(_03272_));
 sg13g2_nor2_1 _24490_ (.A(net9110),
    .B(_03273_),
    .Y(_03274_));
 sg13g2_mux4_1 _24491_ (.S0(net9659),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][14] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][14] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][14] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][14] ),
    .S1(net9598),
    .X(_03275_));
 sg13g2_o21ai_1 _24492_ (.B1(net9555),
    .Y(_03276_),
    .A1(net9569),
    .A2(_03275_));
 sg13g2_a21oi_1 _24493_ (.A1(_03271_),
    .A2(_03274_),
    .Y(_03277_),
    .B1(_03276_));
 sg13g2_mux4_1 _24494_ (.S0(net9656),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][14] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][14] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][14] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][14] ),
    .S1(net9598),
    .X(_03278_));
 sg13g2_mux4_1 _24495_ (.S0(net9656),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][14] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][14] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][14] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][14] ),
    .S1(net9598),
    .X(_03279_));
 sg13g2_a221oi_1 _24496_ (.B2(net8811),
    .C1(_03277_),
    .B1(_03279_),
    .A1(net8948),
    .Y(_03280_),
    .A2(_03278_));
 sg13g2_a221oi_1 _24497_ (.B2(net9552),
    .C1(net8597),
    .B1(_03280_),
    .A1(_03266_),
    .Y(_00756_),
    .A2(_03269_));
 sg13g2_mux4_1 _24498_ (.S0(net9647),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][15] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][15] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][15] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][15] ),
    .S1(net9588),
    .X(_03281_));
 sg13g2_nor2_1 _24499_ (.A(net9565),
    .B(_03281_),
    .Y(_03282_));
 sg13g2_nor2_1 _24500_ (.A(net9091),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][15] ),
    .Y(_03283_));
 sg13g2_nor2_1 _24501_ (.A(net9648),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][15] ),
    .Y(_03284_));
 sg13g2_nor3_1 _24502_ (.A(net9588),
    .B(_03283_),
    .C(_03284_),
    .Y(_03285_));
 sg13g2_nor2_1 _24503_ (.A(net9648),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][15] ),
    .Y(_03286_));
 sg13g2_o21ai_1 _24504_ (.B1(net9588),
    .Y(_03287_),
    .A1(net9080),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][15] ));
 sg13g2_o21ai_1 _24505_ (.B1(net9565),
    .Y(_03288_),
    .A1(_03286_),
    .A2(_03287_));
 sg13g2_o21ai_1 _24506_ (.B1(net9553),
    .Y(_03289_),
    .A1(_03285_),
    .A2(_03288_));
 sg13g2_mux4_1 _24507_ (.S0(net9649),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][15] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][15] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][15] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][15] ),
    .S1(net9590),
    .X(_03290_));
 sg13g2_mux2_1 _24508_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][15] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][15] ),
    .S(net9647),
    .X(_03291_));
 sg13g2_mux2_1 _24509_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][15] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][15] ),
    .S(net9647),
    .X(_03292_));
 sg13g2_a21o_1 _24510_ (.A2(_03292_),
    .A1(net8674),
    .B1(net9546),
    .X(_03293_));
 sg13g2_a221oi_1 _24511_ (.B2(_02899_),
    .C1(_03293_),
    .B1(_03291_),
    .A1(net8808),
    .Y(_03294_),
    .A2(_03290_));
 sg13g2_o21ai_1 _24512_ (.B1(_03294_),
    .Y(_03295_),
    .A1(_03282_),
    .A2(_03289_));
 sg13g2_mux4_1 _24513_ (.S0(net9649),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][15] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][15] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][15] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][15] ),
    .S1(net9590),
    .X(_03296_));
 sg13g2_nor2_1 _24514_ (.A(net9565),
    .B(_03296_),
    .Y(_03297_));
 sg13g2_nor2_1 _24515_ (.A(net9085),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][15] ),
    .Y(_03298_));
 sg13g2_nor2_1 _24516_ (.A(net9652),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][15] ),
    .Y(_03299_));
 sg13g2_nor3_1 _24517_ (.A(net9596),
    .B(_03298_),
    .C(_03299_),
    .Y(_03300_));
 sg13g2_nor2_1 _24518_ (.A(net9655),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][15] ),
    .Y(_03301_));
 sg13g2_o21ai_1 _24519_ (.B1(net9596),
    .Y(_03302_),
    .A1(net9085),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][15] ));
 sg13g2_o21ai_1 _24520_ (.B1(net9567),
    .Y(_03303_),
    .A1(_03301_),
    .A2(_03302_));
 sg13g2_o21ai_1 _24521_ (.B1(net9554),
    .Y(_03304_),
    .A1(_03300_),
    .A2(_03303_));
 sg13g2_mux4_1 _24522_ (.S0(net9652),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][15] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][15] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][15] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][15] ),
    .S1(net9593),
    .X(_03305_));
 sg13g2_mux4_1 _24523_ (.S0(net9655),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][15] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][15] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][15] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][15] ),
    .S1(net9593),
    .X(_03306_));
 sg13g2_a22oi_1 _24524_ (.Y(_03307_),
    .B1(_03306_),
    .B2(net8810),
    .A2(_03305_),
    .A1(net8947));
 sg13g2_o21ai_1 _24525_ (.B1(_03307_),
    .Y(_03308_),
    .A1(_03297_),
    .A2(_03304_));
 sg13g2_o21ai_1 _24526_ (.B1(_03295_),
    .Y(_03309_),
    .A1(net9111),
    .A2(_03308_));
 sg13g2_nor2_1 _24527_ (.A(net8597),
    .B(_03309_),
    .Y(_00757_));
 sg13g2_nor2_1 _24528_ (.A(net9079),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][16] ),
    .Y(_03310_));
 sg13g2_nor2_1 _24529_ (.A(net9645),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][16] ),
    .Y(_03311_));
 sg13g2_nor3_1 _24530_ (.A(net9585),
    .B(_03310_),
    .C(_03311_),
    .Y(_03312_));
 sg13g2_nor2_1 _24531_ (.A(net9644),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][16] ),
    .Y(_03313_));
 sg13g2_o21ai_1 _24532_ (.B1(net9586),
    .Y(_03314_),
    .A1(net9079),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][16] ));
 sg13g2_o21ai_1 _24533_ (.B1(net9564),
    .Y(_03315_),
    .A1(_03313_),
    .A2(_03314_));
 sg13g2_mux4_1 _24534_ (.S0(net9642),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][16] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][16] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][16] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][16] ),
    .S1(net9583),
    .X(_03316_));
 sg13g2_nor2_1 _24535_ (.A(net9564),
    .B(_03316_),
    .Y(_03317_));
 sg13g2_o21ai_1 _24536_ (.B1(net9553),
    .Y(_03318_),
    .A1(_03312_),
    .A2(_03315_));
 sg13g2_mux4_1 _24537_ (.S0(net9642),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][16] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][16] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][16] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][16] ),
    .S1(net9584),
    .X(_03319_));
 sg13g2_mux4_1 _24538_ (.S0(net9643),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][16] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][16] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][16] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][16] ),
    .S1(net9584),
    .X(_03320_));
 sg13g2_a221oi_1 _24539_ (.B2(net8808),
    .C1(net9546),
    .B1(_03320_),
    .A1(net8946),
    .Y(_03321_),
    .A2(_03319_));
 sg13g2_o21ai_1 _24540_ (.B1(_03321_),
    .Y(_03322_),
    .A1(_03317_),
    .A2(_03318_));
 sg13g2_a21oi_1 _24541_ (.A1(net9081),
    .A2(_10758_),
    .Y(_03323_),
    .B1(net9592));
 sg13g2_o21ai_1 _24542_ (.B1(_03323_),
    .Y(_03324_),
    .A1(net9081),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][16] ));
 sg13g2_nor2_1 _24543_ (.A(net9081),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][16] ),
    .Y(_03325_));
 sg13g2_a21oi_1 _24544_ (.A1(net9081),
    .A2(_10759_),
    .Y(_03326_),
    .B1(_03325_));
 sg13g2_a21oi_1 _24545_ (.A1(net9591),
    .A2(_03326_),
    .Y(_03327_),
    .B1(net9110));
 sg13g2_mux4_1 _24546_ (.S0(net9647),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][16] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][16] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][16] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][16] ),
    .S1(net9588),
    .X(_03328_));
 sg13g2_o21ai_1 _24547_ (.B1(net9554),
    .Y(_03329_),
    .A1(net9565),
    .A2(_03328_));
 sg13g2_a21o_1 _24548_ (.A2(_03327_),
    .A1(_03324_),
    .B1(_03329_),
    .X(_03330_));
 sg13g2_mux4_1 _24549_ (.S0(net9648),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][16] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][16] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][16] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][16] ),
    .S1(net9589),
    .X(_03331_));
 sg13g2_mux4_1 _24550_ (.S0(net9644),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][16] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][16] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][16] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][16] ),
    .S1(net9585),
    .X(_03332_));
 sg13g2_a221oi_1 _24551_ (.B2(net8809),
    .C1(net9111),
    .B1(_03332_),
    .A1(net8947),
    .Y(_03333_),
    .A2(_03331_));
 sg13g2_nand2_1 _24552_ (.Y(_03334_),
    .A(net8594),
    .B(_03322_));
 sg13g2_a21oi_2 _24553_ (.B1(_03334_),
    .Y(_00758_),
    .A2(_03333_),
    .A1(_03330_));
 sg13g2_mux4_1 _24554_ (.S0(net9647),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][17] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][17] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][17] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][17] ),
    .S1(net9588),
    .X(_03335_));
 sg13g2_nor2_1 _24555_ (.A(net9081),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][17] ),
    .Y(_03336_));
 sg13g2_nor2_1 _24556_ (.A(net9650),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][17] ),
    .Y(_03337_));
 sg13g2_nor3_1 _24557_ (.A(net9591),
    .B(_03336_),
    .C(_03337_),
    .Y(_03338_));
 sg13g2_nor2_1 _24558_ (.A(net9650),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][17] ),
    .Y(_03339_));
 sg13g2_o21ai_1 _24559_ (.B1(net9591),
    .Y(_03340_),
    .A1(net9080),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][17] ));
 sg13g2_o21ai_1 _24560_ (.B1(net9565),
    .Y(_03341_),
    .A1(_03339_),
    .A2(_03340_));
 sg13g2_o21ai_1 _24561_ (.B1(net9554),
    .Y(_03342_),
    .A1(_03338_),
    .A2(_03341_));
 sg13g2_inv_1 _24562_ (.Y(_03343_),
    .A(_03342_));
 sg13g2_o21ai_1 _24563_ (.B1(_03343_),
    .Y(_03344_),
    .A1(net9565),
    .A2(_03335_));
 sg13g2_mux4_1 _24564_ (.S0(net9648),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][17] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][17] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][17] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][17] ),
    .S1(net9589),
    .X(_03345_));
 sg13g2_mux4_1 _24565_ (.S0(net9644),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][17] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][17] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][17] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][17] ),
    .S1(net9585),
    .X(_03346_));
 sg13g2_a221oi_1 _24566_ (.B2(net8809),
    .C1(net9111),
    .B1(_03346_),
    .A1(net8947),
    .Y(_03347_),
    .A2(_03345_));
 sg13g2_a21oi_1 _24567_ (.A1(net9079),
    .A2(_10761_),
    .Y(_03348_),
    .B1(net9584));
 sg13g2_o21ai_1 _24568_ (.B1(_03348_),
    .Y(_03349_),
    .A1(net9079),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][17] ));
 sg13g2_mux2_1 _24569_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][17] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][17] ),
    .S(net9643),
    .X(_03350_));
 sg13g2_a21oi_1 _24570_ (.A1(net9586),
    .A2(_03350_),
    .Y(_03351_),
    .B1(net9110));
 sg13g2_mux4_1 _24571_ (.S0(net9643),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][17] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][17] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][17] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][17] ),
    .S1(net9584),
    .X(_03352_));
 sg13g2_o21ai_1 _24572_ (.B1(net9553),
    .Y(_03353_),
    .A1(net9564),
    .A2(_03352_));
 sg13g2_a21oi_1 _24573_ (.A1(_03349_),
    .A2(_03351_),
    .Y(_03354_),
    .B1(_03353_));
 sg13g2_mux4_1 _24574_ (.S0(net9643),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][17] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][17] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][17] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][17] ),
    .S1(net9584),
    .X(_03355_));
 sg13g2_mux4_1 _24575_ (.S0(net9643),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][17] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][17] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][17] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][17] ),
    .S1(net9584),
    .X(_03356_));
 sg13g2_a221oi_1 _24576_ (.B2(net8808),
    .C1(_03354_),
    .B1(_03356_),
    .A1(net8946),
    .Y(_03357_),
    .A2(_03355_));
 sg13g2_a221oi_1 _24577_ (.B2(net9111),
    .C1(net8597),
    .B1(_03357_),
    .A1(_03344_),
    .Y(_00759_),
    .A2(_03347_));
 sg13g2_mux4_1 _24578_ (.S0(net9644),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][18] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][18] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][18] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][18] ),
    .S1(net9585),
    .X(_03358_));
 sg13g2_nor2_1 _24579_ (.A(net9566),
    .B(_03358_),
    .Y(_03359_));
 sg13g2_nor2_1 _24580_ (.A(net9080),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][18] ),
    .Y(_03360_));
 sg13g2_nor2_1 _24581_ (.A(net9643),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][18] ),
    .Y(_03361_));
 sg13g2_nor3_1 _24582_ (.A(net9583),
    .B(_03360_),
    .C(_03361_),
    .Y(_03362_));
 sg13g2_nor2_1 _24583_ (.A(net9646),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][18] ),
    .Y(_03363_));
 sg13g2_o21ai_1 _24584_ (.B1(net9587),
    .Y(_03364_),
    .A1(net9080),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][18] ));
 sg13g2_o21ai_1 _24585_ (.B1(net9564),
    .Y(_03365_),
    .A1(_03363_),
    .A2(_03364_));
 sg13g2_o21ai_1 _24586_ (.B1(net9553),
    .Y(_03366_),
    .A1(_03362_),
    .A2(_03365_));
 sg13g2_mux4_1 _24587_ (.S0(net9646),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][18] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][18] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][18] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][18] ),
    .S1(net9587),
    .X(_03367_));
 sg13g2_mux4_1 _24588_ (.S0(net9646),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][18] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][18] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][18] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][18] ),
    .S1(net9587),
    .X(_03368_));
 sg13g2_a221oi_1 _24589_ (.B2(net8946),
    .C1(net9546),
    .B1(_03368_),
    .A1(net8808),
    .Y(_03369_),
    .A2(_03367_));
 sg13g2_o21ai_1 _24590_ (.B1(_03369_),
    .Y(_03370_),
    .A1(_03359_),
    .A2(_03366_));
 sg13g2_nor2_1 _24591_ (.A(net9082),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][18] ),
    .Y(_03371_));
 sg13g2_nor2_1 _24592_ (.A(net9654),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][18] ),
    .Y(_03372_));
 sg13g2_nor3_1 _24593_ (.A(net9594),
    .B(_03371_),
    .C(_03372_),
    .Y(_03373_));
 sg13g2_nor2_1 _24594_ (.A(net9654),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][18] ),
    .Y(_03374_));
 sg13g2_o21ai_1 _24595_ (.B1(net9594),
    .Y(_03375_),
    .A1(net9082),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][18] ));
 sg13g2_o21ai_1 _24596_ (.B1(net9567),
    .Y(_03376_),
    .A1(_03374_),
    .A2(_03375_));
 sg13g2_mux4_1 _24597_ (.S0(net9650),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][18] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][18] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][18] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][18] ),
    .S1(net9591),
    .X(_03377_));
 sg13g2_nor2_1 _24598_ (.A(net9567),
    .B(_03377_),
    .Y(_03378_));
 sg13g2_o21ai_1 _24599_ (.B1(net9556),
    .Y(_03379_),
    .A1(_03373_),
    .A2(_03376_));
 sg13g2_a22oi_1 _24600_ (.Y(_03380_),
    .B1(_02899_),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][18] ),
    .A2(net8674),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][18] ));
 sg13g2_o21ai_1 _24601_ (.B1(net9547),
    .Y(_03381_),
    .A1(net9653),
    .A2(_03380_));
 sg13g2_mux4_1 _24602_ (.S0(net9651),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][18] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][18] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][18] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][18] ),
    .S1(net9592),
    .X(_03382_));
 sg13g2_a22oi_1 _24603_ (.Y(_03383_),
    .B1(_02899_),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][18] ),
    .A2(net8674),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][18] ));
 sg13g2_inv_1 _24604_ (.Y(_03384_),
    .A(_03383_));
 sg13g2_a221oi_1 _24605_ (.B2(net9653),
    .C1(_03381_),
    .B1(_03384_),
    .A1(net8810),
    .Y(_03385_),
    .A2(_03382_));
 sg13g2_o21ai_1 _24606_ (.B1(_03385_),
    .Y(_03386_),
    .A1(_03378_),
    .A2(_03379_));
 sg13g2_and3_2 _24607_ (.X(_00760_),
    .A(net8594),
    .B(_03370_),
    .C(_03386_));
 sg13g2_nor2_1 _24608_ (.A(net9086),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][19] ),
    .Y(_03387_));
 sg13g2_nor2_1 _24609_ (.A(net9656),
    .B(net3124),
    .Y(_03388_));
 sg13g2_nor3_1 _24610_ (.A(net9597),
    .B(_03387_),
    .C(_03388_),
    .Y(_03389_));
 sg13g2_nor2_1 _24611_ (.A(net9656),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][19] ),
    .Y(_03390_));
 sg13g2_o21ai_1 _24612_ (.B1(net9597),
    .Y(_03391_),
    .A1(net9086),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][19] ));
 sg13g2_o21ai_1 _24613_ (.B1(net9569),
    .Y(_03392_),
    .A1(_03390_),
    .A2(_03391_));
 sg13g2_a21oi_1 _24614_ (.A1(net9086),
    .A2(_10766_),
    .Y(_03393_),
    .B1(net9597));
 sg13g2_o21ai_1 _24615_ (.B1(_03393_),
    .Y(_03394_),
    .A1(net9086),
    .A2(net5563));
 sg13g2_mux2_1 _24616_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][19] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][19] ),
    .S(net9656),
    .X(_03395_));
 sg13g2_a21oi_1 _24617_ (.A1(net9597),
    .A2(_03395_),
    .Y(_03396_),
    .B1(net9569));
 sg13g2_a21oi_1 _24618_ (.A1(_03394_),
    .A2(_03396_),
    .Y(_03397_),
    .B1(_10462_));
 sg13g2_o21ai_1 _24619_ (.B1(_03397_),
    .Y(_03398_),
    .A1(_03389_),
    .A2(_03392_));
 sg13g2_mux4_1 _24620_ (.S0(net9653),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][19] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][19] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][19] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][19] ),
    .S1(net9594),
    .X(_03399_));
 sg13g2_mux4_1 _24621_ (.S0(net9656),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][19] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][19] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][19] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][19] ),
    .S1(net9597),
    .X(_03400_));
 sg13g2_a221oi_1 _24622_ (.B2(net8810),
    .C1(net9546),
    .B1(_03400_),
    .A1(net8947),
    .Y(_03401_),
    .A2(_03399_));
 sg13g2_a21oi_1 _24623_ (.A1(net9082),
    .A2(_10769_),
    .Y(_03402_),
    .B1(net9597));
 sg13g2_o21ai_1 _24624_ (.B1(_03402_),
    .Y(_03403_),
    .A1(net9082),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][19] ));
 sg13g2_nor2_1 _24625_ (.A(net9082),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][19] ),
    .Y(_03404_));
 sg13g2_a21oi_1 _24626_ (.A1(net9086),
    .A2(_10770_),
    .Y(_03405_),
    .B1(_03404_));
 sg13g2_a21oi_1 _24627_ (.A1(net9597),
    .A2(_03405_),
    .Y(_03406_),
    .B1(net9110));
 sg13g2_mux4_1 _24628_ (.S0(net9653),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][19] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][19] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][19] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][19] ),
    .S1(net9594),
    .X(_03407_));
 sg13g2_o21ai_1 _24629_ (.B1(net9554),
    .Y(_03408_),
    .A1(net9567),
    .A2(_03407_));
 sg13g2_a21o_1 _24630_ (.A2(_03406_),
    .A1(_03403_),
    .B1(_03408_),
    .X(_03409_));
 sg13g2_a22oi_1 _24631_ (.Y(_03410_),
    .B1(_02899_),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][19] ),
    .A2(net8674),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][19] ));
 sg13g2_a22oi_1 _24632_ (.Y(_03411_),
    .B1(_02899_),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][19] ),
    .A2(net8674),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][19] ));
 sg13g2_mux2_1 _24633_ (.A0(_03410_),
    .A1(_03411_),
    .S(net9082),
    .X(_03412_));
 sg13g2_mux4_1 _24634_ (.S0(net9653),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][19] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][19] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][19] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][19] ),
    .S1(net9594),
    .X(_03413_));
 sg13g2_nand3_1 _24635_ (.B(_03409_),
    .C(_03412_),
    .A(net9546),
    .Y(_03414_));
 sg13g2_a21oi_1 _24636_ (.A1(net8810),
    .A2(_03413_),
    .Y(_03415_),
    .B1(_03414_));
 sg13g2_a221oi_1 _24637_ (.B2(_03401_),
    .C1(_03415_),
    .B1(_03398_),
    .A1(net8674),
    .Y(_00761_),
    .A2(_02903_));
 sg13g2_a21oi_1 _24638_ (.A1(net9097),
    .A2(_10771_),
    .Y(_03416_),
    .B1(net9619));
 sg13g2_o21ai_1 _24639_ (.B1(_03416_),
    .Y(_03417_),
    .A1(net9097),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][20] ));
 sg13g2_mux2_1 _24640_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][20] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][20] ),
    .S(net9677),
    .X(_03418_));
 sg13g2_a21oi_1 _24641_ (.A1(net9619),
    .A2(_03418_),
    .Y(_03419_),
    .B1(net9575));
 sg13g2_nor2_1 _24642_ (.A(net9097),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][20] ),
    .Y(_03420_));
 sg13g2_nor2_1 _24643_ (.A(net9677),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][20] ),
    .Y(_03421_));
 sg13g2_nor3_1 _24644_ (.A(net9619),
    .B(_03420_),
    .C(_03421_),
    .Y(_03422_));
 sg13g2_nor2_1 _24645_ (.A(net9677),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][20] ),
    .Y(_03423_));
 sg13g2_o21ai_1 _24646_ (.B1(net9619),
    .Y(_03424_),
    .A1(net9097),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][20] ));
 sg13g2_o21ai_1 _24647_ (.B1(net9575),
    .Y(_03425_),
    .A1(_03423_),
    .A2(_03424_));
 sg13g2_o21ai_1 _24648_ (.B1(net9559),
    .Y(_03426_),
    .A1(_03422_),
    .A2(_03425_));
 sg13g2_a21o_1 _24649_ (.A2(_03419_),
    .A1(_03417_),
    .B1(_03426_),
    .X(_03427_));
 sg13g2_mux4_1 _24650_ (.S0(net9673),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][20] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][20] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][20] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][20] ),
    .S1(net9618),
    .X(_03428_));
 sg13g2_mux4_1 _24651_ (.S0(net9673),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][20] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][20] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][20] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][20] ),
    .S1(net9616),
    .X(_03429_));
 sg13g2_a221oi_1 _24652_ (.B2(net8951),
    .C1(net9549),
    .B1(_03429_),
    .A1(net8813),
    .Y(_03430_),
    .A2(_03428_));
 sg13g2_a21oi_1 _24653_ (.A1(net9096),
    .A2(_10773_),
    .Y(_03431_),
    .B1(net9621));
 sg13g2_o21ai_1 _24654_ (.B1(_03431_),
    .Y(_03432_),
    .A1(net9096),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][20] ));
 sg13g2_nor2_1 _24655_ (.A(net9096),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][20] ),
    .Y(_03433_));
 sg13g2_a21oi_1 _24656_ (.A1(net9096),
    .A2(_10774_),
    .Y(_03434_),
    .B1(_03433_));
 sg13g2_a21oi_1 _24657_ (.A1(net9619),
    .A2(_03434_),
    .Y(_03435_),
    .B1(net9109));
 sg13g2_mux4_1 _24658_ (.S0(net9677),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][20] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][20] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][20] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][20] ),
    .S1(net9619),
    .X(_03436_));
 sg13g2_o21ai_1 _24659_ (.B1(net9559),
    .Y(_03437_),
    .A1(net9575),
    .A2(_03436_));
 sg13g2_a21o_1 _24660_ (.A2(_03435_),
    .A1(_03432_),
    .B1(_03437_),
    .X(_03438_));
 sg13g2_mux4_1 _24661_ (.S0(net9673),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][20] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][20] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][20] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][20] ),
    .S1(net9616),
    .X(_03439_));
 sg13g2_mux4_1 _24662_ (.S0(net9674),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][20] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][20] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][20] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][20] ),
    .S1(net9617),
    .X(_03440_));
 sg13g2_a221oi_1 _24663_ (.B2(net8813),
    .C1(net9115),
    .B1(_03440_),
    .A1(net8950),
    .Y(_03441_),
    .A2(_03439_));
 sg13g2_a221oi_1 _24664_ (.B2(_03441_),
    .C1(net8597),
    .B1(_03438_),
    .A1(_03427_),
    .Y(_00762_),
    .A2(_03430_));
 sg13g2_nor2_1 _24665_ (.A(net9092),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][21] ),
    .Y(_03442_));
 sg13g2_nor2_1 _24666_ (.A(net9666),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][21] ),
    .Y(_03443_));
 sg13g2_nor3_1 _24667_ (.A(net9608),
    .B(_03442_),
    .C(_03443_),
    .Y(_03444_));
 sg13g2_nor2_1 _24668_ (.A(net9665),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][21] ),
    .Y(_03445_));
 sg13g2_o21ai_1 _24669_ (.B1(net9608),
    .Y(_03446_),
    .A1(net9092),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][21] ));
 sg13g2_o21ai_1 _24670_ (.B1(net9571),
    .Y(_03447_),
    .A1(_03445_),
    .A2(_03446_));
 sg13g2_mux4_1 _24671_ (.S0(net9665),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][21] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][21] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][21] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][21] ),
    .S1(net9609),
    .X(_03448_));
 sg13g2_nor2_1 _24672_ (.A(net9571),
    .B(_03448_),
    .Y(_03449_));
 sg13g2_o21ai_1 _24673_ (.B1(net9557),
    .Y(_03450_),
    .A1(_03444_),
    .A2(_03447_));
 sg13g2_mux4_1 _24674_ (.S0(net9665),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][21] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][21] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][21] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][21] ),
    .S1(net9609),
    .X(_03451_));
 sg13g2_mux4_1 _24675_ (.S0(net9666),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][21] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][21] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][21] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][21] ),
    .S1(net9608),
    .X(_03452_));
 sg13g2_a221oi_1 _24676_ (.B2(net8812),
    .C1(net9548),
    .B1(_03452_),
    .A1(net8950),
    .Y(_03453_),
    .A2(_03451_));
 sg13g2_o21ai_1 _24677_ (.B1(_03453_),
    .Y(_03454_),
    .A1(_03449_),
    .A2(_03450_));
 sg13g2_a21oi_1 _24678_ (.A1(net9089),
    .A2(_10777_),
    .Y(_03455_),
    .B1(net9605));
 sg13g2_o21ai_1 _24679_ (.B1(_03455_),
    .Y(_03456_),
    .A1(net9089),
    .A2(net3547));
 sg13g2_nor2_1 _24680_ (.A(net9089),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][21] ),
    .Y(_03457_));
 sg13g2_a21oi_1 _24681_ (.A1(net9089),
    .A2(_10778_),
    .Y(_03458_),
    .B1(_03457_));
 sg13g2_a21oi_1 _24682_ (.A1(net9605),
    .A2(_03458_),
    .Y(_03459_),
    .B1(net9108));
 sg13g2_mux4_1 _24683_ (.S0(net9666),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][21] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][21] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][21] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][21] ),
    .S1(net9608),
    .X(_03460_));
 sg13g2_o21ai_1 _24684_ (.B1(net9555),
    .Y(_03461_),
    .A1(net9570),
    .A2(_03460_));
 sg13g2_a21o_1 _24685_ (.A2(_03459_),
    .A1(_03456_),
    .B1(_03461_),
    .X(_03462_));
 sg13g2_mux4_1 _24686_ (.S0(net9666),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][21] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][21] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][21] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][21] ),
    .S1(net9608),
    .X(_03463_));
 sg13g2_mux4_1 _24687_ (.S0(net9662),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][21] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][21] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][21] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][21] ),
    .S1(net9605),
    .X(_03464_));
 sg13g2_a221oi_1 _24688_ (.B2(net8811),
    .C1(net9112),
    .B1(_03464_),
    .A1(net8948),
    .Y(_03465_),
    .A2(_03463_));
 sg13g2_nand2_1 _24689_ (.Y(_03466_),
    .A(net8596),
    .B(_03454_));
 sg13g2_a21oi_1 _24690_ (.A1(_03462_),
    .A2(_03465_),
    .Y(_00763_),
    .B1(_03466_));
 sg13g2_mux4_1 _24691_ (.S0(net9692),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][22] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][22] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][22] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][22] ),
    .S1(net9636),
    .X(_03467_));
 sg13g2_nor2_1 _24692_ (.A(net9578),
    .B(_03467_),
    .Y(_03468_));
 sg13g2_nor2_1 _24693_ (.A(net9103),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][22] ),
    .Y(_03469_));
 sg13g2_nor2_1 _24694_ (.A(net9692),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][22] ),
    .Y(_03470_));
 sg13g2_nor3_1 _24695_ (.A(net9636),
    .B(_03469_),
    .C(_03470_),
    .Y(_03471_));
 sg13g2_nor2_1 _24696_ (.A(net9692),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][22] ),
    .Y(_03472_));
 sg13g2_o21ai_1 _24697_ (.B1(net9636),
    .Y(_03473_),
    .A1(net9103),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][22] ));
 sg13g2_o21ai_1 _24698_ (.B1(net9579),
    .Y(_03474_),
    .A1(_03472_),
    .A2(_03473_));
 sg13g2_o21ai_1 _24699_ (.B1(net9560),
    .Y(_03475_),
    .A1(_03471_),
    .A2(_03474_));
 sg13g2_mux4_1 _24700_ (.S0(net9692),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][22] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][22] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][22] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][22] ),
    .S1(net9636),
    .X(_03476_));
 sg13g2_mux4_1 _24701_ (.S0(net9692),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][22] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][22] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][22] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][22] ),
    .S1(net9637),
    .X(_03477_));
 sg13g2_a221oi_1 _24702_ (.B2(net8952),
    .C1(net9550),
    .B1(_03477_),
    .A1(net8815),
    .Y(_03478_),
    .A2(_03476_));
 sg13g2_o21ai_1 _24703_ (.B1(_03478_),
    .Y(_03479_),
    .A1(_03468_),
    .A2(_03475_));
 sg13g2_mux4_1 _24704_ (.S0(net9687),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][22] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][22] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][22] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][22] ),
    .S1(net9630),
    .X(_03480_));
 sg13g2_nor2_1 _24705_ (.A(net9578),
    .B(_03480_),
    .Y(_03481_));
 sg13g2_nor2_1 _24706_ (.A(net9104),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][22] ),
    .Y(_03482_));
 sg13g2_nor2_1 _24707_ (.A(net9691),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][22] ),
    .Y(_03483_));
 sg13g2_nor3_1 _24708_ (.A(net9638),
    .B(_03482_),
    .C(_03483_),
    .Y(_03484_));
 sg13g2_nor2_1 _24709_ (.A(net9691),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][22] ),
    .Y(_03485_));
 sg13g2_o21ai_1 _24710_ (.B1(net9638),
    .Y(_03486_),
    .A1(net9104),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][22] ));
 sg13g2_o21ai_1 _24711_ (.B1(net9578),
    .Y(_03487_),
    .A1(_03485_),
    .A2(_03486_));
 sg13g2_o21ai_1 _24712_ (.B1(net9560),
    .Y(_03488_),
    .A1(_03484_),
    .A2(_03487_));
 sg13g2_mux4_1 _24713_ (.S0(net9686),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][22] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][22] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][22] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][22] ),
    .S1(net9631),
    .X(_03489_));
 sg13g2_mux4_1 _24714_ (.S0(net9687),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][22] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][22] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][22] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][22] ),
    .S1(net9630),
    .X(_03490_));
 sg13g2_a221oi_1 _24715_ (.B2(net8953),
    .C1(net9114),
    .B1(_03490_),
    .A1(net8815),
    .Y(_03491_),
    .A2(_03489_));
 sg13g2_o21ai_1 _24716_ (.B1(_03491_),
    .Y(_03492_),
    .A1(_03481_),
    .A2(_03488_));
 sg13g2_and3_2 _24717_ (.X(_00764_),
    .A(net8595),
    .B(_03479_),
    .C(_03492_));
 sg13g2_a21oi_1 _24718_ (.A1(net9080),
    .A2(_10785_),
    .Y(_03493_),
    .B1(net9590));
 sg13g2_o21ai_1 _24719_ (.B1(_03493_),
    .Y(_03494_),
    .A1(net9080),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][23] ));
 sg13g2_mux2_1 _24720_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][23] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][23] ),
    .S(net9649),
    .X(_03495_));
 sg13g2_a21oi_1 _24721_ (.A1(net9590),
    .A2(_03495_),
    .Y(_03496_),
    .B1(net9110));
 sg13g2_mux4_1 _24722_ (.S0(net9647),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][23] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][23] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][23] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][23] ),
    .S1(net9588),
    .X(_03497_));
 sg13g2_o21ai_1 _24723_ (.B1(net9553),
    .Y(_03498_),
    .A1(net9566),
    .A2(_03497_));
 sg13g2_a21o_1 _24724_ (.A2(_03496_),
    .A1(_03494_),
    .B1(_03498_),
    .X(_03499_));
 sg13g2_mux4_1 _24725_ (.S0(net9647),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][23] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][23] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][23] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][23] ),
    .S1(net9588),
    .X(_03500_));
 sg13g2_mux4_1 _24726_ (.S0(net9649),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][23] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][23] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][23] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][23] ),
    .S1(net9590),
    .X(_03501_));
 sg13g2_a221oi_1 _24727_ (.B2(net8808),
    .C1(net9546),
    .B1(_03501_),
    .A1(net8946),
    .Y(_03502_),
    .A2(_03500_));
 sg13g2_mux4_1 _24728_ (.S0(net9649),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][23] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][23] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][23] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][23] ),
    .S1(net9590),
    .X(_03503_));
 sg13g2_nor2_1 _24729_ (.A(net9080),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][23] ),
    .Y(_03504_));
 sg13g2_nor2_1 _24730_ (.A(net9652),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][23] ),
    .Y(_03505_));
 sg13g2_nor3_1 _24731_ (.A(net9593),
    .B(_03504_),
    .C(_03505_),
    .Y(_03506_));
 sg13g2_nor2_1 _24732_ (.A(net9652),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][23] ),
    .Y(_03507_));
 sg13g2_o21ai_1 _24733_ (.B1(net9593),
    .Y(_03508_),
    .A1(net9081),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][23] ));
 sg13g2_o21ai_1 _24734_ (.B1(net9567),
    .Y(_03509_),
    .A1(_03507_),
    .A2(_03508_));
 sg13g2_o21ai_1 _24735_ (.B1(net9553),
    .Y(_03510_),
    .A1(_03506_),
    .A2(_03509_));
 sg13g2_inv_1 _24736_ (.Y(_03511_),
    .A(_03510_));
 sg13g2_o21ai_1 _24737_ (.B1(_03511_),
    .Y(_03512_),
    .A1(net9566),
    .A2(_03503_));
 sg13g2_mux4_1 _24738_ (.S0(net9652),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][23] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][23] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][23] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][23] ),
    .S1(net9593),
    .X(_03513_));
 sg13g2_mux4_1 _24739_ (.S0(net9650),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][23] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][23] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][23] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][23] ),
    .S1(net9591),
    .X(_03514_));
 sg13g2_a221oi_1 _24740_ (.B2(net8808),
    .C1(net9111),
    .B1(_03514_),
    .A1(net8946),
    .Y(_03515_),
    .A2(_03513_));
 sg13g2_a221oi_1 _24741_ (.B2(_03515_),
    .C1(net8597),
    .B1(_03512_),
    .A1(_03499_),
    .Y(_00765_),
    .A2(_03502_));
 sg13g2_nor2_1 _24742_ (.A(net9092),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][24] ),
    .Y(_03516_));
 sg13g2_nor2_1 _24743_ (.A(net9667),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][24] ),
    .Y(_03517_));
 sg13g2_nor3_1 _24744_ (.A(net9610),
    .B(_03516_),
    .C(_03517_),
    .Y(_03518_));
 sg13g2_nor2_1 _24745_ (.A(net9667),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][24] ),
    .Y(_03519_));
 sg13g2_o21ai_1 _24746_ (.B1(net9610),
    .Y(_03520_),
    .A1(net9092),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][24] ));
 sg13g2_o21ai_1 _24747_ (.B1(net9574),
    .Y(_03521_),
    .A1(_03519_),
    .A2(_03520_));
 sg13g2_mux4_1 _24748_ (.S0(net9667),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][24] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][24] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][24] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][24] ),
    .S1(net9610),
    .X(_03522_));
 sg13g2_nor2_1 _24749_ (.A(net9571),
    .B(_03522_),
    .Y(_03523_));
 sg13g2_o21ai_1 _24750_ (.B1(net9557),
    .Y(_03524_),
    .A1(_03518_),
    .A2(_03521_));
 sg13g2_mux4_1 _24751_ (.S0(net9667),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][24] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][24] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][24] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][24] ),
    .S1(net9610),
    .X(_03525_));
 sg13g2_mux4_1 _24752_ (.S0(net9668),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][24] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][24] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][24] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][24] ),
    .S1(net9611),
    .X(_03526_));
 sg13g2_a221oi_1 _24753_ (.B2(net8812),
    .C1(net9548),
    .B1(_03526_),
    .A1(net8950),
    .Y(_03527_),
    .A2(_03525_));
 sg13g2_o21ai_1 _24754_ (.B1(_03527_),
    .Y(_03528_),
    .A1(_03523_),
    .A2(_03524_));
 sg13g2_mux4_1 _24755_ (.S0(net9665),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][24] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][24] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][24] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][24] ),
    .S1(net9609),
    .X(_03529_));
 sg13g2_nor2_1 _24756_ (.A(net9092),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][24] ),
    .Y(_03530_));
 sg13g2_nor2_1 _24757_ (.A(net9665),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][24] ),
    .Y(_03531_));
 sg13g2_nor3_1 _24758_ (.A(net9609),
    .B(_03530_),
    .C(_03531_),
    .Y(_03532_));
 sg13g2_nor2_1 _24759_ (.A(net9665),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][24] ),
    .Y(_03533_));
 sg13g2_o21ai_1 _24760_ (.B1(net9609),
    .Y(_03534_),
    .A1(net9092),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][24] ));
 sg13g2_o21ai_1 _24761_ (.B1(net9571),
    .Y(_03535_),
    .A1(_03533_),
    .A2(_03534_));
 sg13g2_o21ai_1 _24762_ (.B1(net9557),
    .Y(_03536_),
    .A1(_03532_),
    .A2(_03535_));
 sg13g2_inv_1 _24763_ (.Y(_03537_),
    .A(_03536_));
 sg13g2_o21ai_1 _24764_ (.B1(_03537_),
    .Y(_03538_),
    .A1(net9571),
    .A2(_03529_));
 sg13g2_mux4_1 _24765_ (.S0(net9665),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][24] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][24] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][24] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][24] ),
    .S1(net9608),
    .X(_03539_));
 sg13g2_mux4_1 _24766_ (.S0(net9666),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][24] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][24] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][24] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][24] ),
    .S1(net9608),
    .X(_03540_));
 sg13g2_a221oi_1 _24767_ (.B2(net8812),
    .C1(net9115),
    .B1(_03540_),
    .A1(net8950),
    .Y(_03541_),
    .A2(_03539_));
 sg13g2_nand2_1 _24768_ (.Y(_03542_),
    .A(net8595),
    .B(_03528_));
 sg13g2_a21oi_2 _24769_ (.B1(_03542_),
    .Y(_00766_),
    .A2(_03541_),
    .A1(_03538_));
 sg13g2_mux4_1 _24770_ (.S0(net9678),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][25] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][25] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][25] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][25] ),
    .S1(net9622),
    .X(_03543_));
 sg13g2_nor2_1 _24771_ (.A(net9098),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][25] ),
    .Y(_03544_));
 sg13g2_nor2_1 _24772_ (.A(net9678),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][25] ),
    .Y(_03545_));
 sg13g2_nor3_1 _24773_ (.A(net9622),
    .B(_03544_),
    .C(_03545_),
    .Y(_03546_));
 sg13g2_nor2_1 _24774_ (.A(net9678),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][25] ),
    .Y(_03547_));
 sg13g2_o21ai_1 _24775_ (.B1(net9622),
    .Y(_03548_),
    .A1(net9098),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][25] ));
 sg13g2_o21ai_1 _24776_ (.B1(net9575),
    .Y(_03549_),
    .A1(_03547_),
    .A2(_03548_));
 sg13g2_o21ai_1 _24777_ (.B1(net9559),
    .Y(_03550_),
    .A1(_03546_),
    .A2(_03549_));
 sg13g2_inv_1 _24778_ (.Y(_03551_),
    .A(_03550_));
 sg13g2_o21ai_1 _24779_ (.B1(_03551_),
    .Y(_03552_),
    .A1(net9575),
    .A2(_03543_));
 sg13g2_mux4_1 _24780_ (.S0(net9677),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][25] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][25] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][25] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][25] ),
    .S1(net9619),
    .X(_03553_));
 sg13g2_mux4_1 _24781_ (.S0(net9678),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][25] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][25] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][25] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][25] ),
    .S1(net9622),
    .X(_03554_));
 sg13g2_a221oi_1 _24782_ (.B2(net8951),
    .C1(net9114),
    .B1(_03554_),
    .A1(net8813),
    .Y(_03555_),
    .A2(_03553_));
 sg13g2_mux4_1 _24783_ (.S0(net9673),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][25] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][25] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][25] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][25] ),
    .S1(net9616),
    .X(_03556_));
 sg13g2_nor2_1 _24784_ (.A(net9572),
    .B(_03556_),
    .Y(_03557_));
 sg13g2_nor2_1 _24785_ (.A(net9094),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][25] ),
    .Y(_03558_));
 sg13g2_nor2_1 _24786_ (.A(net9675),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][25] ),
    .Y(_03559_));
 sg13g2_nor3_1 _24787_ (.A(net9618),
    .B(_03558_),
    .C(_03559_),
    .Y(_03560_));
 sg13g2_nor2_1 _24788_ (.A(net9675),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][25] ),
    .Y(_03561_));
 sg13g2_o21ai_1 _24789_ (.B1(net9618),
    .Y(_03562_),
    .A1(net9094),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][25] ));
 sg13g2_o21ai_1 _24790_ (.B1(net9572),
    .Y(_03563_),
    .A1(_03561_),
    .A2(_03562_));
 sg13g2_o21ai_1 _24791_ (.B1(net9558),
    .Y(_03564_),
    .A1(_03560_),
    .A2(_03563_));
 sg13g2_mux4_1 _24792_ (.S0(net9678),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][25] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][25] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][25] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][25] ),
    .S1(net9622),
    .X(_03565_));
 sg13g2_mux4_1 _24793_ (.S0(net9676),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][25] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][25] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][25] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][25] ),
    .S1(net9621),
    .X(_03566_));
 sg13g2_a22oi_1 _24794_ (.Y(_03567_),
    .B1(_03566_),
    .B2(net8954),
    .A2(_03565_),
    .A1(net8814));
 sg13g2_o21ai_1 _24795_ (.B1(_03567_),
    .Y(_03568_),
    .A1(_03557_),
    .A2(_03564_));
 sg13g2_o21ai_1 _24796_ (.B1(net8595),
    .Y(_03569_),
    .A1(net9549),
    .A2(_03568_));
 sg13g2_a21oi_1 _24797_ (.A1(_03552_),
    .A2(_03555_),
    .Y(_00767_),
    .B1(_03569_));
 sg13g2_mux4_1 _24798_ (.S0(net9693),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][26] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][26] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][26] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][26] ),
    .S1(net9637),
    .X(_03570_));
 sg13g2_nor2_1 _24799_ (.A(net9578),
    .B(_03570_),
    .Y(_03571_));
 sg13g2_nor2_1 _24800_ (.A(net9103),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][26] ),
    .Y(_03572_));
 sg13g2_nor2_1 _24801_ (.A(net9692),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][26] ),
    .Y(_03573_));
 sg13g2_nor3_1 _24802_ (.A(net9637),
    .B(_03572_),
    .C(_03573_),
    .Y(_03574_));
 sg13g2_nor2_1 _24803_ (.A(net9693),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][26] ),
    .Y(_03575_));
 sg13g2_o21ai_1 _24804_ (.B1(net9637),
    .Y(_03576_),
    .A1(net9103),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][26] ));
 sg13g2_o21ai_1 _24805_ (.B1(net9579),
    .Y(_03577_),
    .A1(_03575_),
    .A2(_03576_));
 sg13g2_o21ai_1 _24806_ (.B1(net9562),
    .Y(_03578_),
    .A1(_03574_),
    .A2(_03577_));
 sg13g2_mux4_1 _24807_ (.S0(net9693),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][26] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][26] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][26] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][26] ),
    .S1(net9636),
    .X(_03579_));
 sg13g2_mux4_1 _24808_ (.S0(net9692),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][26] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][26] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][26] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][26] ),
    .S1(net9636),
    .X(_03580_));
 sg13g2_a221oi_1 _24809_ (.B2(net8952),
    .C1(net9550),
    .B1(_03580_),
    .A1(net8815),
    .Y(_03581_),
    .A2(_03579_));
 sg13g2_o21ai_1 _24810_ (.B1(_03581_),
    .Y(_03582_),
    .A1(_03571_),
    .A2(_03578_));
 sg13g2_mux4_1 _24811_ (.S0(net9687),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][26] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][26] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][26] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][26] ),
    .S1(net9630),
    .X(_03583_));
 sg13g2_nor2_1 _24812_ (.A(net9578),
    .B(_03583_),
    .Y(_03584_));
 sg13g2_nor2_1 _24813_ (.A(net9104),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][26] ),
    .Y(_03585_));
 sg13g2_nor2_1 _24814_ (.A(net9691),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][26] ),
    .Y(_03586_));
 sg13g2_nor3_1 _24815_ (.A(net9638),
    .B(_03585_),
    .C(_03586_),
    .Y(_03587_));
 sg13g2_nor2_1 _24816_ (.A(net9691),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][26] ),
    .Y(_03588_));
 sg13g2_o21ai_1 _24817_ (.B1(net9630),
    .Y(_03589_),
    .A1(net9104),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][26] ));
 sg13g2_o21ai_1 _24818_ (.B1(net9578),
    .Y(_03590_),
    .A1(_03588_),
    .A2(_03589_));
 sg13g2_o21ai_1 _24819_ (.B1(net9561),
    .Y(_03591_),
    .A1(_03587_),
    .A2(_03590_));
 sg13g2_mux4_1 _24820_ (.S0(net9687),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][26] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][26] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][26] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][26] ),
    .S1(net9630),
    .X(_03592_));
 sg13g2_mux4_1 _24821_ (.S0(net9694),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][26] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][26] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][26] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][26] ),
    .S1(net9638),
    .X(_03593_));
 sg13g2_a22oi_1 _24822_ (.Y(_03594_),
    .B1(_03593_),
    .B2(net8952),
    .A2(_03592_),
    .A1(net8815));
 sg13g2_o21ai_1 _24823_ (.B1(_03594_),
    .Y(_03595_),
    .A1(_03584_),
    .A2(_03591_));
 sg13g2_o21ai_1 _24824_ (.B1(_03582_),
    .Y(_03596_),
    .A1(net9114),
    .A2(_03595_));
 sg13g2_nor2_1 _24825_ (.A(net8597),
    .B(_03596_),
    .Y(_00768_));
 sg13g2_nor2_1 _24826_ (.A(net9090),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][27] ),
    .Y(_03597_));
 sg13g2_nor2_1 _24827_ (.A(net9661),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][27] ),
    .Y(_03598_));
 sg13g2_nor3_1 _24828_ (.A(net9602),
    .B(_03597_),
    .C(_03598_),
    .Y(_03599_));
 sg13g2_nor2_1 _24829_ (.A(net9660),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][27] ),
    .Y(_03600_));
 sg13g2_o21ai_1 _24830_ (.B1(net9602),
    .Y(_03601_),
    .A1(net9090),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][27] ));
 sg13g2_o21ai_1 _24831_ (.B1(net9568),
    .Y(_03602_),
    .A1(_03600_),
    .A2(_03601_));
 sg13g2_mux4_1 _24832_ (.S0(net9661),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][27] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][27] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][27] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][27] ),
    .S1(net9603),
    .X(_03603_));
 sg13g2_nor2_1 _24833_ (.A(net9568),
    .B(_03603_),
    .Y(_03604_));
 sg13g2_o21ai_1 _24834_ (.B1(net9556),
    .Y(_03605_),
    .A1(_03599_),
    .A2(_03602_));
 sg13g2_mux4_1 _24835_ (.S0(net9660),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][27] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][27] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][27] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][27] ),
    .S1(net9603),
    .X(_03606_));
 sg13g2_mux4_1 _24836_ (.S0(net9661),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][27] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][27] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][27] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][27] ),
    .S1(net9603),
    .X(_03607_));
 sg13g2_a221oi_1 _24837_ (.B2(net8818),
    .C1(net9547),
    .B1(_03607_),
    .A1(net8949),
    .Y(_03608_),
    .A2(_03606_));
 sg13g2_o21ai_1 _24838_ (.B1(_03608_),
    .Y(_03609_),
    .A1(_03604_),
    .A2(_03605_));
 sg13g2_mux4_1 _24839_ (.S0(net9661),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][27] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][27] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][27] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][27] ),
    .S1(net9603),
    .X(_03610_));
 sg13g2_nor2_1 _24840_ (.A(net9090),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][27] ),
    .Y(_03611_));
 sg13g2_nor2_1 _24841_ (.A(net9661),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][27] ),
    .Y(_03612_));
 sg13g2_nor3_1 _24842_ (.A(net9603),
    .B(_03611_),
    .C(_03612_),
    .Y(_03613_));
 sg13g2_nor2_1 _24843_ (.A(net9661),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][27] ),
    .Y(_03614_));
 sg13g2_o21ai_1 _24844_ (.B1(net9603),
    .Y(_03615_),
    .A1(net9090),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][27] ));
 sg13g2_o21ai_1 _24845_ (.B1(net9568),
    .Y(_03616_),
    .A1(_03614_),
    .A2(_03615_));
 sg13g2_o21ai_1 _24846_ (.B1(net9556),
    .Y(_03617_),
    .A1(_03613_),
    .A2(_03616_));
 sg13g2_inv_1 _24847_ (.Y(_03618_),
    .A(_03617_));
 sg13g2_o21ai_1 _24848_ (.B1(_03618_),
    .Y(_03619_),
    .A1(net9568),
    .A2(_03610_));
 sg13g2_mux4_1 _24849_ (.S0(net9660),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][27] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][27] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][27] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][27] ),
    .S1(net9602),
    .X(_03620_));
 sg13g2_mux4_1 _24850_ (.S0(net9660),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][27] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][27] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][27] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][27] ),
    .S1(net9602),
    .X(_03621_));
 sg13g2_a221oi_1 _24851_ (.B2(net8811),
    .C1(net9112),
    .B1(_03621_),
    .A1(net8949),
    .Y(_03622_),
    .A2(_03620_));
 sg13g2_nand2_1 _24852_ (.Y(_03623_),
    .A(net8594),
    .B(_03609_));
 sg13g2_a21oi_1 _24853_ (.A1(_03619_),
    .A2(_03622_),
    .Y(_00769_),
    .B1(_03623_));
 sg13g2_nor2_1 _24854_ (.A(net9088),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][28] ),
    .Y(_03624_));
 sg13g2_nor2_1 _24855_ (.A(net9662),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][28] ),
    .Y(_03625_));
 sg13g2_nor3_1 _24856_ (.A(net9604),
    .B(_03624_),
    .C(_03625_),
    .Y(_03626_));
 sg13g2_nor2_1 _24857_ (.A(net9662),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][28] ),
    .Y(_03627_));
 sg13g2_o21ai_1 _24858_ (.B1(net9604),
    .Y(_03628_),
    .A1(net9088),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][28] ));
 sg13g2_o21ai_1 _24859_ (.B1(net9568),
    .Y(_03629_),
    .A1(_03627_),
    .A2(_03628_));
 sg13g2_a21oi_1 _24860_ (.A1(net9088),
    .A2(_10802_),
    .Y(_03630_),
    .B1(net9605));
 sg13g2_o21ai_1 _24861_ (.B1(_03630_),
    .Y(_03631_),
    .A1(net9088),
    .A2(net5575));
 sg13g2_mux2_1 _24862_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][28] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][28] ),
    .S(net9662),
    .X(_03632_));
 sg13g2_a21oi_1 _24863_ (.A1(net9605),
    .A2(_03632_),
    .Y(_03633_),
    .B1(net9568));
 sg13g2_a21oi_1 _24864_ (.A1(_03631_),
    .A2(_03633_),
    .Y(_03634_),
    .B1(_10462_));
 sg13g2_o21ai_1 _24865_ (.B1(_03634_),
    .Y(_03635_),
    .A1(_03626_),
    .A2(_03629_));
 sg13g2_mux4_1 _24866_ (.S0(net9662),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][28] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][28] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][28] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][28] ),
    .S1(net9604),
    .X(_03636_));
 sg13g2_mux4_1 _24867_ (.S0(net9662),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][28] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][28] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][28] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][28] ),
    .S1(net9604),
    .X(_03637_));
 sg13g2_a221oi_1 _24868_ (.B2(net8811),
    .C1(net9547),
    .B1(_03637_),
    .A1(net8948),
    .Y(_03638_),
    .A2(_03636_));
 sg13g2_a21oi_1 _24869_ (.A1(net9088),
    .A2(_10805_),
    .Y(_03639_),
    .B1(net9604));
 sg13g2_o21ai_1 _24870_ (.B1(_03639_),
    .Y(_03640_),
    .A1(net9088),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][28] ));
 sg13g2_nor2_1 _24871_ (.A(net9088),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][28] ),
    .Y(_03641_));
 sg13g2_a21oi_1 _24872_ (.A1(net9088),
    .A2(_10806_),
    .Y(_03642_),
    .B1(_03641_));
 sg13g2_a21oi_1 _24873_ (.A1(net9604),
    .A2(_03642_),
    .Y(_03643_),
    .B1(net9108));
 sg13g2_mux4_1 _24874_ (.S0(net9662),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][28] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][28] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][28] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][28] ),
    .S1(net9604),
    .X(_03644_));
 sg13g2_o21ai_1 _24875_ (.B1(net9555),
    .Y(_03645_),
    .A1(net9568),
    .A2(_03644_));
 sg13g2_a21oi_1 _24876_ (.A1(_03640_),
    .A2(_03643_),
    .Y(_03646_),
    .B1(_03645_));
 sg13g2_mux4_1 _24877_ (.S0(net9662),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][28] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][28] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][28] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][28] ),
    .S1(net9604),
    .X(_03647_));
 sg13g2_mux4_1 _24878_ (.S0(net9663),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][28] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][28] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][28] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][28] ),
    .S1(net9605),
    .X(_03648_));
 sg13g2_a221oi_1 _24879_ (.B2(net8811),
    .C1(_03646_),
    .B1(_03648_),
    .A1(net8948),
    .Y(_03649_),
    .A2(_03647_));
 sg13g2_a221oi_1 _24880_ (.B2(net9547),
    .C1(net8598),
    .B1(_03649_),
    .A1(net5576),
    .Y(_00770_),
    .A2(_03638_));
 sg13g2_nor2_1 _24881_ (.A(net9094),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][29] ),
    .Y(_03650_));
 sg13g2_nor2_1 _24882_ (.A(net9671),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][29] ),
    .Y(_03651_));
 sg13g2_nor3_1 _24883_ (.A(net9615),
    .B(_03650_),
    .C(_03651_),
    .Y(_03652_));
 sg13g2_nor2_1 _24884_ (.A(net9670),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][29] ),
    .Y(_03653_));
 sg13g2_o21ai_1 _24885_ (.B1(net9613),
    .Y(_03654_),
    .A1(net9093),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][29] ));
 sg13g2_o21ai_1 _24886_ (.B1(net9572),
    .Y(_03655_),
    .A1(_03653_),
    .A2(_03654_));
 sg13g2_a21oi_1 _24887_ (.A1(net9093),
    .A2(_10807_),
    .Y(_03656_),
    .B1(net9611));
 sg13g2_o21ai_1 _24888_ (.B1(_03656_),
    .Y(_03657_),
    .A1(net9093),
    .A2(net5579));
 sg13g2_mux2_1 _24889_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][29] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][29] ),
    .S(net9672),
    .X(_03658_));
 sg13g2_a21oi_1 _24890_ (.A1(net9615),
    .A2(_03658_),
    .Y(_03659_),
    .B1(net9572));
 sg13g2_a21oi_1 _24891_ (.A1(_03657_),
    .A2(_03659_),
    .Y(_03660_),
    .B1(_10462_));
 sg13g2_o21ai_1 _24892_ (.B1(_03660_),
    .Y(_03661_),
    .A1(_03652_),
    .A2(_03655_));
 sg13g2_mux4_1 _24893_ (.S0(net9670),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][29] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][29] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][29] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][29] ),
    .S1(net9613),
    .X(_03662_));
 sg13g2_mux4_1 _24894_ (.S0(net9670),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][29] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][29] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][29] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][29] ),
    .S1(net9613),
    .X(_03663_));
 sg13g2_a221oi_1 _24895_ (.B2(net8812),
    .C1(net9548),
    .B1(_03663_),
    .A1(net8950),
    .Y(_03664_),
    .A2(_03662_));
 sg13g2_mux4_1 _24896_ (.S0(net9672),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][29] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][29] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][29] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][29] ),
    .S1(net9615),
    .X(_03665_));
 sg13g2_nor2_1 _24897_ (.A(net9572),
    .B(_03665_),
    .Y(_03666_));
 sg13g2_nor2_1 _24898_ (.A(net9093),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][29] ),
    .Y(_03667_));
 sg13g2_nor2_1 _24899_ (.A(net9671),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][29] ),
    .Y(_03668_));
 sg13g2_nor3_1 _24900_ (.A(net9614),
    .B(_03667_),
    .C(_03668_),
    .Y(_03669_));
 sg13g2_nor2_1 _24901_ (.A(net9672),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][29] ),
    .Y(_03670_));
 sg13g2_o21ai_1 _24902_ (.B1(net9615),
    .Y(_03671_),
    .A1(net9094),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][29] ));
 sg13g2_o21ai_1 _24903_ (.B1(net9572),
    .Y(_03672_),
    .A1(_03670_),
    .A2(_03671_));
 sg13g2_o21ai_1 _24904_ (.B1(net9558),
    .Y(_03673_),
    .A1(_03669_),
    .A2(_03672_));
 sg13g2_mux4_1 _24905_ (.S0(net9672),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][29] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][29] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][29] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][29] ),
    .S1(net9614),
    .X(_03674_));
 sg13g2_mux4_1 _24906_ (.S0(net9670),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][29] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][29] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][29] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][29] ),
    .S1(net9615),
    .X(_03675_));
 sg13g2_a22oi_1 _24907_ (.Y(_03676_),
    .B1(_03675_),
    .B2(net8951),
    .A2(_03674_),
    .A1(net8812));
 sg13g2_o21ai_1 _24908_ (.B1(_03676_),
    .Y(_03677_),
    .A1(_03666_),
    .A2(_03673_));
 sg13g2_o21ai_1 _24909_ (.B1(net8595),
    .Y(_03678_),
    .A1(net9115),
    .A2(_03677_));
 sg13g2_a21oi_2 _24910_ (.B1(_03678_),
    .Y(_00771_),
    .A2(_03664_),
    .A1(_03661_));
 sg13g2_nor2_1 _24911_ (.A(net9087),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][30] ),
    .Y(_03679_));
 sg13g2_nor2_1 _24912_ (.A(net9658),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][30] ),
    .Y(_03680_));
 sg13g2_nor3_1 _24913_ (.A(net9600),
    .B(_03679_),
    .C(_03680_),
    .Y(_03681_));
 sg13g2_nor2_1 _24914_ (.A(net9660),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][30] ),
    .Y(_03682_));
 sg13g2_o21ai_1 _24915_ (.B1(net9602),
    .Y(_03683_),
    .A1(net9087),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][30] ));
 sg13g2_o21ai_1 _24916_ (.B1(net9569),
    .Y(_03684_),
    .A1(_03682_),
    .A2(_03683_));
 sg13g2_mux4_1 _24917_ (.S0(net9660),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][30] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][30] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][30] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][30] ),
    .S1(net9602),
    .X(_03685_));
 sg13g2_nor2_1 _24918_ (.A(net9569),
    .B(_03685_),
    .Y(_03686_));
 sg13g2_o21ai_1 _24919_ (.B1(net9555),
    .Y(_03687_),
    .A1(_03681_),
    .A2(_03684_));
 sg13g2_mux4_1 _24920_ (.S0(net9658),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][30] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][30] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][30] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][30] ),
    .S1(net9600),
    .X(_03688_));
 sg13g2_mux4_1 _24921_ (.S0(net9658),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][30] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][30] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][30] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][30] ),
    .S1(net9600),
    .X(_03689_));
 sg13g2_a221oi_1 _24922_ (.B2(net8811),
    .C1(net9547),
    .B1(_03689_),
    .A1(net8948),
    .Y(_03690_),
    .A2(_03688_));
 sg13g2_o21ai_1 _24923_ (.B1(_03690_),
    .Y(_03691_),
    .A1(_03686_),
    .A2(_03687_));
 sg13g2_mux4_1 _24924_ (.S0(net9657),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][30] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][30] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][30] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][30] ),
    .S1(net9599),
    .X(_03692_));
 sg13g2_nor2_1 _24925_ (.A(net9087),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][30] ),
    .Y(_03693_));
 sg13g2_nor2_1 _24926_ (.A(net9657),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][30] ),
    .Y(_03694_));
 sg13g2_nor3_1 _24927_ (.A(net9599),
    .B(_03693_),
    .C(_03694_),
    .Y(_03695_));
 sg13g2_nor2_1 _24928_ (.A(net9658),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][30] ),
    .Y(_03696_));
 sg13g2_o21ai_1 _24929_ (.B1(net9600),
    .Y(_03697_),
    .A1(net9087),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][30] ));
 sg13g2_o21ai_1 _24930_ (.B1(net9569),
    .Y(_03698_),
    .A1(_03696_),
    .A2(_03697_));
 sg13g2_o21ai_1 _24931_ (.B1(net9555),
    .Y(_03699_),
    .A1(_03695_),
    .A2(_03698_));
 sg13g2_inv_1 _24932_ (.Y(_03700_),
    .A(_03699_));
 sg13g2_o21ai_1 _24933_ (.B1(_03700_),
    .Y(_03701_),
    .A1(net9569),
    .A2(_03692_));
 sg13g2_mux4_1 _24934_ (.S0(net9657),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][30] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][30] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][30] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][30] ),
    .S1(net9599),
    .X(_03702_));
 sg13g2_mux4_1 _24935_ (.S0(net9657),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][30] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][30] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][30] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][30] ),
    .S1(net9599),
    .X(_03703_));
 sg13g2_a221oi_1 _24936_ (.B2(net8811),
    .C1(net9112),
    .B1(_03703_),
    .A1(net8948),
    .Y(_03704_),
    .A2(_03702_));
 sg13g2_nand2_1 _24937_ (.Y(_03705_),
    .A(net8594),
    .B(_03691_));
 sg13g2_a21oi_2 _24938_ (.B1(_03705_),
    .Y(_00772_),
    .A2(_03704_),
    .A1(_03701_));
 sg13g2_nor2_1 _24939_ (.A(net9083),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][31] ),
    .Y(_03706_));
 sg13g2_nor2_1 _24940_ (.A(net9656),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][31] ),
    .Y(_03707_));
 sg13g2_nor3_1 _24941_ (.A(net9595),
    .B(_03706_),
    .C(_03707_),
    .Y(_03708_));
 sg13g2_nor2_1 _24942_ (.A(net9656),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][31] ),
    .Y(_03709_));
 sg13g2_o21ai_1 _24943_ (.B1(net9597),
    .Y(_03710_),
    .A1(net9083),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][31] ));
 sg13g2_o21ai_1 _24944_ (.B1(net9570),
    .Y(_03711_),
    .A1(_03709_),
    .A2(_03710_));
 sg13g2_a21oi_1 _24945_ (.A1(net9083),
    .A2(_10814_),
    .Y(_03712_),
    .B1(net9595));
 sg13g2_o21ai_1 _24946_ (.B1(_03712_),
    .Y(_03713_),
    .A1(net9083),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][31] ));
 sg13g2_mux2_1 _24947_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][31] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][31] ),
    .S(net9653),
    .X(_03714_));
 sg13g2_a21oi_1 _24948_ (.A1(net9594),
    .A2(_03714_),
    .Y(_03715_),
    .B1(net9567));
 sg13g2_a21oi_1 _24949_ (.A1(_03713_),
    .A2(_03715_),
    .Y(_03716_),
    .B1(_10462_));
 sg13g2_o21ai_1 _24950_ (.B1(_03716_),
    .Y(_03717_),
    .A1(_03708_),
    .A2(_03711_));
 sg13g2_mux4_1 _24951_ (.S0(net9650),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][31] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][31] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][31] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][31] ),
    .S1(net9592),
    .X(_03718_));
 sg13g2_mux4_1 _24952_ (.S0(net9650),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][31] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][31] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][31] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][31] ),
    .S1(net9591),
    .X(_03719_));
 sg13g2_a221oi_1 _24953_ (.B2(net8810),
    .C1(net9547),
    .B1(_03719_),
    .A1(net8947),
    .Y(_03720_),
    .A2(_03718_));
 sg13g2_mux4_1 _24954_ (.S0(net9652),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][31] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][31] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][31] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][31] ),
    .S1(net9593),
    .X(_03721_));
 sg13g2_nor2_1 _24955_ (.A(net9566),
    .B(_03721_),
    .Y(_03722_));
 sg13g2_nor2_1 _24956_ (.A(net9084),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][31] ),
    .Y(_03723_));
 sg13g2_nor2_1 _24957_ (.A(net9655),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][31] ),
    .Y(_03724_));
 sg13g2_nor3_1 _24958_ (.A(net9596),
    .B(_03723_),
    .C(_03724_),
    .Y(_03725_));
 sg13g2_nor2_1 _24959_ (.A(net9654),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][31] ),
    .Y(_03726_));
 sg13g2_o21ai_1 _24960_ (.B1(net9595),
    .Y(_03727_),
    .A1(net9084),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][31] ));
 sg13g2_o21ai_1 _24961_ (.B1(net9567),
    .Y(_03728_),
    .A1(_03726_),
    .A2(_03727_));
 sg13g2_o21ai_1 _24962_ (.B1(net9554),
    .Y(_03729_),
    .A1(_03725_),
    .A2(_03728_));
 sg13g2_mux4_1 _24963_ (.S0(net9651),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][31] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][31] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][31] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][31] ),
    .S1(net9592),
    .X(_03730_));
 sg13g2_mux4_1 _24964_ (.S0(net9651),
    .A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][31] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][31] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][31] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][31] ),
    .S1(net9592),
    .X(_03731_));
 sg13g2_a22oi_1 _24965_ (.Y(_03732_),
    .B1(_03731_),
    .B2(net8947),
    .A2(_03730_),
    .A1(net8810));
 sg13g2_o21ai_1 _24966_ (.B1(_03732_),
    .Y(_03733_),
    .A1(_03722_),
    .A2(_03729_));
 sg13g2_o21ai_1 _24967_ (.B1(net8594),
    .Y(_03734_),
    .A1(net9111),
    .A2(_03733_));
 sg13g2_a21oi_2 _24968_ (.B1(_03734_),
    .Y(_00773_),
    .A2(_03720_),
    .A1(_03717_));
 sg13g2_o21ai_1 _24969_ (.B1(net7389),
    .Y(_03735_),
    .A1(_00241_),
    .A2(net8684));
 sg13g2_nor3_1 _24970_ (.A(net9257),
    .B(net4704),
    .C(net8683),
    .Y(_03736_));
 sg13g2_o21ai_1 _24971_ (.B1(net9343),
    .Y(_03737_),
    .A1(_03735_),
    .A2(_03736_));
 sg13g2_a21oi_1 _24972_ (.A1(_10557_),
    .A2(_03735_),
    .Y(_00774_),
    .B1(_03737_));
 sg13g2_nor2_1 _24973_ (.A(_10556_),
    .B(_10557_),
    .Y(_03738_));
 sg13g2_o21ai_1 _24974_ (.B1(_00241_),
    .Y(_03739_),
    .A1(_11847_),
    .A2(_03738_));
 sg13g2_o21ai_1 _24975_ (.B1(_14278_),
    .Y(_03740_),
    .A1(net8683),
    .A2(_03739_));
 sg13g2_o21ai_1 _24976_ (.B1(net9341),
    .Y(_03741_),
    .A1(_03735_),
    .A2(_03740_));
 sg13g2_a21oi_1 _24977_ (.A1(_10556_),
    .A2(_03735_),
    .Y(_00775_),
    .B1(_03741_));
 sg13g2_nor3_2 _24978_ (.A(net9711),
    .B(\soc_I.kianv_I.Instr[9] ),
    .C(_14369_),
    .Y(_03742_));
 sg13g2_nand2_2 _24979_ (.Y(_03743_),
    .A(_14199_),
    .B(_03742_));
 sg13g2_nand2_1 _24980_ (.Y(_03744_),
    .A(net3055),
    .B(net7891));
 sg13g2_o21ai_1 _24981_ (.B1(_03744_),
    .Y(_00776_),
    .A1(net7486),
    .A2(net7891));
 sg13g2_nand2_1 _24982_ (.Y(_03745_),
    .A(net3748),
    .B(net7889));
 sg13g2_o21ai_1 _24983_ (.B1(_03745_),
    .Y(_00777_),
    .A1(net7666),
    .A2(net7889));
 sg13g2_nand2_1 _24984_ (.Y(_03746_),
    .A(net3292),
    .B(net7891));
 sg13g2_o21ai_1 _24985_ (.B1(_03746_),
    .Y(_00778_),
    .A1(net7615),
    .A2(net7891));
 sg13g2_nand2_1 _24986_ (.Y(_03747_),
    .A(net3510),
    .B(net7892));
 sg13g2_o21ai_1 _24987_ (.B1(_03747_),
    .Y(_00779_),
    .A1(net7609),
    .A2(net7892));
 sg13g2_nand2_1 _24988_ (.Y(_03748_),
    .A(net4187),
    .B(net7888));
 sg13g2_o21ai_1 _24989_ (.B1(_03748_),
    .Y(_00780_),
    .A1(net7588),
    .A2(net7888));
 sg13g2_nand2_1 _24990_ (.Y(_03749_),
    .A(net3893),
    .B(net7887));
 sg13g2_o21ai_1 _24991_ (.B1(_03749_),
    .Y(_00781_),
    .A1(net7601),
    .A2(net7887));
 sg13g2_nand2_1 _24992_ (.Y(_03750_),
    .A(net2994),
    .B(net7890));
 sg13g2_o21ai_1 _24993_ (.B1(_03750_),
    .Y(_00782_),
    .A1(net7593),
    .A2(net7890));
 sg13g2_nand2_1 _24994_ (.Y(_03751_),
    .A(net3392),
    .B(net7884));
 sg13g2_o21ai_1 _24995_ (.B1(_03751_),
    .Y(_00783_),
    .A1(net7606),
    .A2(net7884));
 sg13g2_nand2_1 _24996_ (.Y(_03752_),
    .A(net2972),
    .B(net7887));
 sg13g2_o21ai_1 _24997_ (.B1(_03752_),
    .Y(_00784_),
    .A1(net7557),
    .A2(net7887));
 sg13g2_nand2_1 _24998_ (.Y(_03753_),
    .A(net2978),
    .B(net7889));
 sg13g2_o21ai_1 _24999_ (.B1(_03753_),
    .Y(_00785_),
    .A1(net7576),
    .A2(net7889));
 sg13g2_nand2_1 _25000_ (.Y(_03754_),
    .A(net2886),
    .B(net7890));
 sg13g2_o21ai_1 _25001_ (.B1(_03754_),
    .Y(_00786_),
    .A1(net7546),
    .A2(net7890));
 sg13g2_nand2_1 _25002_ (.Y(_03755_),
    .A(net3669),
    .B(net7883));
 sg13g2_o21ai_1 _25003_ (.B1(_03755_),
    .Y(_00787_),
    .A1(net7571),
    .A2(net7883));
 sg13g2_nand2_1 _25004_ (.Y(_03756_),
    .A(net3458),
    .B(net7890));
 sg13g2_o21ai_1 _25005_ (.B1(_03756_),
    .Y(_00788_),
    .A1(net7541),
    .A2(net7891));
 sg13g2_nand2_1 _25006_ (.Y(_03757_),
    .A(net3387),
    .B(net7890));
 sg13g2_o21ai_1 _25007_ (.B1(_03757_),
    .Y(_00789_),
    .A1(net7556),
    .A2(net7890));
 sg13g2_nand2_1 _25008_ (.Y(_03758_),
    .A(net3155),
    .B(net7885));
 sg13g2_o21ai_1 _25009_ (.B1(_03758_),
    .Y(_00790_),
    .A1(net7580),
    .A2(net7885));
 sg13g2_nand2_1 _25010_ (.Y(_03759_),
    .A(net3545),
    .B(net7884));
 sg13g2_o21ai_1 _25011_ (.B1(_03759_),
    .Y(_00791_),
    .A1(net7566),
    .A2(net7884));
 sg13g2_nand2_1 _25012_ (.Y(_03760_),
    .A(net4200),
    .B(net7883));
 sg13g2_o21ai_1 _25013_ (.B1(_03760_),
    .Y(_00792_),
    .A1(net7526),
    .A2(net7883));
 sg13g2_nand2_1 _25014_ (.Y(_03761_),
    .A(net3579),
    .B(net7883));
 sg13g2_o21ai_1 _25015_ (.B1(_03761_),
    .Y(_00793_),
    .A1(net7537),
    .A2(net7883));
 sg13g2_nand2_1 _25016_ (.Y(_03762_),
    .A(net2838),
    .B(net7885));
 sg13g2_o21ai_1 _25017_ (.B1(_03762_),
    .Y(_00794_),
    .A1(net7532),
    .A2(net7885));
 sg13g2_nand2_1 _25018_ (.Y(_03763_),
    .A(net3680),
    .B(net7885));
 sg13g2_o21ai_1 _25019_ (.B1(_03763_),
    .Y(_00795_),
    .A1(net7518),
    .A2(net7885));
 sg13g2_nand2_1 _25020_ (.Y(_03764_),
    .A(net3373),
    .B(net7888));
 sg13g2_o21ai_1 _25021_ (.B1(_03764_),
    .Y(_00796_),
    .A1(net7504),
    .A2(net7888));
 sg13g2_nand2_1 _25022_ (.Y(_03765_),
    .A(net3878),
    .B(_03743_));
 sg13g2_o21ai_1 _25023_ (.B1(_03765_),
    .Y(_00797_),
    .A1(net7512),
    .A2(net7886));
 sg13g2_nand2_1 _25024_ (.Y(_03766_),
    .A(net3054),
    .B(net7889));
 sg13g2_o21ai_1 _25025_ (.B1(_03766_),
    .Y(_00798_),
    .A1(net7494),
    .A2(net7889));
 sg13g2_nand2_1 _25026_ (.Y(_03767_),
    .A(net4067),
    .B(net7884));
 sg13g2_o21ai_1 _25027_ (.B1(_03767_),
    .Y(_00799_),
    .A1(net7503),
    .A2(net7884));
 sg13g2_nand2_1 _25028_ (.Y(_03768_),
    .A(net3557),
    .B(net7887));
 sg13g2_o21ai_1 _25029_ (.B1(_03768_),
    .Y(_00800_),
    .A1(net7646),
    .A2(net7887));
 sg13g2_nand2_1 _25030_ (.Y(_03769_),
    .A(net3830),
    .B(net7891));
 sg13g2_o21ai_1 _25031_ (.B1(_03769_),
    .Y(_00801_),
    .A1(net7649),
    .A2(net7891));
 sg13g2_nand2_1 _25032_ (.Y(_03770_),
    .A(net3281),
    .B(net7889));
 sg13g2_o21ai_1 _25033_ (.B1(_03770_),
    .Y(_00802_),
    .A1(net7656),
    .A2(net7889));
 sg13g2_nand2_1 _25034_ (.Y(_03771_),
    .A(net3152),
    .B(net7886));
 sg13g2_o21ai_1 _25035_ (.B1(_03771_),
    .Y(_00803_),
    .A1(net7661),
    .A2(net7886));
 sg13g2_nand2_1 _25036_ (.Y(_03772_),
    .A(net3182),
    .B(net7886));
 sg13g2_o21ai_1 _25037_ (.B1(_03772_),
    .Y(_00804_),
    .A1(net7638),
    .A2(net7886));
 sg13g2_nand2_1 _25038_ (.Y(_03773_),
    .A(net3115),
    .B(net7887));
 sg13g2_o21ai_1 _25039_ (.B1(_03773_),
    .Y(_00805_),
    .A1(net7628),
    .A2(net7887));
 sg13g2_nand2_1 _25040_ (.Y(_03774_),
    .A(net3722),
    .B(net7886));
 sg13g2_o21ai_1 _25041_ (.B1(_03774_),
    .Y(_00806_),
    .A1(net7620),
    .A2(net7886));
 sg13g2_nand2_1 _25042_ (.Y(_03775_),
    .A(net3002),
    .B(net7883));
 sg13g2_o21ai_1 _25043_ (.B1(_03775_),
    .Y(_00807_),
    .A1(net7630),
    .A2(net7883));
 sg13g2_nand2_2 _25044_ (.Y(_03776_),
    .A(_12607_),
    .B(_14302_));
 sg13g2_nand2_1 _25045_ (.Y(_03777_),
    .A(net3203),
    .B(net8135));
 sg13g2_o21ai_1 _25046_ (.B1(_03777_),
    .Y(_00808_),
    .A1(net7487),
    .A2(net8135));
 sg13g2_nand2_1 _25047_ (.Y(_03778_),
    .A(net2940),
    .B(net8135));
 sg13g2_o21ai_1 _25048_ (.B1(_03778_),
    .Y(_00809_),
    .A1(net7663),
    .A2(net8135));
 sg13g2_nand2_1 _25049_ (.Y(_03779_),
    .A(net3731),
    .B(net8135));
 sg13g2_o21ai_1 _25050_ (.B1(_03779_),
    .Y(_00810_),
    .A1(net7617),
    .A2(net8135));
 sg13g2_nand2_1 _25051_ (.Y(_03780_),
    .A(net3051),
    .B(net8133));
 sg13g2_o21ai_1 _25052_ (.B1(_03780_),
    .Y(_00811_),
    .A1(net7609),
    .A2(net8133));
 sg13g2_nand2_1 _25053_ (.Y(_03781_),
    .A(net2812),
    .B(net8131));
 sg13g2_o21ai_1 _25054_ (.B1(_03781_),
    .Y(_00812_),
    .A1(net7586),
    .A2(net8131));
 sg13g2_nand2_1 _25055_ (.Y(_03782_),
    .A(net3225),
    .B(net8130));
 sg13g2_o21ai_1 _25056_ (.B1(_03782_),
    .Y(_00813_),
    .A1(net7600),
    .A2(net8130));
 sg13g2_nand2_1 _25057_ (.Y(_03783_),
    .A(net3274),
    .B(net8132));
 sg13g2_o21ai_1 _25058_ (.B1(_03783_),
    .Y(_00814_),
    .A1(net7595),
    .A2(net8132));
 sg13g2_nand2_1 _25059_ (.Y(_03784_),
    .A(net3245),
    .B(net8125));
 sg13g2_o21ai_1 _25060_ (.B1(_03784_),
    .Y(_00815_),
    .A1(net7603),
    .A2(net8125));
 sg13g2_nand2_1 _25061_ (.Y(_03785_),
    .A(net3127),
    .B(net8131));
 sg13g2_o21ai_1 _25062_ (.B1(_03785_),
    .Y(_00816_),
    .A1(net7562),
    .A2(net8131));
 sg13g2_nand2_1 _25063_ (.Y(_03786_),
    .A(net2878),
    .B(net8134));
 sg13g2_o21ai_1 _25064_ (.B1(_03786_),
    .Y(_00817_),
    .A1(net7577),
    .A2(net8134));
 sg13g2_nand2_1 _25065_ (.Y(_03787_),
    .A(net2985),
    .B(net8132));
 sg13g2_o21ai_1 _25066_ (.B1(_03787_),
    .Y(_00818_),
    .A1(net7548),
    .A2(net8132));
 sg13g2_nand2_1 _25067_ (.Y(_03788_),
    .A(net2873),
    .B(net8125));
 sg13g2_o21ai_1 _25068_ (.B1(_03788_),
    .Y(_00819_),
    .A1(net7568),
    .A2(net8125));
 sg13g2_nand2_1 _25069_ (.Y(_03789_),
    .A(net2930),
    .B(net8132));
 sg13g2_o21ai_1 _25070_ (.B1(_03789_),
    .Y(_00820_),
    .A1(net7543),
    .A2(net8132));
 sg13g2_nand2_1 _25071_ (.Y(_03790_),
    .A(net3398),
    .B(net8134));
 sg13g2_o21ai_1 _25072_ (.B1(_03790_),
    .Y(_00821_),
    .A1(net7552),
    .A2(net8134));
 sg13g2_nand2_1 _25073_ (.Y(_03791_),
    .A(net2778),
    .B(net8129));
 sg13g2_o21ai_1 _25074_ (.B1(_03791_),
    .Y(_00822_),
    .A1(net7585),
    .A2(net8129));
 sg13g2_nand2_1 _25075_ (.Y(_03792_),
    .A(net3661),
    .B(net8126));
 sg13g2_o21ai_1 _25076_ (.B1(_03792_),
    .Y(_00823_),
    .A1(net7564),
    .A2(net8126));
 sg13g2_nand2_1 _25077_ (.Y(_03793_),
    .A(net3920),
    .B(net8125));
 sg13g2_o21ai_1 _25078_ (.B1(_03793_),
    .Y(_00824_),
    .A1(net7522),
    .A2(net8125));
 sg13g2_nand2_1 _25079_ (.Y(_03794_),
    .A(net3518),
    .B(net8125));
 sg13g2_o21ai_1 _25080_ (.B1(_03794_),
    .Y(_00825_),
    .A1(net7534),
    .A2(net8125));
 sg13g2_nand2_1 _25081_ (.Y(_03795_),
    .A(net3524),
    .B(net8126));
 sg13g2_o21ai_1 _25082_ (.B1(_03795_),
    .Y(_00826_),
    .A1(net7533),
    .A2(net8126));
 sg13g2_nand2_1 _25083_ (.Y(_03796_),
    .A(net3169),
    .B(net8128));
 sg13g2_o21ai_1 _25084_ (.B1(_03796_),
    .Y(_00827_),
    .A1(net7518),
    .A2(net8128));
 sg13g2_nand2_1 _25085_ (.Y(_03797_),
    .A(net3408),
    .B(net8131));
 sg13g2_o21ai_1 _25086_ (.B1(_03797_),
    .Y(_00828_),
    .A1(net7509),
    .A2(net8131));
 sg13g2_nand2_1 _25087_ (.Y(_03798_),
    .A(net3117),
    .B(net8130));
 sg13g2_o21ai_1 _25088_ (.B1(_03798_),
    .Y(_00829_),
    .A1(net7513),
    .A2(net8130));
 sg13g2_nand2_1 _25089_ (.Y(_03799_),
    .A(net2836),
    .B(net8133));
 sg13g2_o21ai_1 _25090_ (.B1(_03799_),
    .Y(_00830_),
    .A1(net7496),
    .A2(net8133));
 sg13g2_nand2_1 _25091_ (.Y(_03800_),
    .A(net3171),
    .B(net8126));
 sg13g2_o21ai_1 _25092_ (.B1(_03800_),
    .Y(_00831_),
    .A1(net7499),
    .A2(net8126));
 sg13g2_nand2_1 _25093_ (.Y(_03801_),
    .A(net3013),
    .B(net8130));
 sg13g2_o21ai_1 _25094_ (.B1(_03801_),
    .Y(_00832_),
    .A1(net7644),
    .A2(net8130));
 sg13g2_nand2_1 _25095_ (.Y(_03802_),
    .A(net3237),
    .B(net8135));
 sg13g2_o21ai_1 _25096_ (.B1(_03802_),
    .Y(_00833_),
    .A1(net7650),
    .A2(net8135));
 sg13g2_nand2_1 _25097_ (.Y(_03803_),
    .A(net2884),
    .B(net8132));
 sg13g2_o21ai_1 _25098_ (.B1(_03803_),
    .Y(_00834_),
    .A1(net7655),
    .A2(net8132));
 sg13g2_nand2_1 _25099_ (.Y(_03804_),
    .A(net2965),
    .B(net8128));
 sg13g2_o21ai_1 _25100_ (.B1(_03804_),
    .Y(_00835_),
    .A1(net7658),
    .A2(net8128));
 sg13g2_nand2_1 _25101_ (.Y(_03805_),
    .A(net2824),
    .B(net8128));
 sg13g2_o21ai_1 _25102_ (.B1(_03805_),
    .Y(_00836_),
    .A1(net7638),
    .A2(net8128));
 sg13g2_nand2_1 _25103_ (.Y(_03806_),
    .A(net3449),
    .B(net8130));
 sg13g2_o21ai_1 _25104_ (.B1(_03806_),
    .Y(_00837_),
    .A1(net7629),
    .A2(net8130));
 sg13g2_nand2_1 _25105_ (.Y(_03807_),
    .A(net3184),
    .B(net8128));
 sg13g2_o21ai_1 _25106_ (.B1(_03807_),
    .Y(_00838_),
    .A1(net7621),
    .A2(net8128));
 sg13g2_nand2_1 _25107_ (.Y(_03808_),
    .A(net3811),
    .B(net8127));
 sg13g2_o21ai_1 _25108_ (.B1(_03808_),
    .Y(_00839_),
    .A1(net7634),
    .A2(net8127));
 sg13g2_nand4_1 _25109_ (.B(net9203),
    .C(net8975),
    .A(net9202),
    .Y(_03809_),
    .D(net8974));
 sg13g2_nor2b_2 _25110_ (.A(net9202),
    .B_N(net9203),
    .Y(_03810_));
 sg13g2_nand2b_2 _25111_ (.Y(_03811_),
    .B(net9203),
    .A_N(net9202));
 sg13g2_nand2_1 _25112_ (.Y(_03812_),
    .A(_13830_),
    .B(_03810_));
 sg13g2_and2_1 _25113_ (.A(_03809_),
    .B(_03812_),
    .X(_03813_));
 sg13g2_o21ai_1 _25114_ (.B1(_03810_),
    .Y(_03814_),
    .A1(_10842_),
    .A2(_10862_));
 sg13g2_and2_1 _25115_ (.A(_03813_),
    .B(_03814_),
    .X(_03815_));
 sg13g2_nand3_1 _25116_ (.B(net8973),
    .C(_03810_),
    .A(net8975),
    .Y(_03816_));
 sg13g2_nand2_1 _25117_ (.Y(_03817_),
    .A(_03815_),
    .B(_03816_));
 sg13g2_nor2_2 _25118_ (.A(_10866_),
    .B(_03811_),
    .Y(_03818_));
 sg13g2_nor3_2 _25119_ (.A(_10849_),
    .B(_10861_),
    .C(_03811_),
    .Y(_03819_));
 sg13g2_nor2_2 _25120_ (.A(_11731_),
    .B(_03811_),
    .Y(_03820_));
 sg13g2_nand3_1 _25121_ (.B(net8975),
    .C(_03810_),
    .A(_10832_),
    .Y(_03821_));
 sg13g2_nor4_1 _25122_ (.A(net8491),
    .B(net8673),
    .C(_03819_),
    .D(_03820_),
    .Y(_03822_));
 sg13g2_or4_1 _25123_ (.A(net8491),
    .B(net8673),
    .C(_03819_),
    .D(_03820_),
    .X(_03823_));
 sg13g2_nor2b_1 _25124_ (.A(_10921_),
    .B_N(_13290_),
    .Y(_03824_));
 sg13g2_nand2_2 _25125_ (.Y(_03825_),
    .A(_10874_),
    .B(_10923_));
 sg13g2_nand2_1 _25126_ (.Y(_03826_),
    .A(_10878_),
    .B(_13290_));
 sg13g2_nor2b_1 _25127_ (.A(_03826_),
    .B_N(_10917_),
    .Y(_03827_));
 sg13g2_nand2_1 _25128_ (.Y(_03828_),
    .A(_03824_),
    .B(_03825_));
 sg13g2_a21oi_1 _25129_ (.A1(_00188_),
    .A2(net8962),
    .Y(_03829_),
    .B1(_03824_));
 sg13g2_nand3_1 _25130_ (.B(net9703),
    .C(_03829_),
    .A(net9698),
    .Y(_03830_));
 sg13g2_and2_1 _25131_ (.A(_03828_),
    .B(_03830_),
    .X(_03831_));
 sg13g2_nand2_2 _25132_ (.Y(_03832_),
    .A(_03828_),
    .B(_03830_));
 sg13g2_nand2b_1 _25133_ (.Y(_03833_),
    .B(_03827_),
    .A_N(_03824_));
 sg13g2_and2_1 _25134_ (.A(_03825_),
    .B(_03833_),
    .X(_03834_));
 sg13g2_nand2_2 _25135_ (.Y(_03835_),
    .A(_03825_),
    .B(_03833_));
 sg13g2_nor2_1 _25136_ (.A(net9659),
    .B(net8343),
    .Y(_03836_));
 sg13g2_a21oi_1 _25137_ (.A1(_11185_),
    .A2(net8343),
    .Y(_03837_),
    .B1(_03836_));
 sg13g2_nor3_1 _25138_ (.A(_03825_),
    .B(_03827_),
    .C(_03829_),
    .Y(_03838_));
 sg13g2_a221oi_1 _25139_ (.B2(_03829_),
    .C1(_03838_),
    .B1(_03826_),
    .A1(_03824_),
    .Y(_03839_),
    .A2(_03825_));
 sg13g2_nor2_1 _25140_ (.A(_03837_),
    .B(net8334),
    .Y(_03840_));
 sg13g2_a22oi_1 _25141_ (.Y(_03841_),
    .B1(_03840_),
    .B2(\soc_I.kianv_I.datapath_unit_I.CSRData[0] ),
    .A2(_03837_),
    .A1(net8346));
 sg13g2_nor2_1 _25142_ (.A(net8356),
    .B(_03841_),
    .Y(_03842_));
 sg13g2_a21oi_1 _25143_ (.A1(_10919_),
    .A2(_11002_),
    .Y(_03843_),
    .B1(net8597));
 sg13g2_o21ai_1 _25144_ (.B1(_10969_),
    .Y(_03844_),
    .A1(_10918_),
    .A2(_03843_));
 sg13g2_inv_1 _25145_ (.Y(_03845_),
    .A(_03844_));
 sg13g2_nand3_1 _25146_ (.B(_00239_),
    .C(net8711),
    .A(net9427),
    .Y(_03846_));
 sg13g2_o21ai_1 _25147_ (.B1(_00240_),
    .Y(_03847_),
    .A1(net9427),
    .A2(_00239_));
 sg13g2_o21ai_1 _25148_ (.B1(_03846_),
    .Y(_03848_),
    .A1(_11209_),
    .A2(_03847_));
 sg13g2_a21o_1 _25149_ (.A2(_03845_),
    .A1(_12580_),
    .B1(_03848_),
    .X(_03849_));
 sg13g2_nor2_2 _25150_ (.A(_03844_),
    .B(_03849_),
    .Y(_03850_));
 sg13g2_and2_2 _25151_ (.A(net7796),
    .B(net7993),
    .X(_03851_));
 sg13g2_nand2_2 _25152_ (.Y(_03852_),
    .A(net7797),
    .B(net7992));
 sg13g2_nor2_2 _25153_ (.A(net8354),
    .B(_03851_),
    .Y(_03853_));
 sg13g2_nand2_2 _25154_ (.Y(_03854_),
    .A(net8366),
    .B(net7747));
 sg13g2_a21oi_1 _25155_ (.A1(\soc_I.kianv_I.Instr[0] ),
    .A2(net8673),
    .Y(_03855_),
    .B1(net8488));
 sg13g2_a21oi_1 _25156_ (.A1(_10496_),
    .A2(net8488),
    .Y(_03856_),
    .B1(_03855_));
 sg13g2_nor3_1 _25157_ (.A(_03842_),
    .B(net7705),
    .C(_03856_),
    .Y(_03857_));
 sg13g2_o21ai_1 _25158_ (.B1(net9391),
    .Y(_03858_),
    .A1(net4451),
    .A2(net7704));
 sg13g2_nor2_1 _25159_ (.A(_03857_),
    .B(_03858_),
    .Y(_00840_));
 sg13g2_nor2_1 _25160_ (.A(net8300),
    .B(net8340),
    .Y(_03859_));
 sg13g2_a21oi_1 _25161_ (.A1(_00293_),
    .A2(net8339),
    .Y(_03860_),
    .B1(_03859_));
 sg13g2_nor2_1 _25162_ (.A(net8334),
    .B(_03860_),
    .Y(_03861_));
 sg13g2_a22oi_1 _25163_ (.Y(_03862_),
    .B1(_03861_),
    .B2(\soc_I.kianv_I.datapath_unit_I.CSRData[1] ),
    .A2(_03860_),
    .A1(net8346));
 sg13g2_nor2_1 _25164_ (.A(net8356),
    .B(_03862_),
    .Y(_03863_));
 sg13g2_a21oi_1 _25165_ (.A1(\soc_I.kianv_I.Instr[1] ),
    .A2(net8673),
    .Y(_03864_),
    .B1(net8489));
 sg13g2_a21oi_1 _25166_ (.A1(_10495_),
    .A2(net8489),
    .Y(_03865_),
    .B1(_03864_));
 sg13g2_a221oi_1 _25167_ (.B2(_03851_),
    .C1(_03865_),
    .B1(_03863_),
    .A1(net5218),
    .Y(_03866_),
    .A2(net7705));
 sg13g2_nor2_1 _25168_ (.A(net9038),
    .B(_03866_),
    .Y(_00841_));
 sg13g2_nand2_1 _25169_ (.Y(_03867_),
    .A(_00294_),
    .B(net8341));
 sg13g2_o21ai_1 _25170_ (.B1(_03867_),
    .Y(_03868_),
    .A1(_11144_),
    .A2(net8341));
 sg13g2_nor2_1 _25171_ (.A(_03832_),
    .B(_03868_),
    .Y(_03869_));
 sg13g2_nor2b_1 _25172_ (.A(net8337),
    .B_N(_03868_),
    .Y(_03870_));
 sg13g2_a21oi_2 _25173_ (.B1(_03869_),
    .Y(_03871_),
    .A2(_03870_),
    .A1(\soc_I.kianv_I.datapath_unit_I.CSRData[2] ));
 sg13g2_nor2_1 _25174_ (.A(net8354),
    .B(_03871_),
    .Y(_03872_));
 sg13g2_a21oi_1 _25175_ (.A1(\soc_I.kianv_I.Instr[2] ),
    .A2(net8673),
    .Y(_03873_),
    .B1(net8489));
 sg13g2_a21oi_1 _25176_ (.A1(_10494_),
    .A2(net8488),
    .Y(_03874_),
    .B1(_03873_));
 sg13g2_a221oi_1 _25177_ (.B2(_03851_),
    .C1(_03874_),
    .B1(_03872_),
    .A1(net5077),
    .Y(_03875_),
    .A2(net7705));
 sg13g2_nor2_1 _25178_ (.A(net9038),
    .B(_03875_),
    .Y(_00842_));
 sg13g2_nand2_1 _25179_ (.Y(_03876_),
    .A(_00295_),
    .B(net8339));
 sg13g2_o21ai_1 _25180_ (.B1(_03876_),
    .Y(_03877_),
    .A1(_11132_),
    .A2(net8339));
 sg13g2_nor2_1 _25181_ (.A(_03832_),
    .B(_03877_),
    .Y(_03878_));
 sg13g2_nor2b_1 _25182_ (.A(net8334),
    .B_N(_03877_),
    .Y(_03879_));
 sg13g2_a21oi_2 _25183_ (.B1(_03878_),
    .Y(_03880_),
    .A2(_03879_),
    .A1(\soc_I.kianv_I.datapath_unit_I.CSRData[3] ));
 sg13g2_nor2_1 _25184_ (.A(net8356),
    .B(_03880_),
    .Y(_03881_));
 sg13g2_a21oi_1 _25185_ (.A1(\soc_I.kianv_I.Instr[3] ),
    .A2(net8673),
    .Y(_03882_),
    .B1(net8489));
 sg13g2_a21oi_1 _25186_ (.A1(_10493_),
    .A2(net8489),
    .Y(_03883_),
    .B1(_03882_));
 sg13g2_nor3_1 _25187_ (.A(net7705),
    .B(_03881_),
    .C(_03883_),
    .Y(_03884_));
 sg13g2_o21ai_1 _25188_ (.B1(net9378),
    .Y(_03885_),
    .A1(net4660),
    .A2(net7704));
 sg13g2_nor2_1 _25189_ (.A(_03884_),
    .B(_03885_),
    .Y(_00843_));
 sg13g2_nor2_1 _25190_ (.A(_11118_),
    .B(net8341),
    .Y(_03886_));
 sg13g2_a21oi_1 _25191_ (.A1(_00296_),
    .A2(net8341),
    .Y(_03887_),
    .B1(_03886_));
 sg13g2_nor2_1 _25192_ (.A(net8337),
    .B(_03887_),
    .Y(_03888_));
 sg13g2_a22oi_1 _25193_ (.Y(_03889_),
    .B1(_03888_),
    .B2(\soc_I.kianv_I.datapath_unit_I.CSRData[4] ),
    .A2(_03887_),
    .A1(net8347));
 sg13g2_nor2_1 _25194_ (.A(net8354),
    .B(_03889_),
    .Y(_03890_));
 sg13g2_a21oi_1 _25195_ (.A1(net9715),
    .A2(_03818_),
    .Y(_03891_),
    .B1(net8489));
 sg13g2_a21oi_1 _25196_ (.A1(_10492_),
    .A2(net8488),
    .Y(_03892_),
    .B1(_03891_));
 sg13g2_a221oi_1 _25197_ (.B2(_03851_),
    .C1(_03892_),
    .B1(_03890_),
    .A1(net5059),
    .Y(_03893_),
    .A2(net7705));
 sg13g2_nor2_1 _25198_ (.A(net9046),
    .B(_03893_),
    .Y(_00844_));
 sg13g2_and2_1 _25199_ (.A(net8306),
    .B(net8344),
    .X(_03894_));
 sg13g2_nor2_1 _25200_ (.A(net8336),
    .B(_03894_),
    .Y(_03895_));
 sg13g2_a22oi_1 _25201_ (.Y(_03896_),
    .B1(_03895_),
    .B2(\soc_I.kianv_I.datapath_unit_I.CSRData[5] ),
    .A2(_03894_),
    .A1(net8346));
 sg13g2_nor2_1 _25202_ (.A(net8356),
    .B(_03896_),
    .Y(_03897_));
 sg13g2_a21oi_1 _25203_ (.A1(net9714),
    .A2(net8673),
    .Y(_03898_),
    .B1(net8488));
 sg13g2_a21oi_1 _25204_ (.A1(_10491_),
    .A2(net8488),
    .Y(_03899_),
    .B1(_03898_));
 sg13g2_nor3_1 _25205_ (.A(net7705),
    .B(_03897_),
    .C(_03899_),
    .Y(_03900_));
 sg13g2_o21ai_1 _25206_ (.B1(net9376),
    .Y(_03901_),
    .A1(net4562),
    .A2(net7704));
 sg13g2_nor2_1 _25207_ (.A(_03900_),
    .B(_03901_),
    .Y(_00845_));
 sg13g2_nor2_2 _25208_ (.A(_11097_),
    .B(net8342),
    .Y(_03902_));
 sg13g2_nor2_1 _25209_ (.A(net8337),
    .B(_03902_),
    .Y(_03903_));
 sg13g2_a22oi_1 _25210_ (.Y(_03904_),
    .B1(_03903_),
    .B2(\soc_I.kianv_I.datapath_unit_I.CSRData[6] ),
    .A2(_03902_),
    .A1(net8347));
 sg13g2_nor2_1 _25211_ (.A(net8354),
    .B(_03904_),
    .Y(_03905_));
 sg13g2_a21oi_1 _25212_ (.A1(net9712),
    .A2(_03818_),
    .Y(_03906_),
    .B1(net8488));
 sg13g2_a21oi_1 _25213_ (.A1(_10490_),
    .A2(net8488),
    .Y(_03907_),
    .B1(_03906_));
 sg13g2_a221oi_1 _25214_ (.B2(_03851_),
    .C1(_03907_),
    .B1(_03905_),
    .A1(net5124),
    .Y(_03908_),
    .A2(net7705));
 sg13g2_nor2_1 _25215_ (.A(net9046),
    .B(_03908_),
    .Y(_00846_));
 sg13g2_nand3_1 _25216_ (.B(net8346),
    .C(net8343),
    .A(_11086_),
    .Y(_03909_));
 sg13g2_a21oi_1 _25217_ (.A1(_11086_),
    .A2(net8343),
    .Y(_03910_),
    .B1(net8334));
 sg13g2_nand2_1 _25218_ (.Y(_03911_),
    .A(\soc_I.kianv_I.datapath_unit_I.CSRData[7] ),
    .B(_03910_));
 sg13g2_nand2_1 _25219_ (.Y(_03912_),
    .A(_03909_),
    .B(_03911_));
 sg13g2_inv_2 _25220_ (.Y(_03913_),
    .A(_03912_));
 sg13g2_nor2_1 _25221_ (.A(net8350),
    .B(_03913_),
    .Y(_03914_));
 sg13g2_inv_1 _25222_ (.Y(_03915_),
    .A(_03914_));
 sg13g2_a21oi_1 _25223_ (.A1(net4526),
    .A2(net8487),
    .Y(_03916_),
    .B1(net7706));
 sg13g2_o21ai_1 _25224_ (.B1(net9349),
    .Y(_03917_),
    .A1(net4620),
    .A2(net7702));
 sg13g2_a21oi_1 _25225_ (.A1(_03915_),
    .A2(_03916_),
    .Y(_00847_),
    .B1(_03917_));
 sg13g2_nor3_1 _25226_ (.A(_11207_),
    .B(_03832_),
    .C(net8341),
    .Y(_03918_));
 sg13g2_a21oi_1 _25227_ (.A1(_11208_),
    .A2(net8344),
    .Y(_03919_),
    .B1(net8337));
 sg13g2_a21o_2 _25228_ (.A2(_03919_),
    .A1(\soc_I.kianv_I.datapath_unit_I.CSRData[8] ),
    .B1(_03918_),
    .X(_03920_));
 sg13g2_inv_2 _25229_ (.Y(_03921_),
    .A(_03920_));
 sg13g2_nor2_1 _25230_ (.A(net8350),
    .B(_03921_),
    .Y(_03922_));
 sg13g2_a221oi_1 _25231_ (.B2(_03920_),
    .C1(net7706),
    .B1(net8362),
    .A1(\soc_I.kianv_I.datapath_unit_I.OldPC[8] ),
    .Y(_03923_),
    .A2(net8487));
 sg13g2_o21ai_1 _25232_ (.B1(net9374),
    .Y(_03924_),
    .A1(net4396),
    .A2(net7702));
 sg13g2_nor2_1 _25233_ (.A(_03923_),
    .B(_03924_),
    .Y(_00848_));
 sg13g2_nor2_1 _25234_ (.A(_11246_),
    .B(net8341),
    .Y(_03925_));
 sg13g2_nor2_1 _25235_ (.A(net8337),
    .B(_03925_),
    .Y(_03926_));
 sg13g2_a22oi_1 _25236_ (.Y(_03927_),
    .B1(_03926_),
    .B2(\soc_I.kianv_I.datapath_unit_I.CSRData[9] ),
    .A2(_03925_),
    .A1(net8347));
 sg13g2_nor2_1 _25237_ (.A(net8349),
    .B(_03927_),
    .Y(_03928_));
 sg13g2_a221oi_1 _25238_ (.B2(net7747),
    .C1(_03928_),
    .B1(net8362),
    .A1(\soc_I.kianv_I.datapath_unit_I.OldPC[9] ),
    .Y(_03929_),
    .A2(net8487));
 sg13g2_o21ai_1 _25239_ (.B1(net9349),
    .Y(_03930_),
    .A1(net4580),
    .A2(net7702));
 sg13g2_nor2_1 _25240_ (.A(_03929_),
    .B(_03930_),
    .Y(_00849_));
 sg13g2_nor2_2 _25241_ (.A(_11221_),
    .B(net8342),
    .Y(_03931_));
 sg13g2_nor2_1 _25242_ (.A(net8334),
    .B(_03931_),
    .Y(_03932_));
 sg13g2_a22oi_1 _25243_ (.Y(_03933_),
    .B1(_03932_),
    .B2(\soc_I.kianv_I.datapath_unit_I.CSRData[10] ),
    .A2(_03931_),
    .A1(net8346));
 sg13g2_nand2b_1 _25244_ (.Y(_03934_),
    .B(net8361),
    .A_N(_03933_));
 sg13g2_inv_1 _25245_ (.Y(_03935_),
    .A(_03934_));
 sg13g2_a21oi_1 _25246_ (.A1(\soc_I.kianv_I.datapath_unit_I.OldPC[10] ),
    .A2(net8487),
    .Y(_03936_),
    .B1(net7706));
 sg13g2_o21ai_1 _25247_ (.B1(net9348),
    .Y(_03937_),
    .A1(net4257),
    .A2(net7702));
 sg13g2_a21oi_1 _25248_ (.A1(_03934_),
    .A2(_03936_),
    .Y(_00850_),
    .B1(_03937_));
 sg13g2_and2_1 _25249_ (.A(_11234_),
    .B(net8343),
    .X(_03938_));
 sg13g2_nor2_1 _25250_ (.A(net8334),
    .B(_03938_),
    .Y(_03939_));
 sg13g2_a22oi_1 _25251_ (.Y(_03940_),
    .B1(_03939_),
    .B2(\soc_I.kianv_I.datapath_unit_I.CSRData[11] ),
    .A2(_03938_),
    .A1(net8346));
 sg13g2_nor2_2 _25252_ (.A(net8349),
    .B(_03940_),
    .Y(_03941_));
 sg13g2_a221oi_1 _25253_ (.B2(net7747),
    .C1(_03941_),
    .B1(net8361),
    .A1(net4330),
    .Y(_03942_),
    .A2(net8487));
 sg13g2_o21ai_1 _25254_ (.B1(net9348),
    .Y(_03943_),
    .A1(net4757),
    .A2(net7702));
 sg13g2_nor2_1 _25255_ (.A(_03942_),
    .B(_03943_),
    .Y(_00851_));
 sg13g2_nor2_2 _25256_ (.A(_11292_),
    .B(net8342),
    .Y(_03944_));
 sg13g2_nor2_1 _25257_ (.A(net8334),
    .B(_03944_),
    .Y(_03945_));
 sg13g2_a22oi_1 _25258_ (.Y(_03946_),
    .B1(_03945_),
    .B2(\soc_I.kianv_I.datapath_unit_I.CSRData[12] ),
    .A2(_03944_),
    .A1(net8346));
 sg13g2_nor2_2 _25259_ (.A(net8349),
    .B(_03946_),
    .Y(_03947_));
 sg13g2_a221oi_1 _25260_ (.B2(net7747),
    .C1(_03947_),
    .B1(net8362),
    .A1(\soc_I.kianv_I.datapath_unit_I.OldPC[12] ),
    .Y(_03948_),
    .A2(net8487));
 sg13g2_o21ai_1 _25261_ (.B1(net9363),
    .Y(_03949_),
    .A1(net4744),
    .A2(net7702));
 sg13g2_nor2_1 _25262_ (.A(_03948_),
    .B(_03949_),
    .Y(_00852_));
 sg13g2_nor2_1 _25263_ (.A(net8291),
    .B(net8339),
    .Y(_03950_));
 sg13g2_nor2_1 _25264_ (.A(net8334),
    .B(_03950_),
    .Y(_03951_));
 sg13g2_a22oi_1 _25265_ (.Y(_03952_),
    .B1(_03951_),
    .B2(\soc_I.kianv_I.datapath_unit_I.CSRData[13] ),
    .A2(_03950_),
    .A1(net8346));
 sg13g2_nor2_1 _25266_ (.A(net8351),
    .B(_03952_),
    .Y(_03953_));
 sg13g2_a221oi_1 _25267_ (.B2(net7747),
    .C1(_03953_),
    .B1(net8363),
    .A1(\soc_I.kianv_I.datapath_unit_I.OldPC[13] ),
    .Y(_03954_),
    .A2(net8486));
 sg13g2_o21ai_1 _25268_ (.B1(net9364),
    .Y(_03955_),
    .A1(net4605),
    .A2(net7701));
 sg13g2_nor2_1 _25269_ (.A(_03954_),
    .B(_03955_),
    .Y(_00853_));
 sg13g2_nor2_2 _25270_ (.A(net8295),
    .B(net8340),
    .Y(_03956_));
 sg13g2_nor2_1 _25271_ (.A(net8336),
    .B(_03956_),
    .Y(_03957_));
 sg13g2_a22oi_1 _25272_ (.Y(_03958_),
    .B1(_03957_),
    .B2(\soc_I.kianv_I.datapath_unit_I.CSRData[14] ),
    .A2(_03956_),
    .A1(net8345));
 sg13g2_nor2_1 _25273_ (.A(net8351),
    .B(_03958_),
    .Y(_03959_));
 sg13g2_a221oi_1 _25274_ (.B2(net7747),
    .C1(_03959_),
    .B1(net8363),
    .A1(\soc_I.kianv_I.datapath_unit_I.OldPC[14] ),
    .Y(_03960_),
    .A2(net8486));
 sg13g2_o21ai_1 _25275_ (.B1(net9362),
    .Y(_03961_),
    .A1(net4623),
    .A2(net7701));
 sg13g2_nor2_1 _25276_ (.A(_03960_),
    .B(_03961_),
    .Y(_00854_));
 sg13g2_and2_1 _25277_ (.A(_11280_),
    .B(net8343),
    .X(_03962_));
 sg13g2_nor2_1 _25278_ (.A(net8335),
    .B(_03962_),
    .Y(_03963_));
 sg13g2_a22oi_1 _25279_ (.Y(_03964_),
    .B1(_03963_),
    .B2(\soc_I.kianv_I.datapath_unit_I.CSRData[15] ),
    .A2(_03962_),
    .A1(net8345));
 sg13g2_nand2b_1 _25280_ (.Y(_03965_),
    .B(net8363),
    .A_N(_03964_));
 sg13g2_inv_1 _25281_ (.Y(_03966_),
    .A(_03965_));
 sg13g2_a21oi_1 _25282_ (.A1(net4226),
    .A2(net8486),
    .Y(_03967_),
    .B1(net7706));
 sg13g2_o21ai_1 _25283_ (.B1(net9356),
    .Y(_03968_),
    .A1(net4349),
    .A2(net7701));
 sg13g2_a21oi_1 _25284_ (.A1(_03965_),
    .A2(_03967_),
    .Y(_00855_),
    .B1(_03968_));
 sg13g2_nor2_2 _25285_ (.A(net8283),
    .B(net8340),
    .Y(_03969_));
 sg13g2_nor2_1 _25286_ (.A(net8336),
    .B(_03969_),
    .Y(_03970_));
 sg13g2_a22oi_1 _25287_ (.Y(_03971_),
    .B1(_03970_),
    .B2(\soc_I.kianv_I.datapath_unit_I.CSRData[16] ),
    .A2(_03969_),
    .A1(net8345));
 sg13g2_nand2b_1 _25288_ (.Y(_03972_),
    .B(net8364),
    .A_N(_03971_));
 sg13g2_inv_1 _25289_ (.Y(_03973_),
    .A(_03972_));
 sg13g2_a21oi_1 _25290_ (.A1(\soc_I.kianv_I.datapath_unit_I.OldPC[16] ),
    .A2(net8486),
    .Y(_03974_),
    .B1(net7706));
 sg13g2_o21ai_1 _25291_ (.B1(net9365),
    .Y(_03975_),
    .A1(net4459),
    .A2(net7701));
 sg13g2_a21oi_1 _25292_ (.A1(_03972_),
    .A2(_03974_),
    .Y(_00856_),
    .B1(_03975_));
 sg13g2_nand3_1 _25293_ (.B(net8345),
    .C(net8343),
    .A(net8278),
    .Y(_03976_));
 sg13g2_a21oi_1 _25294_ (.A1(net8278),
    .A2(net8343),
    .Y(_03977_),
    .B1(net8335));
 sg13g2_nand2_1 _25295_ (.Y(_03978_),
    .A(\soc_I.kianv_I.datapath_unit_I.CSRData[17] ),
    .B(_03977_));
 sg13g2_nand2_2 _25296_ (.Y(_03979_),
    .A(_03976_),
    .B(_03978_));
 sg13g2_inv_2 _25297_ (.Y(_03980_),
    .A(_03979_));
 sg13g2_nand2_1 _25298_ (.Y(_03981_),
    .A(net8364),
    .B(_03979_));
 sg13g2_inv_1 _25299_ (.Y(_03982_),
    .A(_03981_));
 sg13g2_a21oi_1 _25300_ (.A1(\soc_I.kianv_I.datapath_unit_I.OldPC[17] ),
    .A2(net8486),
    .Y(_03983_),
    .B1(net7706));
 sg13g2_o21ai_1 _25301_ (.B1(net9365),
    .Y(_03984_),
    .A1(net4357),
    .A2(net7701));
 sg13g2_a21oi_1 _25302_ (.A1(_03981_),
    .A2(_03983_),
    .Y(_00857_),
    .B1(_03984_));
 sg13g2_nor2_1 _25303_ (.A(net8282),
    .B(net8339),
    .Y(_03985_));
 sg13g2_nor2_1 _25304_ (.A(net8335),
    .B(_03985_),
    .Y(_03986_));
 sg13g2_a22oi_1 _25305_ (.Y(_03987_),
    .B1(_03986_),
    .B2(\soc_I.kianv_I.datapath_unit_I.CSRData[18] ),
    .A2(_03985_),
    .A1(net8345));
 sg13g2_nor2_1 _25306_ (.A(net8351),
    .B(_03987_),
    .Y(_03988_));
 sg13g2_a221oi_1 _25307_ (.B2(net7747),
    .C1(_03988_),
    .B1(net8364),
    .A1(\soc_I.kianv_I.datapath_unit_I.OldPC[18] ),
    .Y(_03989_),
    .A2(net8486));
 sg13g2_o21ai_1 _25308_ (.B1(net9368),
    .Y(_03990_),
    .A1(net4868),
    .A2(net7701));
 sg13g2_nor2_1 _25309_ (.A(_03989_),
    .B(_03990_),
    .Y(_00858_));
 sg13g2_nand3_1 _25310_ (.B(net8348),
    .C(net8344),
    .A(_11401_),
    .Y(_03991_));
 sg13g2_a21oi_1 _25311_ (.A1(_11401_),
    .A2(net8344),
    .Y(_03992_),
    .B1(net8336));
 sg13g2_nand2_1 _25312_ (.Y(_03993_),
    .A(\soc_I.kianv_I.datapath_unit_I.CSRData[19] ),
    .B(_03992_));
 sg13g2_nand2_2 _25313_ (.Y(_03994_),
    .A(_03991_),
    .B(_03993_));
 sg13g2_inv_2 _25314_ (.Y(_03995_),
    .A(_03994_));
 sg13g2_nand2_1 _25315_ (.Y(_03996_),
    .A(net8363),
    .B(_03994_));
 sg13g2_inv_1 _25316_ (.Y(_03997_),
    .A(_03996_));
 sg13g2_a21oi_1 _25317_ (.A1(\soc_I.kianv_I.datapath_unit_I.OldPC[19] ),
    .A2(net8486),
    .Y(_03998_),
    .B1(net7706));
 sg13g2_o21ai_1 _25318_ (.B1(net9368),
    .Y(_03999_),
    .A1(net4788),
    .A2(net7701));
 sg13g2_a21oi_1 _25319_ (.A1(_03996_),
    .A2(_03998_),
    .Y(_00859_),
    .B1(_03999_));
 sg13g2_nor2_2 _25320_ (.A(net8286),
    .B(net8342),
    .Y(_04000_));
 sg13g2_nor2_1 _25321_ (.A(net8335),
    .B(_04000_),
    .Y(_04001_));
 sg13g2_a22oi_1 _25322_ (.Y(_04002_),
    .B1(_04001_),
    .B2(\soc_I.kianv_I.datapath_unit_I.CSRData[20] ),
    .A2(_04000_),
    .A1(net8347));
 sg13g2_nor2_1 _25323_ (.A(net8359),
    .B(_04002_),
    .Y(_04003_));
 sg13g2_a221oi_1 _25324_ (.B2(net7748),
    .C1(_04003_),
    .B1(net8369),
    .A1(\soc_I.kianv_I.datapath_unit_I.OldPC[20] ),
    .Y(_04004_),
    .A2(net8490));
 sg13g2_o21ai_1 _25325_ (.B1(net9389),
    .Y(_04005_),
    .A1(net4678),
    .A2(net7703));
 sg13g2_nor2_1 _25326_ (.A(_04004_),
    .B(_04005_),
    .Y(_00860_));
 sg13g2_and2_1 _25327_ (.A(net8285),
    .B(net8344),
    .X(_04006_));
 sg13g2_nor2_1 _25328_ (.A(net8337),
    .B(_04006_),
    .Y(_04007_));
 sg13g2_a22oi_1 _25329_ (.Y(_04008_),
    .B1(_04007_),
    .B2(\soc_I.kianv_I.datapath_unit_I.CSRData[21] ),
    .A2(_04006_),
    .A1(net8347));
 sg13g2_nor2_1 _25330_ (.A(net8358),
    .B(_04008_),
    .Y(_04009_));
 sg13g2_a221oi_1 _25331_ (.B2(net7748),
    .C1(_04009_),
    .B1(net8367),
    .A1(\soc_I.kianv_I.datapath_unit_I.OldPC[21] ),
    .Y(_04010_),
    .A2(net8490));
 sg13g2_o21ai_1 _25332_ (.B1(net9400),
    .Y(_04011_),
    .A1(net4727),
    .A2(net7704));
 sg13g2_nor2_1 _25333_ (.A(_04010_),
    .B(_04011_),
    .Y(_00861_));
 sg13g2_nor2_1 _25334_ (.A(net8289),
    .B(net8342),
    .Y(_04012_));
 sg13g2_nor2_1 _25335_ (.A(net8338),
    .B(_04012_),
    .Y(_04013_));
 sg13g2_a22oi_1 _25336_ (.Y(_04014_),
    .B1(_04013_),
    .B2(\soc_I.kianv_I.datapath_unit_I.CSRData[22] ),
    .A2(_04012_),
    .A1(net8347));
 sg13g2_nor2_1 _25337_ (.A(net8358),
    .B(_04014_),
    .Y(_04015_));
 sg13g2_a221oi_1 _25338_ (.B2(_03852_),
    .C1(_04015_),
    .B1(net8367),
    .A1(\soc_I.kianv_I.datapath_unit_I.OldPC[22] ),
    .Y(_04016_),
    .A2(net8490));
 sg13g2_o21ai_1 _25339_ (.B1(net9399),
    .Y(_04017_),
    .A1(net4741),
    .A2(net7703));
 sg13g2_nor2_1 _25340_ (.A(_04016_),
    .B(_04017_),
    .Y(_00862_));
 sg13g2_nor2_2 _25341_ (.A(_11336_),
    .B(net8342),
    .Y(_04018_));
 sg13g2_nor2_1 _25342_ (.A(net8335),
    .B(_04018_),
    .Y(_04019_));
 sg13g2_a22oi_1 _25343_ (.Y(_04020_),
    .B1(_04019_),
    .B2(\soc_I.kianv_I.datapath_unit_I.CSRData[23] ),
    .A2(_04018_),
    .A1(net8348));
 sg13g2_nor2_1 _25344_ (.A(net8359),
    .B(_04020_),
    .Y(_04021_));
 sg13g2_a221oi_1 _25345_ (.B2(_03852_),
    .C1(_04021_),
    .B1(net8369),
    .A1(net4588),
    .Y(_04022_),
    .A2(net8490));
 sg13g2_o21ai_1 _25346_ (.B1(net9388),
    .Y(_04023_),
    .A1(net4663),
    .A2(net7703));
 sg13g2_nor2_1 _25347_ (.A(_04022_),
    .B(_04023_),
    .Y(_00863_));
 sg13g2_nor3_1 _25348_ (.A(net8272),
    .B(_03832_),
    .C(net8341),
    .Y(_04024_));
 sg13g2_a21oi_1 _25349_ (.A1(_11463_),
    .A2(net8344),
    .Y(_04025_),
    .B1(net8337));
 sg13g2_a21o_2 _25350_ (.A2(_04025_),
    .A1(\soc_I.kianv_I.datapath_unit_I.CSRData[24] ),
    .B1(_04024_),
    .X(_04026_));
 sg13g2_inv_2 _25351_ (.Y(_04027_),
    .A(_04026_));
 sg13g2_nor2_1 _25352_ (.A(net8357),
    .B(_04027_),
    .Y(_04028_));
 sg13g2_a221oi_1 _25353_ (.B2(_04026_),
    .C1(net7705),
    .B1(net8367),
    .A1(\soc_I.kianv_I.datapath_unit_I.OldPC[24] ),
    .Y(_04029_),
    .A2(net8490));
 sg13g2_o21ai_1 _25354_ (.B1(net9389),
    .Y(_04030_),
    .A1(net4577),
    .A2(net7703));
 sg13g2_nor2_1 _25355_ (.A(_04029_),
    .B(_04030_),
    .Y(_00864_));
 sg13g2_nor2_2 _25356_ (.A(net8270),
    .B(net8341),
    .Y(_04031_));
 sg13g2_nor2_1 _25357_ (.A(net8338),
    .B(_04031_),
    .Y(_04032_));
 sg13g2_a22oi_1 _25358_ (.Y(_04033_),
    .B1(_04032_),
    .B2(\soc_I.kianv_I.datapath_unit_I.CSRData[25] ),
    .A2(_04031_),
    .A1(net8347));
 sg13g2_nor2_1 _25359_ (.A(net8357),
    .B(_04033_),
    .Y(_04034_));
 sg13g2_a221oi_1 _25360_ (.B2(net7748),
    .C1(_04034_),
    .B1(net8367),
    .A1(\soc_I.kianv_I.datapath_unit_I.OldPC[25] ),
    .Y(_04035_),
    .A2(net8490));
 sg13g2_o21ai_1 _25361_ (.B1(net9389),
    .Y(_04036_),
    .A1(net4652),
    .A2(net7703));
 sg13g2_nor2_1 _25362_ (.A(_04035_),
    .B(_04036_),
    .Y(_00865_));
 sg13g2_nor2_1 _25363_ (.A(net8275),
    .B(net8342),
    .Y(_04037_));
 sg13g2_nor2_1 _25364_ (.A(net8338),
    .B(_04037_),
    .Y(_04038_));
 sg13g2_a22oi_1 _25365_ (.Y(_04039_),
    .B1(_04038_),
    .B2(\soc_I.kianv_I.datapath_unit_I.CSRData[26] ),
    .A2(_04037_),
    .A1(net8347));
 sg13g2_nor2_1 _25366_ (.A(net8357),
    .B(_04039_),
    .Y(_04040_));
 sg13g2_a221oi_1 _25367_ (.B2(net7748),
    .C1(_04040_),
    .B1(net8367),
    .A1(\soc_I.kianv_I.datapath_unit_I.OldPC[26] ),
    .Y(_04041_),
    .A2(net8490));
 sg13g2_o21ai_1 _25368_ (.B1(net9400),
    .Y(_04042_),
    .A1(net4730),
    .A2(net7703));
 sg13g2_nor2_1 _25369_ (.A(_04041_),
    .B(_04042_),
    .Y(_00866_));
 sg13g2_and2_1 _25370_ (.A(net8274),
    .B(net8344),
    .X(_04043_));
 sg13g2_nor2_1 _25371_ (.A(net8338),
    .B(_04043_),
    .Y(_04044_));
 sg13g2_a22oi_1 _25372_ (.Y(_04045_),
    .B1(_04044_),
    .B2(\soc_I.kianv_I.datapath_unit_I.CSRData[27] ),
    .A2(_04043_),
    .A1(net8348));
 sg13g2_nand2b_1 _25373_ (.Y(_04046_),
    .B(net8369),
    .A_N(_04045_));
 sg13g2_inv_1 _25374_ (.Y(_04047_),
    .A(_04046_));
 sg13g2_a21oi_1 _25375_ (.A1(\soc_I.kianv_I.datapath_unit_I.OldPC[27] ),
    .A2(net8490),
    .Y(_04048_),
    .B1(_03853_));
 sg13g2_o21ai_1 _25376_ (.B1(net9387),
    .Y(_04049_),
    .A1(net4456),
    .A2(net7703));
 sg13g2_a21oi_1 _25377_ (.A1(_04046_),
    .A2(_04048_),
    .Y(_00867_),
    .B1(_04049_));
 sg13g2_nor2_1 _25378_ (.A(net8269),
    .B(net8340),
    .Y(_04050_));
 sg13g2_nor2_1 _25379_ (.A(net8337),
    .B(_04050_),
    .Y(_04051_));
 sg13g2_a22oi_1 _25380_ (.Y(_04052_),
    .B1(_04051_),
    .B2(\soc_I.kianv_I.datapath_unit_I.CSRData[28] ),
    .A2(_04050_),
    .A1(net8348));
 sg13g2_nor2_1 _25381_ (.A(net8352),
    .B(_04052_),
    .Y(_04053_));
 sg13g2_a221oi_1 _25382_ (.B2(net7748),
    .C1(_04053_),
    .B1(net8365),
    .A1(\soc_I.kianv_I.datapath_unit_I.OldPC[28] ),
    .Y(_04054_),
    .A2(net8492));
 sg13g2_o21ai_1 _25383_ (.B1(net9384),
    .Y(_04055_),
    .A1(net4572),
    .A2(_03854_));
 sg13g2_nor2_1 _25384_ (.A(_04054_),
    .B(_04055_),
    .Y(_00868_));
 sg13g2_nor2_1 _25385_ (.A(net8308),
    .B(net8339),
    .Y(_04056_));
 sg13g2_nor2_1 _25386_ (.A(net8335),
    .B(_04056_),
    .Y(_04057_));
 sg13g2_a22oi_1 _25387_ (.Y(_04058_),
    .B1(_04057_),
    .B2(\soc_I.kianv_I.datapath_unit_I.CSRData[29] ),
    .A2(_04056_),
    .A1(net8345));
 sg13g2_nor2_2 _25388_ (.A(net8352),
    .B(_04058_),
    .Y(_04059_));
 sg13g2_a221oi_1 _25389_ (.B2(net7748),
    .C1(_04059_),
    .B1(net8369),
    .A1(\soc_I.kianv_I.datapath_unit_I.OldPC[29] ),
    .Y(_04060_),
    .A2(net8492));
 sg13g2_o21ai_1 _25390_ (.B1(net9383),
    .Y(_04061_),
    .A1(net4461),
    .A2(net7703));
 sg13g2_nor2_1 _25391_ (.A(_04060_),
    .B(_04061_),
    .Y(_00869_));
 sg13g2_nor2_1 _25392_ (.A(_11052_),
    .B(net8339),
    .Y(_04062_));
 sg13g2_nor2_1 _25393_ (.A(net8335),
    .B(_04062_),
    .Y(_04063_));
 sg13g2_a22oi_1 _25394_ (.Y(_04064_),
    .B1(_04063_),
    .B2(\soc_I.kianv_I.datapath_unit_I.CSRData[30] ),
    .A2(_04062_),
    .A1(net8345));
 sg13g2_nor2_1 _25395_ (.A(net8353),
    .B(_04064_),
    .Y(_04065_));
 sg13g2_a221oi_1 _25396_ (.B2(net7747),
    .C1(_04065_),
    .B1(net8366),
    .A1(\soc_I.kianv_I.datapath_unit_I.OldPC[30] ),
    .Y(_04066_),
    .A2(net8487));
 sg13g2_o21ai_1 _25397_ (.B1(net9384),
    .Y(_04067_),
    .A1(net4505),
    .A2(net7702));
 sg13g2_nor2_1 _25398_ (.A(_04066_),
    .B(_04067_),
    .Y(_00870_));
 sg13g2_nor2_1 _25399_ (.A(_10992_),
    .B(net8339),
    .Y(_04068_));
 sg13g2_nor2_1 _25400_ (.A(net8335),
    .B(_04068_),
    .Y(_04069_));
 sg13g2_a22oi_1 _25401_ (.Y(_04070_),
    .B1(_04069_),
    .B2(\soc_I.kianv_I.datapath_unit_I.CSRData[31] ),
    .A2(_04068_),
    .A1(net8345));
 sg13g2_nor2_1 _25402_ (.A(net8352),
    .B(_04070_),
    .Y(_04071_));
 sg13g2_a221oi_1 _25403_ (.B2(net7748),
    .C1(_04071_),
    .B1(net8365),
    .A1(\soc_I.kianv_I.datapath_unit_I.OldPC[31] ),
    .Y(_04072_),
    .A2(net8486));
 sg13g2_o21ai_1 _25404_ (.B1(net9363),
    .Y(_04073_),
    .A1(net4650),
    .A2(net7701));
 sg13g2_nor2_1 _25405_ (.A(_04072_),
    .B(_04073_),
    .Y(_00871_));
 sg13g2_and2_1 _25406_ (.A(net7809),
    .B(net7991),
    .X(_04074_));
 sg13g2_nor2_1 _25407_ (.A(net8359),
    .B(net7744),
    .Y(_04075_));
 sg13g2_nand2b_2 _25408_ (.Y(_04076_),
    .B(net8361),
    .A_N(net7743));
 sg13g2_nand2b_1 _25409_ (.Y(_04077_),
    .B(_03819_),
    .A_N(_00240_));
 sg13g2_nand3_1 _25410_ (.B(_03821_),
    .C(_04077_),
    .A(_03813_),
    .Y(_04078_));
 sg13g2_nor3_1 _25411_ (.A(_03842_),
    .B(net7698),
    .C(_04078_),
    .Y(_04079_));
 sg13g2_o21ai_1 _25412_ (.B1(net9373),
    .Y(_04080_),
    .A1(net4743),
    .A2(_04076_));
 sg13g2_nor2_1 _25413_ (.A(_04079_),
    .B(_04080_),
    .Y(_00872_));
 sg13g2_nand2b_1 _25414_ (.Y(_04081_),
    .B(_03819_),
    .A_N(_00239_));
 sg13g2_a21oi_2 _25415_ (.B1(net8368),
    .Y(_04082_),
    .A2(_04081_),
    .A1(net9198));
 sg13g2_nor3_1 _25416_ (.A(_03863_),
    .B(net7698),
    .C(_04082_),
    .Y(_04083_));
 sg13g2_o21ai_1 _25417_ (.B1(net9372),
    .Y(_04084_),
    .A1(net4522),
    .A2(_04076_));
 sg13g2_nor2_1 _25418_ (.A(_04083_),
    .B(_04084_),
    .Y(_00873_));
 sg13g2_nand3_1 _25419_ (.B(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[7] ),
    .C(\soc_I.kianv_I.control_unit_I.main_fsm_I.mip[7] ),
    .A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[3] ),
    .Y(_04085_));
 sg13g2_o21ai_1 _25420_ (.B1(_03815_),
    .Y(_04086_),
    .A1(_03821_),
    .A2(_04085_));
 sg13g2_a221oi_1 _25421_ (.B2(net4762),
    .C1(_04086_),
    .B1(net7698),
    .A1(_03872_),
    .Y(_04087_),
    .A2(net7745));
 sg13g2_nor2_1 _25422_ (.A(net9038),
    .B(_04087_),
    .Y(_00874_));
 sg13g2_nor3_1 _25423_ (.A(_03819_),
    .B(_03881_),
    .C(net7698),
    .Y(_04088_));
 sg13g2_o21ai_1 _25424_ (.B1(net9372),
    .Y(_04089_),
    .A1(net4655),
    .A2(_04076_));
 sg13g2_nor2_1 _25425_ (.A(_04088_),
    .B(_04089_),
    .Y(_00875_));
 sg13g2_a22oi_1 _25426_ (.Y(_04090_),
    .B1(net7698),
    .B2(net2635),
    .A2(net7745),
    .A1(_03890_));
 sg13g2_nor2_1 _25427_ (.A(net9046),
    .B(_04090_),
    .Y(_00876_));
 sg13g2_a22oi_1 _25428_ (.Y(_04091_),
    .B1(net7698),
    .B2(net2630),
    .A2(net7745),
    .A1(_03897_));
 sg13g2_nor2_1 _25429_ (.A(net9038),
    .B(_04091_),
    .Y(_00877_));
 sg13g2_a22oi_1 _25430_ (.Y(_04092_),
    .B1(net7698),
    .B2(net2805),
    .A2(net7745),
    .A1(_03905_));
 sg13g2_nor2_1 _25431_ (.A(net9046),
    .B(_04092_),
    .Y(_00878_));
 sg13g2_a22oi_1 _25432_ (.Y(_04093_),
    .B1(net7697),
    .B2(net2725),
    .A2(net7743),
    .A1(_03914_));
 sg13g2_nor2_1 _25433_ (.A(net9026),
    .B(_04093_),
    .Y(_00879_));
 sg13g2_a22oi_1 _25434_ (.Y(_04094_),
    .B1(net7697),
    .B2(net2802),
    .A2(net7743),
    .A1(_03922_));
 sg13g2_nor2_1 _25435_ (.A(net9035),
    .B(_04094_),
    .Y(_00880_));
 sg13g2_a22oi_1 _25436_ (.Y(_04095_),
    .B1(net7697),
    .B2(net2715),
    .A2(net7743),
    .A1(_03928_));
 sg13g2_nor2_1 _25437_ (.A(net9023),
    .B(_04095_),
    .Y(_00881_));
 sg13g2_a22oi_1 _25438_ (.Y(_04096_),
    .B1(net7697),
    .B2(net3215),
    .A2(net7743),
    .A1(_03935_));
 sg13g2_nor2_1 _25439_ (.A(net9022),
    .B(_04096_),
    .Y(_00882_));
 sg13g2_a22oi_1 _25440_ (.Y(_04097_),
    .B1(net7697),
    .B2(net2656),
    .A2(net7743),
    .A1(_03941_));
 sg13g2_nor2_1 _25441_ (.A(net9025),
    .B(_04097_),
    .Y(_00883_));
 sg13g2_a22oi_1 _25442_ (.Y(_04098_),
    .B1(net7697),
    .B2(net2696),
    .A2(net7743),
    .A1(_03947_));
 sg13g2_nor2_1 _25443_ (.A(net9025),
    .B(_04098_),
    .Y(_00884_));
 sg13g2_a22oi_1 _25444_ (.Y(_04099_),
    .B1(net7696),
    .B2(net2901),
    .A2(net7742),
    .A1(_03953_));
 sg13g2_nor2_1 _25445_ (.A(net9031),
    .B(_04099_),
    .Y(_00885_));
 sg13g2_a22oi_1 _25446_ (.Y(_04100_),
    .B1(net7696),
    .B2(net2740),
    .A2(net7742),
    .A1(_03959_));
 sg13g2_nor2_1 _25447_ (.A(net9031),
    .B(_04100_),
    .Y(_00886_));
 sg13g2_a22oi_1 _25448_ (.Y(_04101_),
    .B1(net7696),
    .B2(net2803),
    .A2(net7742),
    .A1(_03966_));
 sg13g2_nor2_1 _25449_ (.A(net9031),
    .B(_04101_),
    .Y(_00887_));
 sg13g2_a22oi_1 _25450_ (.Y(_04102_),
    .B1(net7696),
    .B2(net2741),
    .A2(net7742),
    .A1(_03973_));
 sg13g2_nor2_1 _25451_ (.A(net9031),
    .B(_04102_),
    .Y(_00888_));
 sg13g2_a22oi_1 _25452_ (.Y(_04103_),
    .B1(net7696),
    .B2(net2777),
    .A2(net7742),
    .A1(_03982_));
 sg13g2_nor2_1 _25453_ (.A(net9030),
    .B(_04103_),
    .Y(_00889_));
 sg13g2_a22oi_1 _25454_ (.Y(_04104_),
    .B1(net7696),
    .B2(net2687),
    .A2(net7742),
    .A1(_03988_));
 sg13g2_nor2_1 _25455_ (.A(net9030),
    .B(_04104_),
    .Y(_00890_));
 sg13g2_a22oi_1 _25456_ (.Y(_04105_),
    .B1(net7696),
    .B2(net2818),
    .A2(net7742),
    .A1(_03997_));
 sg13g2_nor2_1 _25457_ (.A(net9030),
    .B(_04105_),
    .Y(_00891_));
 sg13g2_a22oi_1 _25458_ (.Y(_04106_),
    .B1(net7699),
    .B2(net2638),
    .A2(net7744),
    .A1(_04003_));
 sg13g2_nor2_1 _25459_ (.A(net9044),
    .B(_04106_),
    .Y(_00892_));
 sg13g2_a22oi_1 _25460_ (.Y(_04107_),
    .B1(net7699),
    .B2(net2667),
    .A2(net7745),
    .A1(_04009_));
 sg13g2_nor2_1 _25461_ (.A(net9050),
    .B(_04107_),
    .Y(_00893_));
 sg13g2_a22oi_1 _25462_ (.Y(_04108_),
    .B1(net7699),
    .B2(net2668),
    .A2(net7744),
    .A1(_04015_));
 sg13g2_nor2_1 _25463_ (.A(net9050),
    .B(_04108_),
    .Y(_00894_));
 sg13g2_a22oi_1 _25464_ (.Y(_04109_),
    .B1(net7699),
    .B2(net2660),
    .A2(net7744),
    .A1(_04021_));
 sg13g2_nor2_1 _25465_ (.A(net9044),
    .B(_04109_),
    .Y(_00895_));
 sg13g2_a22oi_1 _25466_ (.Y(_04110_),
    .B1(net7699),
    .B2(net2772),
    .A2(net7744),
    .A1(_04028_));
 sg13g2_nor2_1 _25467_ (.A(net9044),
    .B(_04110_),
    .Y(_00896_));
 sg13g2_a22oi_1 _25468_ (.Y(_04111_),
    .B1(net7699),
    .B2(net2703),
    .A2(net7744),
    .A1(_04034_));
 sg13g2_nor2_1 _25469_ (.A(net9044),
    .B(_04111_),
    .Y(_00897_));
 sg13g2_a22oi_1 _25470_ (.Y(_04112_),
    .B1(net7698),
    .B2(net2650),
    .A2(net7744),
    .A1(_04040_));
 sg13g2_nor2_1 _25471_ (.A(net9050),
    .B(_04112_),
    .Y(_00898_));
 sg13g2_a22oi_1 _25472_ (.Y(_04113_),
    .B1(net7699),
    .B2(net2746),
    .A2(net7744),
    .A1(_04047_));
 sg13g2_nor2_1 _25473_ (.A(net9044),
    .B(_04113_),
    .Y(_00899_));
 sg13g2_a22oi_1 _25474_ (.Y(_04114_),
    .B1(net7700),
    .B2(net2665),
    .A2(net7746),
    .A1(_04053_));
 sg13g2_nor2_1 _25475_ (.A(net9042),
    .B(_04114_),
    .Y(_00900_));
 sg13g2_a22oi_1 _25476_ (.Y(_04115_),
    .B1(net7700),
    .B2(net2643),
    .A2(net7742),
    .A1(_04059_));
 sg13g2_nor2_1 _25477_ (.A(net9041),
    .B(_04115_),
    .Y(_00901_));
 sg13g2_a22oi_1 _25478_ (.Y(_04116_),
    .B1(net7697),
    .B2(net2739),
    .A2(net7746),
    .A1(_04065_));
 sg13g2_nor2_1 _25479_ (.A(net9031),
    .B(_04116_),
    .Y(_00902_));
 sg13g2_nor3_1 _25480_ (.A(_03820_),
    .B(_04071_),
    .C(net7696),
    .Y(_04117_));
 sg13g2_o21ai_1 _25481_ (.B1(net9363),
    .Y(_04118_),
    .A1(net4774),
    .A2(_04076_));
 sg13g2_nor2_1 _25482_ (.A(_04117_),
    .B(_04118_),
    .Y(_00903_));
 sg13g2_nand3_1 _25483_ (.B(_03842_),
    .C(net7993),
    .A(net7802),
    .Y(_04119_));
 sg13g2_a21oi_1 _25484_ (.A1(net7803),
    .A2(net7993),
    .Y(_04120_),
    .B1(net8357));
 sg13g2_a21o_1 _25485_ (.A2(net7992),
    .A1(net7804),
    .B1(net8360),
    .X(_04121_));
 sg13g2_a22oi_1 _25486_ (.Y(_04122_),
    .B1(net7740),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[0] ),
    .A2(net8355),
    .A1(net3999));
 sg13g2_a21oi_1 _25487_ (.A1(_04119_),
    .A2(net4000),
    .Y(_00904_),
    .B1(net9038));
 sg13g2_nand3_1 _25488_ (.B(net7993),
    .C(_03863_),
    .A(net7802),
    .Y(_04123_));
 sg13g2_a22oi_1 _25489_ (.Y(_04124_),
    .B1(net7740),
    .B2(net4878),
    .A2(net8354),
    .A1(net4541));
 sg13g2_a21oi_1 _25490_ (.A1(_04123_),
    .A2(_04124_),
    .Y(_00905_),
    .B1(net9038));
 sg13g2_nand3_1 _25491_ (.B(net7993),
    .C(_03872_),
    .A(net7806),
    .Y(_04125_));
 sg13g2_a22oi_1 _25492_ (.Y(_04126_),
    .B1(net7740),
    .B2(net4667),
    .A2(net8355),
    .A1(net4590));
 sg13g2_a21oi_1 _25493_ (.A1(_04125_),
    .A2(_04126_),
    .Y(_00906_),
    .B1(net9046));
 sg13g2_a21oi_1 _25494_ (.A1(net4452),
    .A2(net8356),
    .Y(_04127_),
    .B1(_03881_));
 sg13g2_o21ai_1 _25495_ (.B1(net9372),
    .Y(_04128_),
    .A1(net4891),
    .A2(net7736));
 sg13g2_a21oi_1 _25496_ (.A1(net7736),
    .A2(_04127_),
    .Y(_00907_),
    .B1(_04128_));
 sg13g2_a21oi_1 _25497_ (.A1(\soc_I.kianv_I.datapath_unit_I.OldPC[4] ),
    .A2(net8354),
    .Y(_04129_),
    .B1(_03890_));
 sg13g2_o21ai_1 _25498_ (.B1(net9393),
    .Y(_04130_),
    .A1(net4853),
    .A2(net7736));
 sg13g2_a21oi_1 _25499_ (.A1(net7736),
    .A2(_04129_),
    .Y(_00908_),
    .B1(_04130_));
 sg13g2_a21oi_1 _25500_ (.A1(\soc_I.kianv_I.datapath_unit_I.OldPC[5] ),
    .A2(net8356),
    .Y(_04131_),
    .B1(_03897_));
 sg13g2_o21ai_1 _25501_ (.B1(net9378),
    .Y(_04132_),
    .A1(net4695),
    .A2(net7736));
 sg13g2_a21oi_1 _25502_ (.A1(net7736),
    .A2(_04131_),
    .Y(_00909_),
    .B1(_04132_));
 sg13g2_a21oi_1 _25503_ (.A1(\soc_I.kianv_I.datapath_unit_I.OldPC[6] ),
    .A2(net8355),
    .Y(_04133_),
    .B1(_03905_));
 sg13g2_o21ai_1 _25504_ (.B1(net9393),
    .Y(_04134_),
    .A1(net4732),
    .A2(net7736));
 sg13g2_a21oi_1 _25505_ (.A1(net7736),
    .A2(_04133_),
    .Y(_00910_),
    .B1(_04134_));
 sg13g2_a21oi_1 _25506_ (.A1(net4526),
    .A2(net8350),
    .Y(_04135_),
    .B1(net7738));
 sg13g2_o21ai_1 _25507_ (.B1(net9349),
    .Y(_04136_),
    .A1(net5064),
    .A2(net7734));
 sg13g2_a21oi_1 _25508_ (.A1(_03915_),
    .A2(_04135_),
    .Y(_00911_),
    .B1(_04136_));
 sg13g2_nand3_1 _25509_ (.B(net7990),
    .C(_03922_),
    .A(net7798),
    .Y(_04137_));
 sg13g2_a22oi_1 _25510_ (.Y(_04138_),
    .B1(net7738),
    .B2(net4670),
    .A2(net8350),
    .A1(\soc_I.kianv_I.datapath_unit_I.OldPC[8] ));
 sg13g2_a21oi_1 _25511_ (.A1(_04137_),
    .A2(net4671),
    .Y(_00912_),
    .B1(net9036));
 sg13g2_a21oi_1 _25512_ (.A1(\soc_I.kianv_I.datapath_unit_I.OldPC[9] ),
    .A2(net8349),
    .Y(_04139_),
    .B1(_03928_));
 sg13g2_o21ai_1 _25513_ (.B1(net9348),
    .Y(_04140_),
    .A1(net4780),
    .A2(net7734));
 sg13g2_a21oi_1 _25514_ (.A1(net7734),
    .A2(_04139_),
    .Y(_00913_),
    .B1(_04140_));
 sg13g2_o21ai_1 _25515_ (.B1(net9348),
    .Y(_04141_),
    .A1(net4055),
    .A2(net7734));
 sg13g2_a21oi_1 _25516_ (.A1(net4797),
    .A2(net8349),
    .Y(_04142_),
    .B1(net7738));
 sg13g2_a21oi_1 _25517_ (.A1(_03934_),
    .A2(_04142_),
    .Y(_00914_),
    .B1(_04141_));
 sg13g2_nand3_1 _25518_ (.B(net7990),
    .C(_03941_),
    .A(net7798),
    .Y(_04143_));
 sg13g2_a22oi_1 _25519_ (.Y(_04144_),
    .B1(net7738),
    .B2(net4598),
    .A2(net8349),
    .A1(net4330));
 sg13g2_a21oi_1 _25520_ (.A1(_04143_),
    .A2(_04144_),
    .Y(_00915_),
    .B1(net9025));
 sg13g2_nand3_1 _25521_ (.B(net7990),
    .C(_03947_),
    .A(net7798),
    .Y(_04145_));
 sg13g2_a22oi_1 _25522_ (.Y(_04146_),
    .B1(net7738),
    .B2(net4295),
    .A2(net8350),
    .A1(\soc_I.kianv_I.datapath_unit_I.OldPC[12] ));
 sg13g2_a21oi_1 _25523_ (.A1(_04145_),
    .A2(net4296),
    .Y(_00916_),
    .B1(net9025));
 sg13g2_a21oi_1 _25524_ (.A1(\soc_I.kianv_I.datapath_unit_I.OldPC[13] ),
    .A2(net8351),
    .Y(_04147_),
    .B1(_03953_));
 sg13g2_o21ai_1 _25525_ (.B1(net9364),
    .Y(_04148_),
    .A1(net4798),
    .A2(net7735));
 sg13g2_a21oi_1 _25526_ (.A1(net7735),
    .A2(_04147_),
    .Y(_00917_),
    .B1(_04148_));
 sg13g2_a21oi_1 _25527_ (.A1(\soc_I.kianv_I.datapath_unit_I.OldPC[14] ),
    .A2(net8351),
    .Y(_04149_),
    .B1(_03959_));
 sg13g2_o21ai_1 _25528_ (.B1(net9361),
    .Y(_04150_),
    .A1(net4881),
    .A2(net7734));
 sg13g2_a21oi_1 _25529_ (.A1(net7734),
    .A2(_04149_),
    .Y(_00918_),
    .B1(_04150_));
 sg13g2_o21ai_1 _25530_ (.B1(net9356),
    .Y(_04151_),
    .A1(net4910),
    .A2(net7734));
 sg13g2_a21oi_1 _25531_ (.A1(net4226),
    .A2(net8351),
    .Y(_04152_),
    .B1(net7739));
 sg13g2_a21oi_1 _25532_ (.A1(_03965_),
    .A2(_04152_),
    .Y(_00919_),
    .B1(_04151_));
 sg13g2_o21ai_1 _25533_ (.B1(net9359),
    .Y(_04153_),
    .A1(net4992),
    .A2(net7734));
 sg13g2_a21oi_1 _25534_ (.A1(\soc_I.kianv_I.datapath_unit_I.OldPC[16] ),
    .A2(net8351),
    .Y(_04154_),
    .B1(net7739));
 sg13g2_a21oi_1 _25535_ (.A1(_03972_),
    .A2(_04154_),
    .Y(_00920_),
    .B1(_04153_));
 sg13g2_o21ai_1 _25536_ (.B1(net9359),
    .Y(_04155_),
    .A1(net4883),
    .A2(net7735));
 sg13g2_a21oi_1 _25537_ (.A1(\soc_I.kianv_I.datapath_unit_I.OldPC[17] ),
    .A2(net8351),
    .Y(_04156_),
    .B1(net7739));
 sg13g2_a21oi_1 _25538_ (.A1(_03981_),
    .A2(_04156_),
    .Y(_00921_),
    .B1(_04155_));
 sg13g2_nand3_1 _25539_ (.B(net7991),
    .C(_03988_),
    .A(net7799),
    .Y(_04157_));
 sg13g2_a22oi_1 _25540_ (.Y(_04158_),
    .B1(net7739),
    .B2(net4932),
    .A2(net8352),
    .A1(\soc_I.kianv_I.datapath_unit_I.OldPC[18] ));
 sg13g2_a21oi_1 _25541_ (.A1(_04157_),
    .A2(net4933),
    .Y(_00922_),
    .B1(net9027));
 sg13g2_o21ai_1 _25542_ (.B1(net9359),
    .Y(_04159_),
    .A1(net4905),
    .A2(net7735));
 sg13g2_a21oi_1 _25543_ (.A1(\soc_I.kianv_I.datapath_unit_I.OldPC[19] ),
    .A2(net8352),
    .Y(_04160_),
    .B1(net7739));
 sg13g2_a21oi_1 _25544_ (.A1(_03996_),
    .A2(_04160_),
    .Y(_00923_),
    .B1(_04159_));
 sg13g2_nand3_1 _25545_ (.B(net7992),
    .C(_04003_),
    .A(net7805),
    .Y(_04161_));
 sg13g2_a22oi_1 _25546_ (.Y(_04162_),
    .B1(net7740),
    .B2(net4643),
    .A2(net8357),
    .A1(\soc_I.kianv_I.datapath_unit_I.OldPC[20] ));
 sg13g2_a21oi_1 _25547_ (.A1(_04161_),
    .A2(net4644),
    .Y(_00924_),
    .B1(net9045));
 sg13g2_nand3_1 _25548_ (.B(net7993),
    .C(_04009_),
    .A(net7804),
    .Y(_04163_));
 sg13g2_a22oi_1 _25549_ (.Y(_04164_),
    .B1(net7740),
    .B2(net5135),
    .A2(net8357),
    .A1(net4785));
 sg13g2_a21oi_1 _25550_ (.A1(_04163_),
    .A2(_04164_),
    .Y(_00925_),
    .B1(net9050));
 sg13g2_nand3_1 _25551_ (.B(net7992),
    .C(_04015_),
    .A(net7803),
    .Y(_04165_));
 sg13g2_a22oi_1 _25552_ (.Y(_04166_),
    .B1(net7740),
    .B2(net4840),
    .A2(net8358),
    .A1(\soc_I.kianv_I.datapath_unit_I.OldPC[22] ));
 sg13g2_a21oi_1 _25553_ (.A1(_04165_),
    .A2(net4841),
    .Y(_00926_),
    .B1(net9050));
 sg13g2_nand3_1 _25554_ (.B(net7992),
    .C(_04021_),
    .A(net7805),
    .Y(_04167_));
 sg13g2_a22oi_1 _25555_ (.Y(_04168_),
    .B1(net7741),
    .B2(net4764),
    .A2(net8359),
    .A1(net4588));
 sg13g2_a21oi_1 _25556_ (.A1(_04167_),
    .A2(_04168_),
    .Y(_00927_),
    .B1(net9044));
 sg13g2_nand3_1 _25557_ (.B(net7992),
    .C(_04028_),
    .A(net7803),
    .Y(_04169_));
 sg13g2_a22oi_1 _25558_ (.Y(_04170_),
    .B1(net7740),
    .B2(net4778),
    .A2(net8358),
    .A1(\soc_I.kianv_I.datapath_unit_I.OldPC[24] ));
 sg13g2_a21oi_1 _25559_ (.A1(_04169_),
    .A2(net4779),
    .Y(_00928_),
    .B1(net9050));
 sg13g2_nand3_1 _25560_ (.B(net7992),
    .C(_04034_),
    .A(net7803),
    .Y(_04171_));
 sg13g2_a22oi_1 _25561_ (.Y(_04172_),
    .B1(net7740),
    .B2(net4861),
    .A2(net8357),
    .A1(\soc_I.kianv_I.datapath_unit_I.OldPC[25] ));
 sg13g2_a21oi_1 _25562_ (.A1(_04171_),
    .A2(net4862),
    .Y(_00929_),
    .B1(net9044));
 sg13g2_a21oi_1 _25563_ (.A1(\soc_I.kianv_I.datapath_unit_I.OldPC[26] ),
    .A2(net8358),
    .Y(_04173_),
    .B1(_04040_));
 sg13g2_o21ai_1 _25564_ (.B1(net9399),
    .Y(_04174_),
    .A1(net4876),
    .A2(net7737));
 sg13g2_a21oi_1 _25565_ (.A1(net7737),
    .A2(_04173_),
    .Y(_00930_),
    .B1(_04174_));
 sg13g2_o21ai_1 _25566_ (.B1(net9387),
    .Y(_04175_),
    .A1(net4801),
    .A2(net7737));
 sg13g2_a21oi_1 _25567_ (.A1(net4783),
    .A2(net8359),
    .Y(_04176_),
    .B1(net7741));
 sg13g2_a21oi_1 _25568_ (.A1(_04046_),
    .A2(_04176_),
    .Y(_00931_),
    .B1(_04175_));
 sg13g2_nand3_1 _25569_ (.B(net7990),
    .C(_04053_),
    .A(net7800),
    .Y(_04177_));
 sg13g2_a22oi_1 _25570_ (.Y(_04178_),
    .B1(net7738),
    .B2(net4397),
    .A2(net8352),
    .A1(\soc_I.kianv_I.datapath_unit_I.OldPC[28] ));
 sg13g2_a21oi_1 _25571_ (.A1(_04177_),
    .A2(net4398),
    .Y(_00932_),
    .B1(net9041));
 sg13g2_nand3_1 _25572_ (.B(net7990),
    .C(_04059_),
    .A(net7800),
    .Y(_04179_));
 sg13g2_a22oi_1 _25573_ (.Y(_04180_),
    .B1(net7741),
    .B2(net4874),
    .A2(net8359),
    .A1(net4994));
 sg13g2_a21oi_1 _25574_ (.A1(_04179_),
    .A2(_04180_),
    .Y(_00933_),
    .B1(net9041));
 sg13g2_nand3_1 _25575_ (.B(net7991),
    .C(_04065_),
    .A(net7800),
    .Y(_04181_));
 sg13g2_a22oi_1 _25576_ (.Y(_04182_),
    .B1(net7738),
    .B2(net4711),
    .A2(net8353),
    .A1(\soc_I.kianv_I.datapath_unit_I.OldPC[30] ));
 sg13g2_a21oi_1 _25577_ (.A1(_04181_),
    .A2(net4712),
    .Y(_00934_),
    .B1(net9040));
 sg13g2_nand3_1 _25578_ (.B(net7990),
    .C(_04071_),
    .A(net7800),
    .Y(_04183_));
 sg13g2_a22oi_1 _25579_ (.Y(_04184_),
    .B1(net7738),
    .B2(net4406),
    .A2(net8352),
    .A1(\soc_I.kianv_I.datapath_unit_I.OldPC[31] ));
 sg13g2_a21oi_1 _25580_ (.A1(_04183_),
    .A2(net4407),
    .Y(_00935_),
    .B1(net9031));
 sg13g2_and2_1 _25581_ (.A(net7783),
    .B(net7991),
    .X(_04185_));
 sg13g2_o21ai_1 _25582_ (.B1(net9374),
    .Y(_04186_),
    .A1(net4925),
    .A2(net7723));
 sg13g2_a21oi_1 _25583_ (.A1(_03841_),
    .A2(net7723),
    .Y(_00936_),
    .B1(_04186_));
 sg13g2_o21ai_1 _25584_ (.B1(net9373),
    .Y(_04187_),
    .A1(net4781),
    .A2(net7730));
 sg13g2_a21oi_1 _25585_ (.A1(_03862_),
    .A2(net7730),
    .Y(_00937_),
    .B1(_04187_));
 sg13g2_o21ai_1 _25586_ (.B1(net9376),
    .Y(_04188_),
    .A1(net5091),
    .A2(net7730));
 sg13g2_a21oi_1 _25587_ (.A1(_03871_),
    .A2(net7733),
    .Y(_00938_),
    .B1(_04188_));
 sg13g2_o21ai_1 _25588_ (.B1(net9374),
    .Y(_04189_),
    .A1(net5339),
    .A2(net7723));
 sg13g2_a21oi_1 _25589_ (.A1(_03880_),
    .A2(net7723),
    .Y(_00939_),
    .B1(_04189_));
 sg13g2_o21ai_1 _25590_ (.B1(net9379),
    .Y(_04190_),
    .A1(net5269),
    .A2(net7730));
 sg13g2_a21oi_1 _25591_ (.A1(_03889_),
    .A2(net7730),
    .Y(_00940_),
    .B1(_04190_));
 sg13g2_o21ai_1 _25592_ (.B1(net9379),
    .Y(_04191_),
    .A1(net5354),
    .A2(net7730));
 sg13g2_a21oi_1 _25593_ (.A1(_03896_),
    .A2(net7730),
    .Y(_00941_),
    .B1(_04191_));
 sg13g2_o21ai_1 _25594_ (.B1(net9378),
    .Y(_04192_),
    .A1(net4995),
    .A2(net7733));
 sg13g2_a21oi_1 _25595_ (.A1(_03904_),
    .A2(net7730),
    .Y(_00942_),
    .B1(_04192_));
 sg13g2_o21ai_1 _25596_ (.B1(net9349),
    .Y(_04193_),
    .A1(net5197),
    .A2(net7723));
 sg13g2_a21oi_1 _25597_ (.A1(_03913_),
    .A2(net7723),
    .Y(_00943_),
    .B1(_04193_));
 sg13g2_o21ai_1 _25598_ (.B1(net9352),
    .Y(_04194_),
    .A1(net4957),
    .A2(net7723));
 sg13g2_a21oi_1 _25599_ (.A1(_03921_),
    .A2(net7723),
    .Y(_00944_),
    .B1(_04194_));
 sg13g2_o21ai_1 _25600_ (.B1(net9352),
    .Y(_04195_),
    .A1(net5027),
    .A2(net7725));
 sg13g2_a21oi_1 _25601_ (.A1(_03927_),
    .A2(net7725),
    .Y(_00945_),
    .B1(_04195_));
 sg13g2_o21ai_1 _25602_ (.B1(net9352),
    .Y(_04196_),
    .A1(net5168),
    .A2(net7725));
 sg13g2_a21oi_1 _25603_ (.A1(_03933_),
    .A2(net7725),
    .Y(_00946_),
    .B1(_04196_));
 sg13g2_o21ai_1 _25604_ (.B1(net9350),
    .Y(_04197_),
    .A1(net4907),
    .A2(net7724));
 sg13g2_a21oi_1 _25605_ (.A1(_03940_),
    .A2(net7724),
    .Y(_00947_),
    .B1(_04197_));
 sg13g2_o21ai_1 _25606_ (.B1(net9362),
    .Y(_04198_),
    .A1(net5026),
    .A2(net7724));
 sg13g2_a21oi_1 _25607_ (.A1(_03946_),
    .A2(net7724),
    .Y(_00948_),
    .B1(_04198_));
 sg13g2_o21ai_1 _25608_ (.B1(net9356),
    .Y(_04199_),
    .A1(net5029),
    .A2(net7726));
 sg13g2_a21oi_1 _25609_ (.A1(_03952_),
    .A2(net7726),
    .Y(_00949_),
    .B1(_04199_));
 sg13g2_o21ai_1 _25610_ (.B1(net9356),
    .Y(_04200_),
    .A1(net5147),
    .A2(net7726));
 sg13g2_a21oi_1 _25611_ (.A1(_03958_),
    .A2(net7726),
    .Y(_00950_),
    .B1(_04200_));
 sg13g2_o21ai_1 _25612_ (.B1(net9362),
    .Y(_04201_),
    .A1(net4900),
    .A2(net7726));
 sg13g2_a21oi_1 _25613_ (.A1(_03964_),
    .A2(net7726),
    .Y(_00951_),
    .B1(_04201_));
 sg13g2_o21ai_1 _25614_ (.B1(net9357),
    .Y(_04202_),
    .A1(net4968),
    .A2(net7727));
 sg13g2_a21oi_1 _25615_ (.A1(_03971_),
    .A2(net7727),
    .Y(_00952_),
    .B1(_04202_));
 sg13g2_o21ai_1 _25616_ (.B1(net9357),
    .Y(_04203_),
    .A1(net5164),
    .A2(net7726));
 sg13g2_a21oi_1 _25617_ (.A1(_03980_),
    .A2(net7726),
    .Y(_00953_),
    .B1(_04203_));
 sg13g2_o21ai_1 _25618_ (.B1(net9358),
    .Y(_04204_),
    .A1(net5141),
    .A2(net7727));
 sg13g2_a21oi_1 _25619_ (.A1(_03987_),
    .A2(net7727),
    .Y(_00954_),
    .B1(_04204_));
 sg13g2_o21ai_1 _25620_ (.B1(net9358),
    .Y(_04205_),
    .A1(net5046),
    .A2(net7727));
 sg13g2_a21oi_1 _25621_ (.A1(_03995_),
    .A2(net7727),
    .Y(_00955_),
    .B1(_04205_));
 sg13g2_o21ai_1 _25622_ (.B1(net9385),
    .Y(_04206_),
    .A1(net5107),
    .A2(net7732));
 sg13g2_a21oi_1 _25623_ (.A1(_04002_),
    .A2(net7732),
    .Y(_00956_),
    .B1(_04206_));
 sg13g2_o21ai_1 _25624_ (.B1(net9401),
    .Y(_04207_),
    .A1(net5209),
    .A2(net7731));
 sg13g2_a21oi_1 _25625_ (.A1(_04008_),
    .A2(net7731),
    .Y(_00957_),
    .B1(_04207_));
 sg13g2_o21ai_1 _25626_ (.B1(net9402),
    .Y(_04208_),
    .A1(net5165),
    .A2(net7731));
 sg13g2_a21oi_1 _25627_ (.A1(_04014_),
    .A2(net7732),
    .Y(_00958_),
    .B1(_04208_));
 sg13g2_o21ai_1 _25628_ (.B1(net9388),
    .Y(_04209_),
    .A1(net5251),
    .A2(net7732));
 sg13g2_a21oi_1 _25629_ (.A1(_04020_),
    .A2(net7732),
    .Y(_00959_),
    .B1(_04209_));
 sg13g2_o21ai_1 _25630_ (.B1(net9389),
    .Y(_04210_),
    .A1(net5517),
    .A2(net7731));
 sg13g2_a21oi_1 _25631_ (.A1(_04027_),
    .A2(net7731),
    .Y(_00960_),
    .B1(_04210_));
 sg13g2_o21ai_1 _25632_ (.B1(net9400),
    .Y(_04211_),
    .A1(net5322),
    .A2(net7731));
 sg13g2_a21oi_1 _25633_ (.A1(_04033_),
    .A2(net7731),
    .Y(_00961_),
    .B1(_04211_));
 sg13g2_o21ai_1 _25634_ (.B1(net9401),
    .Y(_04212_),
    .A1(net5126),
    .A2(net7731));
 sg13g2_a21oi_1 _25635_ (.A1(_04039_),
    .A2(net7732),
    .Y(_00962_),
    .B1(_04212_));
 sg13g2_o21ai_1 _25636_ (.B1(net9385),
    .Y(_04213_),
    .A1(net5190),
    .A2(net7732));
 sg13g2_a21oi_1 _25637_ (.A1(_04045_),
    .A2(net7732),
    .Y(_00963_),
    .B1(_04213_));
 sg13g2_o21ai_1 _25638_ (.B1(net9384),
    .Y(_04214_),
    .A1(net5028),
    .A2(net7728));
 sg13g2_a21oi_1 _25639_ (.A1(_04052_),
    .A2(net7728),
    .Y(_00964_),
    .B1(_04214_));
 sg13g2_o21ai_1 _25640_ (.B1(net9366),
    .Y(_04215_),
    .A1(net5018),
    .A2(net7729));
 sg13g2_a21oi_1 _25641_ (.A1(_04058_),
    .A2(net7729),
    .Y(_00965_),
    .B1(_04215_));
 sg13g2_o21ai_1 _25642_ (.B1(net9366),
    .Y(_04216_),
    .A1(net5133),
    .A2(net7728));
 sg13g2_a21oi_1 _25643_ (.A1(_04064_),
    .A2(net7728),
    .Y(_00966_),
    .B1(_04216_));
 sg13g2_o21ai_1 _25644_ (.B1(net9363),
    .Y(_04217_),
    .A1(net5134),
    .A2(net7728));
 sg13g2_a21oi_1 _25645_ (.A1(_04070_),
    .A2(net7728),
    .Y(_00967_),
    .B1(_04217_));
 sg13g2_and2_1 _25646_ (.A(net7906),
    .B(net7990),
    .X(_04218_));
 sg13g2_o21ai_1 _25647_ (.B1(net9374),
    .Y(_04219_),
    .A1(net4436),
    .A2(net7777));
 sg13g2_a21oi_1 _25648_ (.A1(_03841_),
    .A2(net7777),
    .Y(_00968_),
    .B1(_04219_));
 sg13g2_o21ai_1 _25649_ (.B1(net9372),
    .Y(_04220_),
    .A1(net4291),
    .A2(net7772));
 sg13g2_a21oi_1 _25650_ (.A1(_03862_),
    .A2(net7772),
    .Y(_00969_),
    .B1(_04220_));
 sg13g2_o21ai_1 _25651_ (.B1(net9379),
    .Y(_04221_),
    .A1(net4770),
    .A2(net7780));
 sg13g2_a21oi_1 _25652_ (.A1(_03871_),
    .A2(net7780),
    .Y(_00970_),
    .B1(_04221_));
 sg13g2_o21ai_1 _25653_ (.B1(net9373),
    .Y(_04222_),
    .A1(net4567),
    .A2(net7772));
 sg13g2_a21oi_1 _25654_ (.A1(_03880_),
    .A2(net7772),
    .Y(_00971_),
    .B1(_04222_));
 sg13g2_o21ai_1 _25655_ (.B1(net9395),
    .Y(_04223_),
    .A1(net4617),
    .A2(net7780));
 sg13g2_a21oi_1 _25656_ (.A1(_03889_),
    .A2(net7780),
    .Y(_00972_),
    .B1(_04223_));
 sg13g2_o21ai_1 _25657_ (.B1(net9379),
    .Y(_04224_),
    .A1(net4836),
    .A2(net7780));
 sg13g2_a21oi_1 _25658_ (.A1(_03896_),
    .A2(net7780),
    .Y(_00973_),
    .B1(_04224_));
 sg13g2_o21ai_1 _25659_ (.B1(net9395),
    .Y(_04225_),
    .A1(net4554),
    .A2(net7780));
 sg13g2_a21oi_1 _25660_ (.A1(_03904_),
    .A2(net7780),
    .Y(_00974_),
    .B1(_04225_));
 sg13g2_o21ai_1 _25661_ (.B1(net9350),
    .Y(_04226_),
    .A1(net4529),
    .A2(net7772));
 sg13g2_a21oi_1 _25662_ (.A1(_03913_),
    .A2(net7772),
    .Y(_00975_),
    .B1(_04226_));
 sg13g2_o21ai_1 _25663_ (.B1(net9370),
    .Y(_04227_),
    .A1(net4464),
    .A2(net7772));
 sg13g2_a21oi_1 _25664_ (.A1(_03921_),
    .A2(net7772),
    .Y(_00976_),
    .B1(_04227_));
 sg13g2_o21ai_1 _25665_ (.B1(net9352),
    .Y(_04228_),
    .A1(net4612),
    .A2(net7773));
 sg13g2_a21oi_1 _25666_ (.A1(_03927_),
    .A2(net7773),
    .Y(_00977_),
    .B1(_04228_));
 sg13g2_o21ai_1 _25667_ (.B1(net9346),
    .Y(_04229_),
    .A1(net4680),
    .A2(net7773));
 sg13g2_a21oi_1 _25668_ (.A1(_03933_),
    .A2(net7773),
    .Y(_00978_),
    .B1(_04229_));
 sg13g2_o21ai_1 _25669_ (.B1(net9350),
    .Y(_04230_),
    .A1(net4539),
    .A2(net7773));
 sg13g2_a21oi_1 _25670_ (.A1(_03940_),
    .A2(net7773),
    .Y(_00979_),
    .B1(_04230_));
 sg13g2_o21ai_1 _25671_ (.B1(net9363),
    .Y(_04231_),
    .A1(net4665),
    .A2(net7773));
 sg13g2_a21oi_1 _25672_ (.A1(_03946_),
    .A2(net7773),
    .Y(_00980_),
    .B1(_04231_));
 sg13g2_o21ai_1 _25673_ (.B1(net9355),
    .Y(_04232_),
    .A1(net4517),
    .A2(net7774));
 sg13g2_a21oi_1 _25674_ (.A1(_03952_),
    .A2(net7774),
    .Y(_00981_),
    .B1(_04232_));
 sg13g2_o21ai_1 _25675_ (.B1(net9364),
    .Y(_04233_),
    .A1(net4585),
    .A2(net7774));
 sg13g2_a21oi_1 _25676_ (.A1(_03958_),
    .A2(net7774),
    .Y(_00982_),
    .B1(_04233_));
 sg13g2_o21ai_1 _25677_ (.B1(net9354),
    .Y(_04234_),
    .A1(net4453),
    .A2(net7774));
 sg13g2_a21oi_1 _25678_ (.A1(_03964_),
    .A2(net7774),
    .Y(_00983_),
    .B1(_04234_));
 sg13g2_o21ai_1 _25679_ (.B1(net9365),
    .Y(_04235_),
    .A1(net4611),
    .A2(net7774));
 sg13g2_a21oi_1 _25680_ (.A1(_03971_),
    .A2(net7774),
    .Y(_00984_),
    .B1(_04235_));
 sg13g2_o21ai_1 _25681_ (.B1(net9365),
    .Y(_04236_),
    .A1(net4445),
    .A2(net7775));
 sg13g2_a21oi_1 _25682_ (.A1(_03980_),
    .A2(net7775),
    .Y(_00985_),
    .B1(_04236_));
 sg13g2_o21ai_1 _25683_ (.B1(net9365),
    .Y(_04237_),
    .A1(net4516),
    .A2(net7775));
 sg13g2_a21oi_1 _25684_ (.A1(_03987_),
    .A2(net7775),
    .Y(_00986_),
    .B1(_04237_));
 sg13g2_o21ai_1 _25685_ (.B1(net9360),
    .Y(_04238_),
    .A1(net4370),
    .A2(net7775));
 sg13g2_a21oi_1 _25686_ (.A1(_03995_),
    .A2(net7775),
    .Y(_00987_),
    .B1(_04238_));
 sg13g2_o21ai_1 _25687_ (.B1(net9387),
    .Y(_04239_),
    .A1(net4538),
    .A2(net7779));
 sg13g2_a21oi_1 _25688_ (.A1(_04002_),
    .A2(net7779),
    .Y(_00988_),
    .B1(_04239_));
 sg13g2_o21ai_1 _25689_ (.B1(net9399),
    .Y(_04240_),
    .A1(net4373),
    .A2(net7778));
 sg13g2_a21oi_1 _25690_ (.A1(_04008_),
    .A2(net7778),
    .Y(_00989_),
    .B1(_04240_));
 sg13g2_o21ai_1 _25691_ (.B1(net9400),
    .Y(_04241_),
    .A1(net4385),
    .A2(net7778));
 sg13g2_a21oi_1 _25692_ (.A1(_04014_),
    .A2(net7778),
    .Y(_00990_),
    .B1(_04241_));
 sg13g2_o21ai_1 _25693_ (.B1(net9388),
    .Y(_04242_),
    .A1(net4525),
    .A2(net7779));
 sg13g2_a21oi_1 _25694_ (.A1(_04020_),
    .A2(net7779),
    .Y(_00991_),
    .B1(_04242_));
 sg13g2_o21ai_1 _25695_ (.B1(net9390),
    .Y(_04243_),
    .A1(net4471),
    .A2(net7778));
 sg13g2_a21oi_1 _25696_ (.A1(_04027_),
    .A2(net7778),
    .Y(_00992_),
    .B1(_04243_));
 sg13g2_o21ai_1 _25697_ (.B1(net9389),
    .Y(_04244_),
    .A1(net4600),
    .A2(net7778));
 sg13g2_a21oi_1 _25698_ (.A1(_04033_),
    .A2(net7778),
    .Y(_00993_),
    .B1(_04244_));
 sg13g2_o21ai_1 _25699_ (.B1(net9399),
    .Y(_04245_),
    .A1(net4515),
    .A2(net7779));
 sg13g2_a21oi_1 _25700_ (.A1(_04039_),
    .A2(net7779),
    .Y(_00994_),
    .B1(_04245_));
 sg13g2_o21ai_1 _25701_ (.B1(net9388),
    .Y(_04246_),
    .A1(net4528),
    .A2(net7779));
 sg13g2_a21oi_1 _25702_ (.A1(_04045_),
    .A2(net7779),
    .Y(_00995_),
    .B1(_04246_));
 sg13g2_o21ai_1 _25703_ (.B1(net9384),
    .Y(_04247_),
    .A1(net4576),
    .A2(net7776));
 sg13g2_a21oi_1 _25704_ (.A1(_04052_),
    .A2(net7776),
    .Y(_00996_),
    .B1(_04247_));
 sg13g2_o21ai_1 _25705_ (.B1(net9366),
    .Y(_04248_),
    .A1(net4309),
    .A2(net7776));
 sg13g2_a21oi_1 _25706_ (.A1(_04058_),
    .A2(net7776),
    .Y(_00997_),
    .B1(_04248_));
 sg13g2_o21ai_1 _25707_ (.B1(net9366),
    .Y(_04249_),
    .A1(net4579),
    .A2(net7777));
 sg13g2_a21oi_1 _25708_ (.A1(_04064_),
    .A2(net7777),
    .Y(_00998_),
    .B1(_04249_));
 sg13g2_o21ai_1 _25709_ (.B1(net9363),
    .Y(_04250_),
    .A1(net4371),
    .A2(net7776));
 sg13g2_a21oi_1 _25710_ (.A1(_04070_),
    .A2(net7776),
    .Y(_00999_),
    .B1(_04250_));
 sg13g2_nor3_1 _25711_ (.A(net8977),
    .B(_10841_),
    .C(_10861_),
    .Y(_04251_));
 sg13g2_nand2_2 _25712_ (.Y(_04252_),
    .A(net8978),
    .B(_13830_));
 sg13g2_nor2_1 _25713_ (.A(net8357),
    .B(net8805),
    .Y(_04253_));
 sg13g2_nand2_2 _25714_ (.Y(_04254_),
    .A(net8365),
    .B(_04252_));
 sg13g2_nor2_1 _25715_ (.A(net9023),
    .B(net8120),
    .Y(_01000_));
 sg13g2_and2_2 _25716_ (.A(net5145),
    .B(net9356),
    .X(_01001_));
 sg13g2_nor2b_1 _25717_ (.A(\soc_I.clint_I.mtime[39] ),
    .B_N(\soc_I.clint_I.mtimecmp[39] ),
    .Y(_04255_));
 sg13g2_nor2_1 _25718_ (.A(_10414_),
    .B(\soc_I.clint_I.mtimecmp[39] ),
    .Y(_04256_));
 sg13g2_nor2_1 _25719_ (.A(_10415_),
    .B(\soc_I.clint_I.mtimecmp[38] ),
    .Y(_04257_));
 sg13g2_a22oi_1 _25720_ (.Y(_04258_),
    .B1(\soc_I.clint_I.mtimecmp[36] ),
    .B2(_10417_),
    .A2(\soc_I.clint_I.mtimecmp[37] ),
    .A1(_10416_));
 sg13g2_a22oi_1 _25721_ (.Y(_04259_),
    .B1(_10447_),
    .B2(\soc_I.clint_I.mtime[35] ),
    .A2(_10446_),
    .A1(\soc_I.clint_I.mtime[36] ));
 sg13g2_a22oi_1 _25722_ (.Y(_04260_),
    .B1(\soc_I.clint_I.mtimecmp[34] ),
    .B2(_10419_),
    .A2(\soc_I.clint_I.mtimecmp[35] ),
    .A1(_10418_));
 sg13g2_nor2_1 _25723_ (.A(\soc_I.clint_I.mtime[33] ),
    .B(_10449_),
    .Y(_04261_));
 sg13g2_nand2b_1 _25724_ (.Y(_04262_),
    .B(\soc_I.clint_I.mtime[32] ),
    .A_N(\soc_I.clint_I.mtimecmp[32] ));
 sg13g2_a22oi_1 _25725_ (.Y(_04263_),
    .B1(_10449_),
    .B2(\soc_I.clint_I.mtime[33] ),
    .A2(_10448_),
    .A1(\soc_I.clint_I.mtime[34] ));
 sg13g2_o21ai_1 _25726_ (.B1(_04263_),
    .Y(_04264_),
    .A1(_04261_),
    .A2(_04262_));
 sg13g2_nand2_1 _25727_ (.Y(_04265_),
    .A(_04260_),
    .B(_04264_));
 sg13g2_and2_1 _25728_ (.A(_04259_),
    .B(_04265_),
    .X(_04266_));
 sg13g2_nand2b_1 _25729_ (.Y(_04267_),
    .B(_04258_),
    .A_N(_04266_));
 sg13g2_nand2b_1 _25730_ (.Y(_04268_),
    .B(\soc_I.clint_I.mtime[37] ),
    .A_N(\soc_I.clint_I.mtimecmp[37] ));
 sg13g2_a22oi_1 _25731_ (.Y(_04269_),
    .B1(_04267_),
    .B2(_04268_),
    .A2(\soc_I.clint_I.mtimecmp[38] ),
    .A1(_10415_));
 sg13g2_nor3_1 _25732_ (.A(_04256_),
    .B(_04257_),
    .C(_04269_),
    .Y(_04270_));
 sg13g2_nor2_1 _25733_ (.A(_04255_),
    .B(_04270_),
    .Y(_04271_));
 sg13g2_nor2b_1 _25734_ (.A(\soc_I.clint_I.mtimecmp[28] ),
    .B_N(\soc_I.clint_I.mtime[28] ),
    .Y(_04272_));
 sg13g2_nor2b_1 _25735_ (.A(\soc_I.clint_I.mtime[27] ),
    .B_N(\soc_I.clint_I.mtimecmp[27] ),
    .Y(_04273_));
 sg13g2_nand2b_1 _25736_ (.Y(_04274_),
    .B(\soc_I.clint_I.mtime[25] ),
    .A_N(\soc_I.clint_I.mtimecmp[25] ));
 sg13g2_o21ai_1 _25737_ (.B1(_04274_),
    .Y(_04275_),
    .A1(_10426_),
    .A2(\soc_I.clint_I.mtimecmp[24] ));
 sg13g2_nor2b_1 _25738_ (.A(\soc_I.clint_I.mtimecmp[27] ),
    .B_N(\soc_I.clint_I.mtime[27] ),
    .Y(_04276_));
 sg13g2_nor2b_1 _25739_ (.A(\soc_I.clint_I.mtime[26] ),
    .B_N(\soc_I.clint_I.mtimecmp[26] ),
    .Y(_04277_));
 sg13g2_nor2_1 _25740_ (.A(_04276_),
    .B(_04277_),
    .Y(_04278_));
 sg13g2_nand2_1 _25741_ (.Y(_04279_),
    .A(_10425_),
    .B(\soc_I.clint_I.mtimecmp[25] ));
 sg13g2_nand3_1 _25742_ (.B(_04278_),
    .C(_04279_),
    .A(_04275_),
    .Y(_04280_));
 sg13g2_nand2b_1 _25743_ (.Y(_04281_),
    .B(\soc_I.clint_I.mtime[26] ),
    .A_N(\soc_I.clint_I.mtimecmp[26] ));
 sg13g2_a21oi_1 _25744_ (.A1(_04280_),
    .A2(_04281_),
    .Y(_04282_),
    .B1(_04273_));
 sg13g2_nor3_1 _25745_ (.A(_04272_),
    .B(_04276_),
    .C(_04282_),
    .Y(_04283_));
 sg13g2_a22oi_1 _25746_ (.Y(_04284_),
    .B1(\soc_I.clint_I.mtimecmp[30] ),
    .B2(_10422_),
    .A2(\soc_I.clint_I.mtimecmp[31] ),
    .A1(_10421_));
 sg13g2_nand2b_1 _25747_ (.Y(_04285_),
    .B(\soc_I.clint_I.mtimecmp[28] ),
    .A_N(\soc_I.clint_I.mtime[28] ));
 sg13g2_nand2_1 _25748_ (.Y(_04286_),
    .A(_10423_),
    .B(\soc_I.clint_I.mtimecmp[29] ));
 sg13g2_nand2_1 _25749_ (.Y(_04287_),
    .A(_04285_),
    .B(_04286_));
 sg13g2_nand3_1 _25750_ (.B(_04285_),
    .C(_04286_),
    .A(_04284_),
    .Y(_04288_));
 sg13g2_a22oi_1 _25751_ (.Y(_04289_),
    .B1(_10560_),
    .B2(\soc_I.clint_I.mtime[29] ),
    .A2(_10559_),
    .A1(\soc_I.clint_I.mtime[30] ));
 sg13g2_o21ai_1 _25752_ (.B1(_04289_),
    .Y(_04290_),
    .A1(_04283_),
    .A2(_04287_));
 sg13g2_nand2_1 _25753_ (.Y(_04291_),
    .A(_10432_),
    .B(\soc_I.clint_I.mtimecmp[15] ));
 sg13g2_nand2b_1 _25754_ (.Y(_04292_),
    .B(\soc_I.clint_I.mtime[15] ),
    .A_N(\soc_I.clint_I.mtimecmp[15] ));
 sg13g2_o21ai_1 _25755_ (.B1(_04292_),
    .Y(_04293_),
    .A1(_10433_),
    .A2(\soc_I.clint_I.mtimecmp[14] ));
 sg13g2_a22oi_1 _25756_ (.Y(_04294_),
    .B1(_10566_),
    .B2(\soc_I.clint_I.mtime[12] ),
    .A2(_10565_),
    .A1(\soc_I.clint_I.mtime[13] ));
 sg13g2_a22oi_1 _25757_ (.Y(_04295_),
    .B1(\soc_I.clint_I.mtimecmp[13] ),
    .B2(_10434_),
    .A2(\soc_I.clint_I.mtimecmp[14] ),
    .A1(_10433_));
 sg13g2_nor2b_1 _25758_ (.A(_04294_),
    .B_N(_04295_),
    .Y(_04296_));
 sg13g2_o21ai_1 _25759_ (.B1(_04291_),
    .Y(_04297_),
    .A1(_04293_),
    .A2(_04296_));
 sg13g2_nand2b_1 _25760_ (.Y(_04298_),
    .B(\soc_I.clint_I.mtimecmp[2] ),
    .A_N(\soc_I.clint_I.mtime[2] ));
 sg13g2_a22oi_1 _25761_ (.Y(_04299_),
    .B1(\soc_I.clint_I.mtimecmp[0] ),
    .B2(_10445_),
    .A2(\soc_I.clint_I.mtimecmp[1] ),
    .A1(_10444_));
 sg13g2_nand2b_1 _25762_ (.Y(_04300_),
    .B(\soc_I.clint_I.mtime[2] ),
    .A_N(\soc_I.clint_I.mtimecmp[2] ));
 sg13g2_o21ai_1 _25763_ (.B1(_04300_),
    .Y(_04301_),
    .A1(_10444_),
    .A2(\soc_I.clint_I.mtimecmp[1] ));
 sg13g2_o21ai_1 _25764_ (.B1(_04298_),
    .Y(_04302_),
    .A1(_04299_),
    .A2(_04301_));
 sg13g2_o21ai_1 _25765_ (.B1(_04302_),
    .Y(_04303_),
    .A1(_10443_),
    .A2(\soc_I.clint_I.mtimecmp[3] ));
 sg13g2_a22oi_1 _25766_ (.Y(_04304_),
    .B1(\soc_I.clint_I.mtimecmp[3] ),
    .B2(_10443_),
    .A2(\soc_I.clint_I.mtimecmp[4] ),
    .A1(_10442_));
 sg13g2_nand2b_1 _25767_ (.Y(_04305_),
    .B(\soc_I.clint_I.mtime[5] ),
    .A_N(\soc_I.clint_I.mtimecmp[5] ));
 sg13g2_o21ai_1 _25768_ (.B1(_04305_),
    .Y(_04306_),
    .A1(_10442_),
    .A2(\soc_I.clint_I.mtimecmp[4] ));
 sg13g2_a21oi_1 _25769_ (.A1(_04303_),
    .A2(_04304_),
    .Y(_04307_),
    .B1(_04306_));
 sg13g2_a221oi_1 _25770_ (.B2(_10441_),
    .C1(_04307_),
    .B1(\soc_I.clint_I.mtimecmp[5] ),
    .A1(_10440_),
    .Y(_04308_),
    .A2(\soc_I.clint_I.mtimecmp[6] ));
 sg13g2_nand2b_1 _25771_ (.Y(_04309_),
    .B(\soc_I.clint_I.mtime[6] ),
    .A_N(\soc_I.clint_I.mtimecmp[6] ));
 sg13g2_o21ai_1 _25772_ (.B1(_04309_),
    .Y(_04310_),
    .A1(_10439_),
    .A2(\soc_I.clint_I.mtimecmp[7] ));
 sg13g2_a22oi_1 _25773_ (.Y(_04311_),
    .B1(\soc_I.clint_I.mtimecmp[7] ),
    .B2(_10439_),
    .A2(\soc_I.clint_I.mtimecmp[8] ),
    .A1(_10438_));
 sg13g2_o21ai_1 _25774_ (.B1(_04311_),
    .Y(_04312_),
    .A1(_04308_),
    .A2(_04310_));
 sg13g2_a22oi_1 _25775_ (.Y(_04313_),
    .B1(_10570_),
    .B2(\soc_I.clint_I.mtime[8] ),
    .A2(_10569_),
    .A1(\soc_I.clint_I.mtime[9] ));
 sg13g2_nand2_1 _25776_ (.Y(_04314_),
    .A(_10435_),
    .B(\soc_I.clint_I.mtimecmp[11] ));
 sg13g2_o21ai_1 _25777_ (.B1(_04314_),
    .Y(_04315_),
    .A1(\soc_I.clint_I.mtime[10] ),
    .A2(_10568_));
 sg13g2_a221oi_1 _25778_ (.B2(_04313_),
    .C1(_04315_),
    .B1(_04312_),
    .A1(_10437_),
    .Y(_04316_),
    .A2(\soc_I.clint_I.mtimecmp[9] ));
 sg13g2_a221oi_1 _25779_ (.B2(\soc_I.clint_I.mtime[10] ),
    .C1(_04316_),
    .B1(_10568_),
    .A1(\soc_I.clint_I.mtime[11] ),
    .Y(_04317_),
    .A2(_10567_));
 sg13g2_o21ai_1 _25780_ (.B1(_04291_),
    .Y(_04318_),
    .A1(\soc_I.clint_I.mtime[12] ),
    .A2(_10566_));
 sg13g2_nor3_2 _25781_ (.A(_10436_),
    .B(\soc_I.clint_I.mtimecmp[10] ),
    .C(_04314_),
    .Y(_04319_));
 sg13g2_nand2_1 _25782_ (.Y(_04320_),
    .A(_04294_),
    .B(_04295_));
 sg13g2_or4_1 _25783_ (.A(_04293_),
    .B(_04318_),
    .C(_04319_),
    .D(_04320_),
    .X(_04321_));
 sg13g2_o21ai_1 _25784_ (.B1(_04297_),
    .Y(_04322_),
    .A1(_04317_),
    .A2(_04321_));
 sg13g2_a22oi_1 _25785_ (.Y(_04323_),
    .B1(_10562_),
    .B2(\soc_I.clint_I.mtime[22] ),
    .A2(_10561_),
    .A1(\soc_I.clint_I.mtime[23] ));
 sg13g2_nor2_1 _25786_ (.A(\soc_I.clint_I.mtime[23] ),
    .B(_10561_),
    .Y(_04324_));
 sg13g2_a21oi_1 _25787_ (.A1(_10430_),
    .A2(\soc_I.clint_I.mtimecmp[18] ),
    .Y(_04325_),
    .B1(_04324_));
 sg13g2_a22oi_1 _25788_ (.Y(_04326_),
    .B1(_10564_),
    .B2(\soc_I.clint_I.mtime[20] ),
    .A2(_10563_),
    .A1(\soc_I.clint_I.mtime[21] ));
 sg13g2_nand2b_1 _25789_ (.Y(_04327_),
    .B(\soc_I.clint_I.mtimecmp[22] ),
    .A_N(\soc_I.clint_I.mtime[22] ));
 sg13g2_o21ai_1 _25790_ (.B1(_04327_),
    .Y(_04328_),
    .A1(\soc_I.clint_I.mtime[21] ),
    .A2(_10563_));
 sg13g2_a22oi_1 _25791_ (.Y(_04329_),
    .B1(\soc_I.clint_I.mtimecmp[19] ),
    .B2(_10429_),
    .A2(\soc_I.clint_I.mtimecmp[20] ),
    .A1(_10428_));
 sg13g2_nand2b_1 _25792_ (.Y(_04330_),
    .B(\soc_I.clint_I.mtime[19] ),
    .A_N(\soc_I.clint_I.mtimecmp[19] ));
 sg13g2_o21ai_1 _25793_ (.B1(_04330_),
    .Y(_04331_),
    .A1(_10430_),
    .A2(\soc_I.clint_I.mtimecmp[18] ));
 sg13g2_nand2_1 _25794_ (.Y(_04332_),
    .A(_04323_),
    .B(_04326_));
 sg13g2_nor3_1 _25795_ (.A(_04328_),
    .B(_04331_),
    .C(_04332_),
    .Y(_04333_));
 sg13g2_nand3_1 _25796_ (.B(_04329_),
    .C(_04333_),
    .A(_04325_),
    .Y(_04334_));
 sg13g2_nand2b_1 _25797_ (.Y(_04335_),
    .B(\soc_I.clint_I.mtime[16] ),
    .A_N(\soc_I.clint_I.mtimecmp[16] ));
 sg13g2_o21ai_1 _25798_ (.B1(_04335_),
    .Y(_04336_),
    .A1(_10431_),
    .A2(\soc_I.clint_I.mtimecmp[17] ));
 sg13g2_nor2b_1 _25799_ (.A(\soc_I.clint_I.mtime[17] ),
    .B_N(\soc_I.clint_I.mtimecmp[17] ),
    .Y(_04337_));
 sg13g2_nor2b_1 _25800_ (.A(\soc_I.clint_I.mtime[16] ),
    .B_N(\soc_I.clint_I.mtimecmp[16] ),
    .Y(_04338_));
 sg13g2_nor4_1 _25801_ (.A(_04334_),
    .B(_04336_),
    .C(_04337_),
    .D(_04338_),
    .Y(_04339_));
 sg13g2_nand2_1 _25802_ (.Y(_04340_),
    .A(_04329_),
    .B(_04331_));
 sg13g2_a21o_1 _25803_ (.A2(_04340_),
    .A1(_04326_),
    .B1(_04328_),
    .X(_04341_));
 sg13g2_a21oi_1 _25804_ (.A1(_04323_),
    .A2(_04341_),
    .Y(_04342_),
    .B1(_04324_));
 sg13g2_nor2_1 _25805_ (.A(_04334_),
    .B(_04337_),
    .Y(_04343_));
 sg13g2_a221oi_1 _25806_ (.B2(_04336_),
    .C1(_04342_),
    .B1(_04343_),
    .A1(_04322_),
    .Y(_04344_),
    .A2(_04339_));
 sg13g2_nor4_1 _25807_ (.A(_04272_),
    .B(_04273_),
    .C(_04276_),
    .D(_04277_),
    .Y(_04345_));
 sg13g2_nand3b_1 _25808_ (.B(_04289_),
    .C(_04345_),
    .Y(_04346_),
    .A_N(_04275_));
 sg13g2_nand2_1 _25809_ (.Y(_04347_),
    .A(_10426_),
    .B(\soc_I.clint_I.mtimecmp[24] ));
 sg13g2_nand3_1 _25810_ (.B(_04281_),
    .C(_04347_),
    .A(_04279_),
    .Y(_04348_));
 sg13g2_nor4_1 _25811_ (.A(_04288_),
    .B(_04344_),
    .C(_04346_),
    .D(_04348_),
    .Y(_04349_));
 sg13g2_a221oi_1 _25812_ (.B2(_04290_),
    .C1(_04349_),
    .B1(_04284_),
    .A1(\soc_I.clint_I.mtime[31] ),
    .Y(_04350_),
    .A2(_10558_));
 sg13g2_nand4_1 _25813_ (.B(_04259_),
    .C(_04260_),
    .A(_04258_),
    .Y(_04351_),
    .D(_04263_));
 sg13g2_a22oi_1 _25814_ (.Y(_04352_),
    .B1(\soc_I.clint_I.mtimecmp[32] ),
    .B2(_10420_),
    .A2(\soc_I.clint_I.mtimecmp[38] ),
    .A1(_10415_));
 sg13g2_nand3_1 _25815_ (.B(_04268_),
    .C(_04352_),
    .A(_04262_),
    .Y(_04353_));
 sg13g2_or4_1 _25816_ (.A(_04255_),
    .B(_04256_),
    .C(_04257_),
    .D(_04261_),
    .X(_04354_));
 sg13g2_nor4_1 _25817_ (.A(_04350_),
    .B(_04351_),
    .C(_04353_),
    .D(_04354_),
    .Y(_04355_));
 sg13g2_nor2_1 _25818_ (.A(\soc_I.clint_I.mtime[40] ),
    .B(_10586_),
    .Y(_04356_));
 sg13g2_nor2_1 _25819_ (.A(\soc_I.clint_I.mtime[41] ),
    .B(_10585_),
    .Y(_04357_));
 sg13g2_nor2_1 _25820_ (.A(_10410_),
    .B(\soc_I.clint_I.mtimecmp[47] ),
    .Y(_04358_));
 sg13g2_nor2_1 _25821_ (.A(_10413_),
    .B(\soc_I.clint_I.mtimecmp[44] ),
    .Y(_04359_));
 sg13g2_or4_1 _25822_ (.A(_04356_),
    .B(_04357_),
    .C(_04358_),
    .D(_04359_),
    .X(_04360_));
 sg13g2_a22oi_1 _25823_ (.Y(_04361_),
    .B1(_10582_),
    .B2(\soc_I.clint_I.mtime[45] ),
    .A2(_10581_),
    .A1(\soc_I.clint_I.mtime[46] ));
 sg13g2_a22oi_1 _25824_ (.Y(_04362_),
    .B1(_10586_),
    .B2(\soc_I.clint_I.mtime[40] ),
    .A2(_10585_),
    .A1(\soc_I.clint_I.mtime[41] ));
 sg13g2_a22oi_1 _25825_ (.Y(_04363_),
    .B1(_10584_),
    .B2(\soc_I.clint_I.mtime[42] ),
    .A2(_10583_),
    .A1(\soc_I.clint_I.mtime[43] ));
 sg13g2_nand2b_1 _25826_ (.Y(_04364_),
    .B(\soc_I.clint_I.mtimecmp[42] ),
    .A_N(\soc_I.clint_I.mtime[42] ));
 sg13g2_nand2b_1 _25827_ (.Y(_04365_),
    .B(\soc_I.clint_I.mtimecmp[43] ),
    .A_N(\soc_I.clint_I.mtime[43] ));
 sg13g2_nand3_1 _25828_ (.B(_04364_),
    .C(_04365_),
    .A(_04363_),
    .Y(_04366_));
 sg13g2_a22oi_1 _25829_ (.Y(_04367_),
    .B1(\soc_I.clint_I.mtimecmp[44] ),
    .B2(_10413_),
    .A2(\soc_I.clint_I.mtimecmp[45] ),
    .A1(_10412_));
 sg13g2_a22oi_1 _25830_ (.Y(_04368_),
    .B1(\soc_I.clint_I.mtimecmp[46] ),
    .B2(_10411_),
    .A2(\soc_I.clint_I.mtimecmp[47] ),
    .A1(_10410_));
 sg13g2_nand4_1 _25831_ (.B(_04362_),
    .C(_04367_),
    .A(_04361_),
    .Y(_04369_),
    .D(_04368_));
 sg13g2_nor3_2 _25832_ (.A(_04360_),
    .B(_04366_),
    .C(_04369_),
    .Y(_04370_));
 sg13g2_o21ai_1 _25833_ (.B1(_04370_),
    .Y(_04371_),
    .A1(_04271_),
    .A2(_04355_));
 sg13g2_nor3_1 _25834_ (.A(_04357_),
    .B(_04362_),
    .C(_04366_),
    .Y(_04372_));
 sg13g2_nor2b_1 _25835_ (.A(_04363_),
    .B_N(_04365_),
    .Y(_04373_));
 sg13g2_nor3_1 _25836_ (.A(_04359_),
    .B(_04372_),
    .C(_04373_),
    .Y(_04374_));
 sg13g2_nand2b_1 _25837_ (.Y(_04375_),
    .B(_04367_),
    .A_N(_04374_));
 sg13g2_nand2_1 _25838_ (.Y(_04376_),
    .A(_04361_),
    .B(_04375_));
 sg13g2_a21oi_2 _25839_ (.B1(_04358_),
    .Y(_04377_),
    .A2(_04376_),
    .A1(_04368_));
 sg13g2_nand2_2 _25840_ (.Y(_04378_),
    .A(_04371_),
    .B(_04377_));
 sg13g2_a22oi_1 _25841_ (.Y(_04379_),
    .B1(_10574_),
    .B2(\soc_I.clint_I.mtime[58] ),
    .A2(_10573_),
    .A1(\soc_I.clint_I.mtime[59] ));
 sg13g2_nand2b_1 _25842_ (.Y(_04380_),
    .B(\soc_I.clint_I.mtimecmp[58] ),
    .A_N(\soc_I.clint_I.mtime[58] ));
 sg13g2_nand2_1 _25843_ (.Y(_04381_),
    .A(_10403_),
    .B(\soc_I.clint_I.mtimecmp[59] ));
 sg13g2_nand3_1 _25844_ (.B(_04380_),
    .C(_04381_),
    .A(_04379_),
    .Y(_04382_));
 sg13g2_a22oi_1 _25845_ (.Y(_04383_),
    .B1(\soc_I.clint_I.mtimecmp[62] ),
    .B2(_10400_),
    .A2(\soc_I.clint_I.mtimecmp[63] ),
    .A1(_10399_));
 sg13g2_a22oi_1 _25846_ (.Y(_04384_),
    .B1(\soc_I.clint_I.mtimecmp[60] ),
    .B2(_10402_),
    .A2(\soc_I.clint_I.mtimecmp[61] ),
    .A1(_10401_));
 sg13g2_nand2_1 _25847_ (.Y(_04385_),
    .A(_04383_),
    .B(_04384_));
 sg13g2_nand2b_1 _25848_ (.Y(_04386_),
    .B(\soc_I.clint_I.mtime[61] ),
    .A_N(\soc_I.clint_I.mtimecmp[61] ));
 sg13g2_o21ai_1 _25849_ (.B1(_04386_),
    .Y(_04387_),
    .A1(_10400_),
    .A2(\soc_I.clint_I.mtimecmp[62] ));
 sg13g2_a21oi_1 _25850_ (.A1(_10405_),
    .A2(\soc_I.clint_I.mtimecmp[56] ),
    .Y(_04388_),
    .B1(_04387_));
 sg13g2_a22oi_1 _25851_ (.Y(_04389_),
    .B1(_10578_),
    .B2(\soc_I.clint_I.mtime[53] ),
    .A2(_10577_),
    .A1(\soc_I.clint_I.mtime[54] ));
 sg13g2_nor2b_1 _25852_ (.A(\soc_I.clint_I.mtime[55] ),
    .B_N(\soc_I.clint_I.mtimecmp[55] ),
    .Y(_04390_));
 sg13g2_nor2_1 _25853_ (.A(\soc_I.clint_I.mtime[54] ),
    .B(_10577_),
    .Y(_04391_));
 sg13g2_nand2b_1 _25854_ (.Y(_04392_),
    .B(\soc_I.clint_I.mtime[51] ),
    .A_N(\soc_I.clint_I.mtimecmp[51] ));
 sg13g2_nand2b_1 _25855_ (.Y(_04393_),
    .B(\soc_I.clint_I.mtimecmp[50] ),
    .A_N(\soc_I.clint_I.mtime[50] ));
 sg13g2_a22oi_1 _25856_ (.Y(_04394_),
    .B1(\soc_I.clint_I.mtimecmp[52] ),
    .B2(_10408_),
    .A2(\soc_I.clint_I.mtimecmp[53] ),
    .A1(_10407_));
 sg13g2_nor2_1 _25857_ (.A(_10402_),
    .B(\soc_I.clint_I.mtimecmp[60] ),
    .Y(_04395_));
 sg13g2_a21o_1 _25858_ (.A2(_10572_),
    .A1(\soc_I.clint_I.mtime[63] ),
    .B1(_04395_),
    .X(_04396_));
 sg13g2_a22oi_1 _25859_ (.Y(_04397_),
    .B1(_10576_),
    .B2(\soc_I.clint_I.mtime[56] ),
    .A2(_10575_),
    .A1(\soc_I.clint_I.mtime[57] ));
 sg13g2_a22oi_1 _25860_ (.Y(_04398_),
    .B1(_10580_),
    .B2(\soc_I.clint_I.mtime[48] ),
    .A2(_10579_),
    .A1(\soc_I.clint_I.mtime[49] ));
 sg13g2_nor2b_1 _25861_ (.A(\soc_I.clint_I.mtimecmp[55] ),
    .B_N(\soc_I.clint_I.mtime[55] ),
    .Y(_04399_));
 sg13g2_nand2_1 _25862_ (.Y(_04400_),
    .A(_10404_),
    .B(\soc_I.clint_I.mtimecmp[57] ));
 sg13g2_nand2b_1 _25863_ (.Y(_04401_),
    .B(\soc_I.clint_I.mtimecmp[51] ),
    .A_N(\soc_I.clint_I.mtime[51] ));
 sg13g2_nand2_1 _25864_ (.Y(_04402_),
    .A(_10409_),
    .B(\soc_I.clint_I.mtimecmp[48] ));
 sg13g2_nand2b_1 _25865_ (.Y(_04403_),
    .B(\soc_I.clint_I.mtimecmp[49] ),
    .A_N(\soc_I.clint_I.mtime[49] ));
 sg13g2_nand2b_1 _25866_ (.Y(_04404_),
    .B(\soc_I.clint_I.mtime[50] ),
    .A_N(\soc_I.clint_I.mtimecmp[50] ));
 sg13g2_nor2_1 _25867_ (.A(_10408_),
    .B(\soc_I.clint_I.mtimecmp[52] ),
    .Y(_04405_));
 sg13g2_nand4_1 _25868_ (.B(_04402_),
    .C(_04403_),
    .A(_04401_),
    .Y(_04406_),
    .D(_04404_));
 sg13g2_nand3_1 _25869_ (.B(_04397_),
    .C(_04400_),
    .A(_04388_),
    .Y(_04407_));
 sg13g2_nor4_1 _25870_ (.A(_04382_),
    .B(_04385_),
    .C(_04390_),
    .D(_04391_),
    .Y(_04408_));
 sg13g2_or3_1 _25871_ (.A(_04399_),
    .B(_04405_),
    .C(_04406_),
    .X(_04409_));
 sg13g2_nand4_1 _25872_ (.B(_04392_),
    .C(_04393_),
    .A(_04389_),
    .Y(_04410_),
    .D(_04398_));
 sg13g2_nor4_1 _25873_ (.A(_04396_),
    .B(_04407_),
    .C(_04409_),
    .D(_04410_),
    .Y(_04411_));
 sg13g2_nand4_1 _25874_ (.B(_04394_),
    .C(_04408_),
    .A(_04378_),
    .Y(_04412_),
    .D(_04411_));
 sg13g2_nand3_1 _25875_ (.B(_04393_),
    .C(_04403_),
    .A(_04392_),
    .Y(_04413_));
 sg13g2_o21ai_1 _25876_ (.B1(_04404_),
    .Y(_04414_),
    .A1(_04398_),
    .A2(_04413_));
 sg13g2_nand2_1 _25877_ (.Y(_04415_),
    .A(_04401_),
    .B(_04414_));
 sg13g2_nand2_1 _25878_ (.Y(_04416_),
    .A(_04392_),
    .B(_04415_));
 sg13g2_o21ai_1 _25879_ (.B1(_04394_),
    .Y(_04417_),
    .A1(_04405_),
    .A2(_04416_));
 sg13g2_a221oi_1 _25880_ (.B2(_04417_),
    .C1(_04390_),
    .B1(_04389_),
    .A1(_10406_),
    .Y(_04418_),
    .A2(\soc_I.clint_I.mtimecmp[54] ));
 sg13g2_o21ai_1 _25881_ (.B1(_04388_),
    .Y(_04419_),
    .A1(_04399_),
    .A2(_04418_));
 sg13g2_a221oi_1 _25882_ (.B2(_04419_),
    .C1(_04382_),
    .B1(_04397_),
    .A1(_10404_),
    .Y(_04420_),
    .A2(\soc_I.clint_I.mtimecmp[57] ));
 sg13g2_nor2b_1 _25883_ (.A(_04379_),
    .B_N(_04381_),
    .Y(_04421_));
 sg13g2_nor3_1 _25884_ (.A(_04395_),
    .B(_04420_),
    .C(_04421_),
    .Y(_04422_));
 sg13g2_nor2_1 _25885_ (.A(_04385_),
    .B(_04422_),
    .Y(_04423_));
 sg13g2_a221oi_1 _25886_ (.B2(_04387_),
    .C1(_04423_),
    .B1(_04383_),
    .A1(\soc_I.clint_I.mtime[63] ),
    .Y(_04424_),
    .A2(_10572_));
 sg13g2_a21oi_2 _25887_ (.B1(net9011),
    .Y(_01002_),
    .A2(_04424_),
    .A1(_04412_));
 sg13g2_a22oi_1 _25888_ (.Y(_04425_),
    .B1(net8122),
    .B2(net3037),
    .A2(net8806),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[0] ));
 sg13g2_nor2_1 _25889_ (.A(net9037),
    .B(net3038),
    .Y(_01003_));
 sg13g2_a22oi_1 _25890_ (.Y(_04426_),
    .B1(net8122),
    .B2(net2807),
    .A2(net8806),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[1] ));
 sg13g2_nor2_1 _25891_ (.A(net9039),
    .B(net2808),
    .Y(_01004_));
 sg13g2_nor2b_1 _25892_ (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[0] ),
    .B_N(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[1] ),
    .Y(_04427_));
 sg13g2_nand2_1 _25893_ (.Y(_04428_),
    .A(_04078_),
    .B(net8945));
 sg13g2_nand2_1 _25894_ (.Y(_04429_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[2] ),
    .B(_04078_));
 sg13g2_xnor2_1 _25895_ (.Y(_04430_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[2] ),
    .B(_04428_));
 sg13g2_nand2_1 _25896_ (.Y(_04431_),
    .A(net8354),
    .B(_04430_));
 sg13g2_a22oi_1 _25897_ (.Y(_04432_),
    .B1(net8122),
    .B2(net4321),
    .A2(net8806),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[2] ));
 sg13g2_a21oi_1 _25898_ (.A1(_04431_),
    .A2(net4322),
    .Y(_01005_),
    .B1(net9046));
 sg13g2_and2_1 _25899_ (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[3] ),
    .B(_04082_),
    .X(_04433_));
 sg13g2_xnor2_1 _25900_ (.Y(_04434_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[3] ),
    .B(_04082_));
 sg13g2_nor2_1 _25901_ (.A(_04429_),
    .B(_04434_),
    .Y(_04435_));
 sg13g2_xor2_1 _25902_ (.B(_04434_),
    .A(_04429_),
    .X(_04436_));
 sg13g2_nor2b_1 _25903_ (.A(net8945),
    .B_N(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[3] ),
    .Y(_04437_));
 sg13g2_a21oi_1 _25904_ (.A1(net8945),
    .A2(_04436_),
    .Y(_04438_),
    .B1(_04437_));
 sg13g2_o21ai_1 _25905_ (.B1(net9372),
    .Y(_04439_),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[3] ),
    .A2(_04252_));
 sg13g2_a221oi_1 _25906_ (.B2(net8356),
    .C1(_04439_),
    .B1(_04438_),
    .A1(_10555_),
    .Y(_01006_),
    .A2(net8122));
 sg13g2_nand2_1 _25907_ (.Y(_04440_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[4] ),
    .B(_04086_));
 sg13g2_xor2_1 _25908_ (.B(_04086_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[4] ),
    .X(_04441_));
 sg13g2_o21ai_1 _25909_ (.B1(_04441_),
    .Y(_04442_),
    .A1(_04433_),
    .A2(_04435_));
 sg13g2_or3_1 _25910_ (.A(_04433_),
    .B(_04435_),
    .C(_04441_),
    .X(_04443_));
 sg13g2_nand2_1 _25911_ (.Y(_04444_),
    .A(_04442_),
    .B(_04443_));
 sg13g2_o21ai_1 _25912_ (.B1(net8354),
    .Y(_04445_),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[4] ),
    .A2(net8945));
 sg13g2_a21oi_1 _25913_ (.A1(net8945),
    .A2(_04444_),
    .Y(_04446_),
    .B1(_04445_));
 sg13g2_a221oi_1 _25914_ (.B2(net4847),
    .C1(_04446_),
    .B1(net8122),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[4] ),
    .Y(_04447_),
    .A2(net8806));
 sg13g2_nor2_1 _25915_ (.A(net9046),
    .B(net4848),
    .Y(_01007_));
 sg13g2_xnor2_1 _25916_ (.Y(_04448_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[5] ),
    .B(_03819_));
 sg13g2_a21oi_1 _25917_ (.A1(_04440_),
    .A2(_04442_),
    .Y(_04449_),
    .B1(_04448_));
 sg13g2_and3_1 _25918_ (.X(_04450_),
    .A(_04440_),
    .B(_04442_),
    .C(_04448_));
 sg13g2_o21ai_1 _25919_ (.B1(_04427_),
    .Y(_04451_),
    .A1(_04449_),
    .A2(_04450_));
 sg13g2_o21ai_1 _25920_ (.B1(_04451_),
    .Y(_04452_),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[5] ),
    .A2(net8945));
 sg13g2_a22oi_1 _25921_ (.Y(_04453_),
    .B1(net8122),
    .B2(net5422),
    .A2(net8806),
    .A1(net4695));
 sg13g2_o21ai_1 _25922_ (.B1(_04453_),
    .Y(_04454_),
    .A1(net8370),
    .A2(_04452_));
 sg13g2_and2_1 _25923_ (.A(net9376),
    .B(net5423),
    .X(_01008_));
 sg13g2_a21o_1 _25924_ (.A2(_03819_),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[5] ),
    .B1(_04449_),
    .X(_04455_));
 sg13g2_and3_2 _25925_ (.X(_04456_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[6] ),
    .B(net8945),
    .C(_04455_));
 sg13g2_a21oi_1 _25926_ (.A1(net8945),
    .A2(_04455_),
    .Y(_04457_),
    .B1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[6] ));
 sg13g2_or3_1 _25927_ (.A(net8370),
    .B(_04456_),
    .C(_04457_),
    .X(_04458_));
 sg13g2_a22oi_1 _25928_ (.Y(_04459_),
    .B1(net8122),
    .B2(net3923),
    .A2(net8806),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[6] ));
 sg13g2_a21oi_1 _25929_ (.A1(_04458_),
    .A2(net3924),
    .Y(_01009_),
    .B1(net9046));
 sg13g2_o21ai_1 _25930_ (.B1(net8350),
    .Y(_04460_),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[7] ),
    .A2(_04456_));
 sg13g2_a21o_1 _25931_ (.A2(_04456_),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[7] ),
    .B1(_04460_),
    .X(_04461_));
 sg13g2_a22oi_1 _25932_ (.Y(_04462_),
    .B1(net8120),
    .B2(net4228),
    .A2(net8804),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[7] ));
 sg13g2_a21oi_1 _25933_ (.A1(_04461_),
    .A2(net4229),
    .Y(_01010_),
    .B1(net9023));
 sg13g2_and3_1 _25934_ (.X(_04463_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[8] ),
    .B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[7] ),
    .C(_04456_));
 sg13g2_a21oi_1 _25935_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[7] ),
    .A2(_04456_),
    .Y(_04464_),
    .B1(net4957));
 sg13g2_nor3_1 _25936_ (.A(net8362),
    .B(_04463_),
    .C(_04464_),
    .Y(_04465_));
 sg13g2_a221oi_1 _25937_ (.B2(net5233),
    .C1(_04465_),
    .B1(net8120),
    .A1(net4670),
    .Y(_04466_),
    .A2(net8801));
 sg13g2_nor2_1 _25938_ (.A(net9024),
    .B(_04466_),
    .Y(_01011_));
 sg13g2_and2_1 _25939_ (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[9] ),
    .B(_04463_),
    .X(_04467_));
 sg13g2_o21ai_1 _25940_ (.B1(net8349),
    .Y(_04468_),
    .A1(net5027),
    .A2(_04463_));
 sg13g2_a22oi_1 _25941_ (.Y(_04469_),
    .B1(net8120),
    .B2(net5330),
    .A2(net8801),
    .A1(net4780));
 sg13g2_o21ai_1 _25942_ (.B1(_04469_),
    .Y(_04470_),
    .A1(_04467_),
    .A2(_04468_));
 sg13g2_and2_1 _25943_ (.A(net9352),
    .B(_04470_),
    .X(_01012_));
 sg13g2_and2_1 _25944_ (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[10] ),
    .B(_04467_),
    .X(_04471_));
 sg13g2_nor2_1 _25945_ (.A(net8361),
    .B(_04471_),
    .Y(_04472_));
 sg13g2_o21ai_1 _25946_ (.B1(_04472_),
    .Y(_04473_),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[10] ),
    .A2(_04467_));
 sg13g2_a22oi_1 _25947_ (.Y(_04474_),
    .B1(net8120),
    .B2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[10] ),
    .A2(net8801),
    .A1(net4055));
 sg13g2_a21oi_1 _25948_ (.A1(_04473_),
    .A2(net4056),
    .Y(_01013_),
    .B1(net9023));
 sg13g2_and2_1 _25949_ (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[11] ),
    .B(_04471_),
    .X(_04475_));
 sg13g2_nor2_1 _25950_ (.A(net8361),
    .B(_04475_),
    .Y(_04476_));
 sg13g2_o21ai_1 _25951_ (.B1(_04476_),
    .Y(_04477_),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[11] ),
    .A2(_04471_));
 sg13g2_a22oi_1 _25952_ (.Y(_04478_),
    .B1(net8120),
    .B2(net4177),
    .A2(net8804),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[11] ));
 sg13g2_a21oi_1 _25953_ (.A1(_04477_),
    .A2(net4178),
    .Y(_01014_),
    .B1(net9026));
 sg13g2_and2_1 _25954_ (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[12] ),
    .B(_04475_),
    .X(_04479_));
 sg13g2_nor2_1 _25955_ (.A(net8361),
    .B(_04479_),
    .Y(_04480_));
 sg13g2_o21ai_1 _25956_ (.B1(_04480_),
    .Y(_04481_),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[12] ),
    .A2(_04475_));
 sg13g2_a22oi_1 _25957_ (.Y(_04482_),
    .B1(net8120),
    .B2(net4133),
    .A2(net8801),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[12] ));
 sg13g2_a21oi_1 _25958_ (.A1(_04481_),
    .A2(net4134),
    .Y(_01015_),
    .B1(net9025));
 sg13g2_and2_1 _25959_ (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[13] ),
    .B(_04479_),
    .X(_04483_));
 sg13g2_nor2_1 _25960_ (.A(net8363),
    .B(_04483_),
    .Y(_04484_));
 sg13g2_o21ai_1 _25961_ (.B1(_04484_),
    .Y(_04485_),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[13] ),
    .A2(_04479_));
 sg13g2_a22oi_1 _25962_ (.Y(_04486_),
    .B1(net8119),
    .B2(net4123),
    .A2(net8802),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[13] ));
 sg13g2_a21oi_1 _25963_ (.A1(_04485_),
    .A2(net4124),
    .Y(_01016_),
    .B1(net9031));
 sg13g2_and2_1 _25964_ (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[14] ),
    .B(_04483_),
    .X(_04487_));
 sg13g2_nor2_1 _25965_ (.A(net8363),
    .B(_04487_),
    .Y(_04488_));
 sg13g2_o21ai_1 _25966_ (.B1(_04488_),
    .Y(_04489_),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[14] ),
    .A2(_04483_));
 sg13g2_a22oi_1 _25967_ (.Y(_04490_),
    .B1(net8119),
    .B2(net4338),
    .A2(net8802),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[14] ));
 sg13g2_a21oi_1 _25968_ (.A1(_04489_),
    .A2(net4339),
    .Y(_01017_),
    .B1(net9029));
 sg13g2_and2_1 _25969_ (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[15] ),
    .B(_04487_),
    .X(_04491_));
 sg13g2_nor2_1 _25970_ (.A(net8363),
    .B(_04491_),
    .Y(_04492_));
 sg13g2_o21ai_1 _25971_ (.B1(_04492_),
    .Y(_04493_),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[15] ),
    .A2(_04487_));
 sg13g2_a22oi_1 _25972_ (.Y(_04494_),
    .B1(net8119),
    .B2(net4139),
    .A2(net8802),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[15] ));
 sg13g2_a21oi_1 _25973_ (.A1(_04493_),
    .A2(net4140),
    .Y(_01018_),
    .B1(net9029));
 sg13g2_and2_1 _25974_ (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[16] ),
    .B(_04491_),
    .X(_04495_));
 sg13g2_nor2_1 _25975_ (.A(net8363),
    .B(_04495_),
    .Y(_04496_));
 sg13g2_o21ai_1 _25976_ (.B1(_04496_),
    .Y(_04497_),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[16] ),
    .A2(_04491_));
 sg13g2_a22oi_1 _25977_ (.Y(_04498_),
    .B1(net8119),
    .B2(net4203),
    .A2(net8802),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[16] ));
 sg13g2_a21oi_1 _25978_ (.A1(_04497_),
    .A2(net4204),
    .Y(_01019_),
    .B1(net9029));
 sg13g2_and2_1 _25979_ (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[17] ),
    .B(_04495_),
    .X(_04499_));
 sg13g2_nor2_1 _25980_ (.A(net8364),
    .B(_04499_),
    .Y(_04500_));
 sg13g2_o21ai_1 _25981_ (.B1(_04500_),
    .Y(_04501_),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[17] ),
    .A2(_04495_));
 sg13g2_a22oi_1 _25982_ (.Y(_04502_),
    .B1(net8119),
    .B2(net4246),
    .A2(net8802),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[17] ));
 sg13g2_a21oi_1 _25983_ (.A1(_04501_),
    .A2(net4247),
    .Y(_01020_),
    .B1(net9027));
 sg13g2_and2_1 _25984_ (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[18] ),
    .B(_04499_),
    .X(_04503_));
 sg13g2_nor2_1 _25985_ (.A(net8364),
    .B(_04503_),
    .Y(_04504_));
 sg13g2_o21ai_1 _25986_ (.B1(_04504_),
    .Y(_04505_),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[18] ),
    .A2(_04499_));
 sg13g2_a22oi_1 _25987_ (.Y(_04506_),
    .B1(net8119),
    .B2(net4415),
    .A2(net8802),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[18] ));
 sg13g2_a21oi_1 _25988_ (.A1(_04505_),
    .A2(net4416),
    .Y(_01021_),
    .B1(net9027));
 sg13g2_and2_2 _25989_ (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[19] ),
    .B(_04503_),
    .X(_04507_));
 sg13g2_nor2_1 _25990_ (.A(net8364),
    .B(_04507_),
    .Y(_04508_));
 sg13g2_o21ai_1 _25991_ (.B1(_04508_),
    .Y(_04509_),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[19] ),
    .A2(_04503_));
 sg13g2_a22oi_1 _25992_ (.Y(_04510_),
    .B1(net8119),
    .B2(net4550),
    .A2(net8802),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[19] ));
 sg13g2_a21oi_1 _25993_ (.A1(_04509_),
    .A2(net4551),
    .Y(_01022_),
    .B1(net9027));
 sg13g2_and2_2 _25994_ (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[20] ),
    .B(_04507_),
    .X(_04511_));
 sg13g2_nor2_1 _25995_ (.A(net8369),
    .B(_04511_),
    .Y(_04512_));
 sg13g2_o21ai_1 _25996_ (.B1(_04512_),
    .Y(_04513_),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[20] ),
    .A2(_04507_));
 sg13g2_a22oi_1 _25997_ (.Y(_04514_),
    .B1(net8123),
    .B2(net4232),
    .A2(net8806),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[20] ));
 sg13g2_a21oi_1 _25998_ (.A1(_04513_),
    .A2(net4233),
    .Y(_01023_),
    .B1(net9045));
 sg13g2_and2_1 _25999_ (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[21] ),
    .B(_04511_),
    .X(_04515_));
 sg13g2_nor2_1 _26000_ (.A(net8368),
    .B(_04515_),
    .Y(_04516_));
 sg13g2_o21ai_1 _26001_ (.B1(_04516_),
    .Y(_04517_),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[21] ),
    .A2(_04511_));
 sg13g2_a22oi_1 _26002_ (.Y(_04518_),
    .B1(net8123),
    .B2(net3968),
    .A2(net8805),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[21] ));
 sg13g2_a21oi_1 _26003_ (.A1(_04517_),
    .A2(net3969),
    .Y(_01024_),
    .B1(net9052));
 sg13g2_and2_1 _26004_ (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[22] ),
    .B(_04515_),
    .X(_04519_));
 sg13g2_nor2_1 _26005_ (.A(net8368),
    .B(_04519_),
    .Y(_04520_));
 sg13g2_o21ai_1 _26006_ (.B1(_04520_),
    .Y(_04521_),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[22] ),
    .A2(_04515_));
 sg13g2_a22oi_1 _26007_ (.Y(_04522_),
    .B1(net8123),
    .B2(net4403),
    .A2(net8807),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[22] ));
 sg13g2_a21oi_1 _26008_ (.A1(_04521_),
    .A2(net4404),
    .Y(_01025_),
    .B1(net9051));
 sg13g2_and2_1 _26009_ (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[23] ),
    .B(_04519_),
    .X(_04523_));
 sg13g2_nor2_1 _26010_ (.A(net8367),
    .B(_04523_),
    .Y(_04524_));
 sg13g2_o21ai_1 _26011_ (.B1(_04524_),
    .Y(_04525_),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[23] ),
    .A2(_04519_));
 sg13g2_a22oi_1 _26012_ (.Y(_04526_),
    .B1(net8123),
    .B2(net4422),
    .A2(net8805),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[23] ));
 sg13g2_a21oi_1 _26013_ (.A1(_04525_),
    .A2(net4423),
    .Y(_01026_),
    .B1(net9044));
 sg13g2_and2_1 _26014_ (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[24] ),
    .B(_04523_),
    .X(_04527_));
 sg13g2_nor2_1 _26015_ (.A(net8367),
    .B(_04527_),
    .Y(_04528_));
 sg13g2_o21ai_1 _26016_ (.B1(_04528_),
    .Y(_04529_),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[24] ),
    .A2(_04523_));
 sg13g2_a22oi_1 _26017_ (.Y(_04530_),
    .B1(net8122),
    .B2(net4119),
    .A2(net8805),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[24] ));
 sg13g2_a21oi_1 _26018_ (.A1(_04529_),
    .A2(net4120),
    .Y(_01027_),
    .B1(net9050));
 sg13g2_and2_1 _26019_ (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[25] ),
    .B(_04527_),
    .X(_04531_));
 sg13g2_nor2_1 _26020_ (.A(net8367),
    .B(_04531_),
    .Y(_04532_));
 sg13g2_o21ai_1 _26021_ (.B1(_04532_),
    .Y(_04533_),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[25] ),
    .A2(_04527_));
 sg13g2_a22oi_1 _26022_ (.Y(_04534_),
    .B1(net8123),
    .B2(net4086),
    .A2(net8805),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[25] ));
 sg13g2_a21oi_1 _26023_ (.A1(_04533_),
    .A2(net4087),
    .Y(_01028_),
    .B1(net9050));
 sg13g2_and2_2 _26024_ (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[26] ),
    .B(_04531_),
    .X(_04535_));
 sg13g2_nor2_1 _26025_ (.A(net8368),
    .B(_04535_),
    .Y(_04536_));
 sg13g2_o21ai_1 _26026_ (.B1(_04536_),
    .Y(_04537_),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[26] ),
    .A2(_04531_));
 sg13g2_a22oi_1 _26027_ (.Y(_04538_),
    .B1(net8123),
    .B2(net4263),
    .A2(net8805),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[26] ));
 sg13g2_a21oi_1 _26028_ (.A1(_04537_),
    .A2(net4264),
    .Y(_01029_),
    .B1(net9051));
 sg13g2_and2_1 _26029_ (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[27] ),
    .B(_04535_),
    .X(_04539_));
 sg13g2_nor2_1 _26030_ (.A(net8805),
    .B(_04539_),
    .Y(_04540_));
 sg13g2_o21ai_1 _26031_ (.B1(_04540_),
    .Y(_04541_),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[27] ),
    .A2(_04535_));
 sg13g2_a21oi_1 _26032_ (.A1(net4801),
    .A2(net8805),
    .Y(_04542_),
    .B1(net8123));
 sg13g2_o21ai_1 _26033_ (.B1(net9383),
    .Y(_04543_),
    .A1(net4963),
    .A2(_04254_));
 sg13g2_a21oi_1 _26034_ (.A1(_04541_),
    .A2(_04542_),
    .Y(_01030_),
    .B1(_04543_));
 sg13g2_and2_1 _26035_ (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[28] ),
    .B(_04539_),
    .X(_04544_));
 sg13g2_nor2_1 _26036_ (.A(net8365),
    .B(_04544_),
    .Y(_04545_));
 sg13g2_o21ai_1 _26037_ (.B1(_04545_),
    .Y(_04546_),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[28] ),
    .A2(_04539_));
 sg13g2_a22oi_1 _26038_ (.Y(_04547_),
    .B1(net8121),
    .B2(net4690),
    .A2(net8803),
    .A1(net4397));
 sg13g2_a21oi_1 _26039_ (.A1(_04546_),
    .A2(_04547_),
    .Y(_01031_),
    .B1(net9041));
 sg13g2_and2_1 _26040_ (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[29] ),
    .B(_04544_),
    .X(_04548_));
 sg13g2_nor2_1 _26041_ (.A(net8802),
    .B(_04548_),
    .Y(_04549_));
 sg13g2_o21ai_1 _26042_ (.B1(_04549_),
    .Y(_04550_),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[29] ),
    .A2(_04544_));
 sg13g2_a21oi_1 _26043_ (.A1(net4874),
    .A2(net8803),
    .Y(_04551_),
    .B1(net8121));
 sg13g2_o21ai_1 _26044_ (.B1(net9383),
    .Y(_04552_),
    .A1(net4672),
    .A2(_04254_));
 sg13g2_a21oi_1 _26045_ (.A1(_04550_),
    .A2(_04551_),
    .Y(_01032_),
    .B1(_04552_));
 sg13g2_and2_1 _26046_ (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[30] ),
    .B(_04548_),
    .X(_04553_));
 sg13g2_nor2_1 _26047_ (.A(net8365),
    .B(_04553_),
    .Y(_04554_));
 sg13g2_o21ai_1 _26048_ (.B1(_04554_),
    .Y(_04555_),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[30] ),
    .A2(_04548_));
 sg13g2_a22oi_1 _26049_ (.Y(_04556_),
    .B1(net8121),
    .B2(net3885),
    .A2(net8803),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[30] ));
 sg13g2_a21oi_1 _26050_ (.A1(_04555_),
    .A2(net3886),
    .Y(_01033_),
    .B1(net9040));
 sg13g2_a21oi_1 _26051_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[31] ),
    .A2(_04553_),
    .Y(_04557_),
    .B1(net8365));
 sg13g2_o21ai_1 _26052_ (.B1(_04557_),
    .Y(_04558_),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[31] ),
    .A2(_04553_));
 sg13g2_a22oi_1 _26053_ (.Y(_04559_),
    .B1(net8119),
    .B2(net4790),
    .A2(net8803),
    .A1(net4406));
 sg13g2_a21oi_1 _26054_ (.A1(_04558_),
    .A2(_04559_),
    .Y(_01034_),
    .B1(net9031));
 sg13g2_and2_1 _26055_ (.A(net7790),
    .B(net7992),
    .X(_04560_));
 sg13g2_o21ai_1 _26056_ (.B1(net9382),
    .Y(_04561_),
    .A1(net4350),
    .A2(net7718));
 sg13g2_a21oi_1 _26057_ (.A1(_03841_),
    .A2(net7718),
    .Y(_01035_),
    .B1(_04561_));
 sg13g2_o21ai_1 _26058_ (.B1(net9372),
    .Y(_04562_),
    .A1(net4231),
    .A2(net7721));
 sg13g2_a21oi_1 _26059_ (.A1(_03862_),
    .A2(net7721),
    .Y(_01036_),
    .B1(_04562_));
 sg13g2_o21ai_1 _26060_ (.B1(net9379),
    .Y(_04563_),
    .A1(net4540),
    .A2(net7721));
 sg13g2_a21oi_1 _26061_ (.A1(_03871_),
    .A2(net7721),
    .Y(_01037_),
    .B1(_04563_));
 sg13g2_o21ai_1 _26062_ (.B1(net9372),
    .Y(_04564_),
    .A1(net5140),
    .A2(net7713));
 sg13g2_a21oi_1 _26063_ (.A1(_03880_),
    .A2(net7713),
    .Y(_01038_),
    .B1(_04564_));
 sg13g2_o21ai_1 _26064_ (.B1(net9376),
    .Y(_04565_),
    .A1(net4794),
    .A2(net7721));
 sg13g2_a21oi_1 _26065_ (.A1(_03889_),
    .A2(net7721),
    .Y(_01039_),
    .B1(_04565_));
 sg13g2_o21ai_1 _26066_ (.B1(net9370),
    .Y(_04566_),
    .A1(net4320),
    .A2(net7713));
 sg13g2_a21oi_1 _26067_ (.A1(_03896_),
    .A2(net7713),
    .Y(_01040_),
    .B1(_04566_));
 sg13g2_o21ai_1 _26068_ (.B1(net9395),
    .Y(_04567_),
    .A1(net4773),
    .A2(net7721));
 sg13g2_a21oi_1 _26069_ (.A1(_03904_),
    .A2(net7721),
    .Y(_01041_),
    .B1(_04567_));
 sg13g2_o21ai_1 _26070_ (.B1(net9349),
    .Y(_04568_),
    .A1(net5088),
    .A2(net7713));
 sg13g2_a21oi_1 _26071_ (.A1(_03913_),
    .A2(net7713),
    .Y(_01042_),
    .B1(_04568_));
 sg13g2_o21ai_1 _26072_ (.B1(net9352),
    .Y(_04569_),
    .A1(net4700),
    .A2(net7713));
 sg13g2_a21oi_1 _26073_ (.A1(_03921_),
    .A2(net7713),
    .Y(_01043_),
    .B1(_04569_));
 sg13g2_o21ai_1 _26074_ (.B1(net9352),
    .Y(_04570_),
    .A1(net4394),
    .A2(net7714));
 sg13g2_a21oi_1 _26075_ (.A1(_03927_),
    .A2(net7714),
    .Y(_01044_),
    .B1(_04570_));
 sg13g2_o21ai_1 _26076_ (.B1(net9353),
    .Y(_04571_),
    .A1(net4402),
    .A2(net7714));
 sg13g2_a21oi_1 _26077_ (.A1(_03933_),
    .A2(net7714),
    .Y(_01045_),
    .B1(_04571_));
 sg13g2_o21ai_1 _26078_ (.B1(net9348),
    .Y(_04572_),
    .A1(net4447),
    .A2(net7718));
 sg13g2_a21oi_1 _26079_ (.A1(_03940_),
    .A2(net7714),
    .Y(_01046_),
    .B1(_04572_));
 sg13g2_o21ai_1 _26080_ (.B1(net9362),
    .Y(_04573_),
    .A1(net4586),
    .A2(net7714));
 sg13g2_a21oi_1 _26081_ (.A1(_03946_),
    .A2(net7714),
    .Y(_01047_),
    .B1(_04573_));
 sg13g2_o21ai_1 _26082_ (.B1(net9354),
    .Y(_04574_),
    .A1(net4482),
    .A2(net7715));
 sg13g2_a21oi_1 _26083_ (.A1(_03952_),
    .A2(net7715),
    .Y(_01048_),
    .B1(_04574_));
 sg13g2_o21ai_1 _26084_ (.B1(net9356),
    .Y(_04575_),
    .A1(net4429),
    .A2(net7715));
 sg13g2_a21oi_1 _26085_ (.A1(_03958_),
    .A2(net7715),
    .Y(_01049_),
    .B1(_04575_));
 sg13g2_o21ai_1 _26086_ (.B1(net9354),
    .Y(_04576_),
    .A1(net4521),
    .A2(net7715));
 sg13g2_a21oi_1 _26087_ (.A1(_03964_),
    .A2(net7715),
    .Y(_01050_),
    .B1(_04576_));
 sg13g2_o21ai_1 _26088_ (.B1(net9357),
    .Y(_04577_),
    .A1(net4303),
    .A2(net7715));
 sg13g2_a21oi_1 _26089_ (.A1(_03971_),
    .A2(net7715),
    .Y(_01051_),
    .B1(_04577_));
 sg13g2_o21ai_1 _26090_ (.B1(net9358),
    .Y(_04578_),
    .A1(net4549),
    .A2(net7716));
 sg13g2_a21oi_1 _26091_ (.A1(_03980_),
    .A2(net7716),
    .Y(_01052_),
    .B1(_04578_));
 sg13g2_o21ai_1 _26092_ (.B1(net9360),
    .Y(_04579_),
    .A1(net4493),
    .A2(net7716));
 sg13g2_a21oi_1 _26093_ (.A1(_03987_),
    .A2(net7716),
    .Y(_01053_),
    .B1(_04579_));
 sg13g2_o21ai_1 _26094_ (.B1(net9358),
    .Y(_04580_),
    .A1(net4581),
    .A2(net7716));
 sg13g2_a21oi_1 _26095_ (.A1(_03995_),
    .A2(net7716),
    .Y(_01054_),
    .B1(_04580_));
 sg13g2_o21ai_1 _26096_ (.B1(net9365),
    .Y(_04581_),
    .A1(net4337),
    .A2(net7716));
 sg13g2_a21oi_1 _26097_ (.A1(_04002_),
    .A2(net7716),
    .Y(_01055_),
    .B1(_04581_));
 sg13g2_o21ai_1 _26098_ (.B1(net9401),
    .Y(_04582_),
    .A1(net4756),
    .A2(net7720));
 sg13g2_a21oi_1 _26099_ (.A1(_04008_),
    .A2(net7720),
    .Y(_01056_),
    .B1(_04582_));
 sg13g2_o21ai_1 _26100_ (.B1(net9402),
    .Y(_04583_),
    .A1(net4631),
    .A2(net7720));
 sg13g2_a21oi_1 _26101_ (.A1(_04014_),
    .A2(net7720),
    .Y(_01057_),
    .B1(_04583_));
 sg13g2_o21ai_1 _26102_ (.B1(net9385),
    .Y(_04584_),
    .A1(net4290),
    .A2(net7719));
 sg13g2_a21oi_1 _26103_ (.A1(_04020_),
    .A2(net7719),
    .Y(_01058_),
    .B1(_04584_));
 sg13g2_o21ai_1 _26104_ (.B1(net9390),
    .Y(_04585_),
    .A1(net4446),
    .A2(net7719));
 sg13g2_a21oi_1 _26105_ (.A1(_04027_),
    .A2(net7719),
    .Y(_01059_),
    .B1(_04585_));
 sg13g2_o21ai_1 _26106_ (.B1(net9390),
    .Y(_04586_),
    .A1(net4629),
    .A2(net7720));
 sg13g2_a21oi_1 _26107_ (.A1(_04033_),
    .A2(net7720),
    .Y(_01060_),
    .B1(_04586_));
 sg13g2_o21ai_1 _26108_ (.B1(net9404),
    .Y(_04587_),
    .A1(net4654),
    .A2(net7719));
 sg13g2_a21oi_1 _26109_ (.A1(_04039_),
    .A2(net7719),
    .Y(_01061_),
    .B1(_04587_));
 sg13g2_o21ai_1 _26110_ (.B1(net9383),
    .Y(_04588_),
    .A1(net4400),
    .A2(net7719));
 sg13g2_a21oi_1 _26111_ (.A1(_04045_),
    .A2(net7719),
    .Y(_01062_),
    .B1(_04588_));
 sg13g2_o21ai_1 _26112_ (.B1(net9384),
    .Y(_04589_),
    .A1(net4463),
    .A2(net7717));
 sg13g2_a21oi_1 _26113_ (.A1(_04052_),
    .A2(net7717),
    .Y(_01063_),
    .B1(_04589_));
 sg13g2_o21ai_1 _26114_ (.B1(net9383),
    .Y(_04590_),
    .A1(net4355),
    .A2(net7718));
 sg13g2_a21oi_1 _26115_ (.A1(_04058_),
    .A2(net7718),
    .Y(_01064_),
    .B1(_04590_));
 sg13g2_o21ai_1 _26116_ (.B1(net9366),
    .Y(_04591_),
    .A1(net4428),
    .A2(net7717));
 sg13g2_a21oi_1 _26117_ (.A1(_04064_),
    .A2(net7717),
    .Y(_01065_),
    .B1(_04591_));
 sg13g2_o21ai_1 _26118_ (.B1(net9382),
    .Y(_04592_),
    .A1(net4481),
    .A2(net7717));
 sg13g2_a21oi_1 _26119_ (.A1(_04070_),
    .A2(net7717),
    .Y(_01066_),
    .B1(_04592_));
 sg13g2_and2_1 _26120_ (.A(net7929),
    .B(net7993),
    .X(_04593_));
 sg13g2_nand2_1 _26121_ (.Y(_04594_),
    .A(net7927),
    .B(net7990));
 sg13g2_nor2_2 _26122_ (.A(_04254_),
    .B(net7762),
    .Y(_04595_));
 sg13g2_a22oi_1 _26123_ (.Y(_04596_),
    .B1(_04595_),
    .B2(net5452),
    .A2(net8801),
    .A1(net4221));
 sg13g2_o21ai_1 _26124_ (.B1(_04596_),
    .Y(_04597_),
    .A1(_03880_),
    .A2(_04594_));
 sg13g2_and2_1 _26125_ (.A(net9374),
    .B(_04597_),
    .X(_01067_));
 sg13g2_o21ai_1 _26126_ (.B1(_04594_),
    .Y(_04598_),
    .A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[3] ),
    .A2(net8361));
 sg13g2_a221oi_1 _26127_ (.B2(_03915_),
    .C1(net9025),
    .B1(_04598_),
    .A1(_10554_),
    .Y(_01068_),
    .A2(_04595_));
 sg13g2_a21oi_1 _26128_ (.A1(net4559),
    .A2(net8349),
    .Y(_04599_),
    .B1(_03941_));
 sg13g2_nor3_1 _26129_ (.A(net8801),
    .B(_04595_),
    .C(_04599_),
    .Y(_04600_));
 sg13g2_a21oi_1 _26130_ (.A1(net5266),
    .A2(_04595_),
    .Y(_04601_),
    .B1(_04600_));
 sg13g2_nand2_1 _26131_ (.Y(_01069_),
    .A(net9350),
    .B(_04601_));
 sg13g2_a21oi_1 _26132_ (.A1(\soc_I.kianv_I.control_unit_I.main_fsm_I.privilege_mode[1] ),
    .A2(net8350),
    .Y(_04602_),
    .B1(_03947_));
 sg13g2_nor3_1 _26133_ (.A(net8801),
    .B(_04595_),
    .C(_04602_),
    .Y(_04603_));
 sg13g2_a21oi_1 _26134_ (.A1(net4745),
    .A2(_04595_),
    .Y(_04604_),
    .B1(_04603_));
 sg13g2_nand2_1 _26135_ (.Y(_01070_),
    .A(net9350),
    .B(net4746));
 sg13g2_nor2_1 _26136_ (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[11] ),
    .B(_04252_),
    .Y(_04605_));
 sg13g2_nor2_1 _26137_ (.A(net4559),
    .B(_04254_),
    .Y(_04606_));
 sg13g2_o21ai_1 _26138_ (.B1(net9374),
    .Y(_01071_),
    .A1(_04605_),
    .A2(_04606_));
 sg13g2_nand2_1 _26139_ (.Y(_04607_),
    .A(net4745),
    .B(net8801));
 sg13g2_a21oi_1 _26140_ (.A1(net4782),
    .A2(_04252_),
    .Y(_04608_),
    .B1(net9037));
 sg13g2_nand3_1 _26141_ (.B(_04607_),
    .C(_04608_),
    .A(net8361),
    .Y(_01072_));
 sg13g2_nand2_1 _26142_ (.Y(_04609_),
    .A(_02798_),
    .B(_02805_));
 sg13g2_nand2_1 _26143_ (.Y(_04610_),
    .A(net2651),
    .B(net8593));
 sg13g2_o21ai_1 _26144_ (.B1(_04610_),
    .Y(_01073_),
    .A1(net9170),
    .A2(net8593));
 sg13g2_mux2_1 _26145_ (.A0(\soc_I.rx_uart_i.fifo_i.din[1] ),
    .A1(net4180),
    .S(net8593),
    .X(_01074_));
 sg13g2_mux2_1 _26146_ (.A0(net3981),
    .A1(net4071),
    .S(_04609_),
    .X(_01075_));
 sg13g2_mux2_1 _26147_ (.A0(net9284),
    .A1(net4158),
    .S(net8593),
    .X(_01076_));
 sg13g2_mux2_1 _26148_ (.A0(\soc_I.rx_uart_i.fifo_i.din[4] ),
    .A1(net4003),
    .S(net8593),
    .X(_01077_));
 sg13g2_mux2_1 _26149_ (.A0(net9279),
    .A1(net4395),
    .S(net8593),
    .X(_01078_));
 sg13g2_mux2_1 _26150_ (.A0(net9278),
    .A1(net4207),
    .S(net8593),
    .X(_01079_));
 sg13g2_mux2_1 _26151_ (.A0(net9275),
    .A1(net4052),
    .S(net8593),
    .X(_01080_));
 sg13g2_nand2_1 _26152_ (.Y(_04611_),
    .A(_02798_),
    .B(_02801_));
 sg13g2_nand2_1 _26153_ (.Y(_04612_),
    .A(net2661),
    .B(net8543));
 sg13g2_o21ai_1 _26154_ (.B1(_04612_),
    .Y(_01081_),
    .A1(net9171),
    .A2(net8543));
 sg13g2_mux2_1 _26155_ (.A0(net9289),
    .A1(net4096),
    .S(net8543),
    .X(_01082_));
 sg13g2_mux2_1 _26156_ (.A0(net9286),
    .A1(net4194),
    .S(_04611_),
    .X(_01083_));
 sg13g2_mux2_1 _26157_ (.A0(net9284),
    .A1(net4152),
    .S(net8543),
    .X(_01084_));
 sg13g2_mux2_1 _26158_ (.A0(net9283),
    .A1(net3988),
    .S(net8543),
    .X(_01085_));
 sg13g2_mux2_1 _26159_ (.A0(net9279),
    .A1(net4063),
    .S(net8543),
    .X(_01086_));
 sg13g2_mux2_1 _26160_ (.A0(net9278),
    .A1(net4084),
    .S(net8543),
    .X(_01087_));
 sg13g2_mux2_1 _26161_ (.A0(net9275),
    .A1(net4163),
    .S(net8543),
    .X(_01088_));
 sg13g2_nand2_1 _26162_ (.Y(_04613_),
    .A(_02798_),
    .B(_02810_));
 sg13g2_nand2_1 _26163_ (.Y(_04614_),
    .A(net2716),
    .B(net8592));
 sg13g2_o21ai_1 _26164_ (.B1(_04614_),
    .Y(_01089_),
    .A1(net9170),
    .A2(net8592));
 sg13g2_mux2_1 _26165_ (.A0(net9289),
    .A1(net4034),
    .S(net8592),
    .X(_01090_));
 sg13g2_mux2_1 _26166_ (.A0(net9286),
    .A1(net4019),
    .S(_04613_),
    .X(_01091_));
 sg13g2_mux2_1 _26167_ (.A0(net9284),
    .A1(net4026),
    .S(net8592),
    .X(_01092_));
 sg13g2_mux2_1 _26168_ (.A0(net9283),
    .A1(net4094),
    .S(net8592),
    .X(_01093_));
 sg13g2_mux2_1 _26169_ (.A0(net9279),
    .A1(net4170),
    .S(net8592),
    .X(_01094_));
 sg13g2_mux2_1 _26170_ (.A0(net9278),
    .A1(net4131),
    .S(net8592),
    .X(_01095_));
 sg13g2_mux2_1 _26171_ (.A0(net9275),
    .A1(net4065),
    .S(net8592),
    .X(_01096_));
 sg13g2_nand3_1 _26172_ (.B(net9273),
    .C(_02805_),
    .A(\soc_I.rx_uart_i.fifo_i.wr_ptr[3] ),
    .Y(_04615_));
 sg13g2_nand2_1 _26173_ (.Y(_04616_),
    .A(net2760),
    .B(_04615_));
 sg13g2_o21ai_1 _26174_ (.B1(_04616_),
    .Y(_01097_),
    .A1(_10396_),
    .A2(_04615_));
 sg13g2_mux2_1 _26175_ (.A0(net9288),
    .A1(net4098),
    .S(net8591),
    .X(_01098_));
 sg13g2_mux2_1 _26176_ (.A0(net9287),
    .A1(net4286),
    .S(net8591),
    .X(_01099_));
 sg13g2_mux2_1 _26177_ (.A0(net9285),
    .A1(net4092),
    .S(net8591),
    .X(_01100_));
 sg13g2_mux2_1 _26178_ (.A0(net9282),
    .A1(net4089),
    .S(net8591),
    .X(_01101_));
 sg13g2_mux2_1 _26179_ (.A0(net9279),
    .A1(net4186),
    .S(net8591),
    .X(_01102_));
 sg13g2_mux2_1 _26180_ (.A0(net9277),
    .A1(net4043),
    .S(net8591),
    .X(_01103_));
 sg13g2_mux2_1 _26181_ (.A0(\soc_I.rx_uart_i.fifo_i.din[7] ),
    .A1(net3974),
    .S(net8591),
    .X(_01104_));
 sg13g2_nand2_2 _26182_ (.Y(_04617_),
    .A(_14165_),
    .B(_14302_));
 sg13g2_nand2_1 _26183_ (.Y(_04618_),
    .A(net3198),
    .B(net8117));
 sg13g2_o21ai_1 _26184_ (.B1(_04618_),
    .Y(_01105_),
    .A1(net7489),
    .A2(net8117));
 sg13g2_nand2_1 _26185_ (.Y(_04619_),
    .A(net3253),
    .B(net8117));
 sg13g2_o21ai_1 _26186_ (.B1(_04619_),
    .Y(_01106_),
    .A1(net7663),
    .A2(net8117));
 sg13g2_nand2_1 _26187_ (.Y(_04620_),
    .A(net3667),
    .B(net8117));
 sg13g2_o21ai_1 _26188_ (.B1(_04620_),
    .Y(_01107_),
    .A1(net7613),
    .A2(net8117));
 sg13g2_nand2_1 _26189_ (.Y(_04621_),
    .A(net3178),
    .B(net8115));
 sg13g2_o21ai_1 _26190_ (.B1(_04621_),
    .Y(_01108_),
    .A1(net7609),
    .A2(net8115));
 sg13g2_nand2_1 _26191_ (.Y(_04622_),
    .A(net3234),
    .B(net8112));
 sg13g2_o21ai_1 _26192_ (.B1(_04622_),
    .Y(_01109_),
    .A1(net7588),
    .A2(net8113));
 sg13g2_nand2_1 _26193_ (.Y(_04623_),
    .A(net3062),
    .B(net8112));
 sg13g2_o21ai_1 _26194_ (.B1(_04623_),
    .Y(_01110_),
    .A1(net7598),
    .A2(net8112));
 sg13g2_nand2_1 _26195_ (.Y(_04624_),
    .A(net3336),
    .B(net8114));
 sg13g2_o21ai_1 _26196_ (.B1(_04624_),
    .Y(_01111_),
    .A1(net7595),
    .A2(net8114));
 sg13g2_nand2_1 _26197_ (.Y(_04625_),
    .A(net3555),
    .B(net8108));
 sg13g2_o21ai_1 _26198_ (.B1(_04625_),
    .Y(_01112_),
    .A1(net7603),
    .A2(net8108));
 sg13g2_nand2_1 _26199_ (.Y(_04626_),
    .A(net3755),
    .B(net8113));
 sg13g2_o21ai_1 _26200_ (.B1(_04626_),
    .Y(_01113_),
    .A1(net7557),
    .A2(net8113));
 sg13g2_nand2_1 _26201_ (.Y(_04627_),
    .A(net2986),
    .B(net8116));
 sg13g2_o21ai_1 _26202_ (.B1(_04627_),
    .Y(_01114_),
    .A1(net7575),
    .A2(net8116));
 sg13g2_nand2_1 _26203_ (.Y(_04628_),
    .A(net3135),
    .B(net8114));
 sg13g2_o21ai_1 _26204_ (.B1(_04628_),
    .Y(_01115_),
    .A1(net7549),
    .A2(net8114));
 sg13g2_nand2_1 _26205_ (.Y(_04629_),
    .A(net3605),
    .B(net8108));
 sg13g2_o21ai_1 _26206_ (.B1(_04629_),
    .Y(_01116_),
    .A1(net7568),
    .A2(net8108));
 sg13g2_nand2_1 _26207_ (.Y(_04630_),
    .A(net3707),
    .B(net8114));
 sg13g2_o21ai_1 _26208_ (.B1(_04630_),
    .Y(_01117_),
    .A1(net7544),
    .A2(net8114));
 sg13g2_nand2_1 _26209_ (.Y(_04631_),
    .A(net3455),
    .B(net8116));
 sg13g2_o21ai_1 _26210_ (.B1(_04631_),
    .Y(_01118_),
    .A1(net7552),
    .A2(net8116));
 sg13g2_nand2_1 _26211_ (.Y(_04632_),
    .A(net3881),
    .B(net8111));
 sg13g2_o21ai_1 _26212_ (.B1(_04632_),
    .Y(_01119_),
    .A1(net7584),
    .A2(net8111));
 sg13g2_nand2_1 _26213_ (.Y(_04633_),
    .A(net3477),
    .B(net8109));
 sg13g2_o21ai_1 _26214_ (.B1(_04633_),
    .Y(_01120_),
    .A1(net7563),
    .A2(net8109));
 sg13g2_nand2_1 _26215_ (.Y(_04634_),
    .A(net3326),
    .B(net8108));
 sg13g2_o21ai_1 _26216_ (.B1(_04634_),
    .Y(_01121_),
    .A1(net7523),
    .A2(net8108));
 sg13g2_nand2_1 _26217_ (.Y(_04635_),
    .A(net2974),
    .B(net8108));
 sg13g2_o21ai_1 _26218_ (.B1(_04635_),
    .Y(_01122_),
    .A1(net7534),
    .A2(net8108));
 sg13g2_nand2_1 _26219_ (.Y(_04636_),
    .A(net3042),
    .B(net8109));
 sg13g2_o21ai_1 _26220_ (.B1(_04636_),
    .Y(_01123_),
    .A1(net7533),
    .A2(net8109));
 sg13g2_nand2_1 _26221_ (.Y(_04637_),
    .A(net3997),
    .B(net8110));
 sg13g2_o21ai_1 _26222_ (.B1(_04637_),
    .Y(_01124_),
    .A1(net7519),
    .A2(net8110));
 sg13g2_nand2_1 _26223_ (.Y(_04638_),
    .A(net3399),
    .B(net8117));
 sg13g2_o21ai_1 _26224_ (.B1(_04638_),
    .Y(_01125_),
    .A1(net7507),
    .A2(net8117));
 sg13g2_nand2_1 _26225_ (.Y(_04639_),
    .A(net3553),
    .B(net8112));
 sg13g2_o21ai_1 _26226_ (.B1(_04639_),
    .Y(_01126_),
    .A1(net7513),
    .A2(net8112));
 sg13g2_nand2_1 _26227_ (.Y(_04640_),
    .A(net3076),
    .B(net8115));
 sg13g2_o21ai_1 _26228_ (.B1(_04640_),
    .Y(_01127_),
    .A1(net7495),
    .A2(net8115));
 sg13g2_nand2_1 _26229_ (.Y(_04641_),
    .A(net3251),
    .B(net8109));
 sg13g2_o21ai_1 _26230_ (.B1(_04641_),
    .Y(_01128_),
    .A1(net7499),
    .A2(net8109));
 sg13g2_nand2_1 _26231_ (.Y(_04642_),
    .A(net3339),
    .B(net8112));
 sg13g2_o21ai_1 _26232_ (.B1(_04642_),
    .Y(_01129_),
    .A1(net7645),
    .A2(net8112));
 sg13g2_nand2_1 _26233_ (.Y(_04643_),
    .A(net2998),
    .B(net8112));
 sg13g2_o21ai_1 _26234_ (.B1(_04643_),
    .Y(_01130_),
    .A1(net7648),
    .A2(net8113));
 sg13g2_nand2_1 _26235_ (.Y(_04644_),
    .A(net3597),
    .B(net8114));
 sg13g2_o21ai_1 _26236_ (.B1(_04644_),
    .Y(_01131_),
    .A1(net7654),
    .A2(net8114));
 sg13g2_nand2_1 _26237_ (.Y(_04645_),
    .A(net3726),
    .B(net8111));
 sg13g2_o21ai_1 _26238_ (.B1(_04645_),
    .Y(_01132_),
    .A1(net7660),
    .A2(net8111));
 sg13g2_nand2_1 _26239_ (.Y(_04646_),
    .A(net3828),
    .B(net8111));
 sg13g2_o21ai_1 _26240_ (.B1(_04646_),
    .Y(_01133_),
    .A1(net7640),
    .A2(net8111));
 sg13g2_nand2_1 _26241_ (.Y(_04647_),
    .A(net3041),
    .B(net8113));
 sg13g2_o21ai_1 _26242_ (.B1(_04647_),
    .Y(_01134_),
    .A1(net7625),
    .A2(net8113));
 sg13g2_nand2_1 _26243_ (.Y(_04648_),
    .A(net3416),
    .B(_04617_));
 sg13g2_o21ai_1 _26244_ (.B1(_04648_),
    .Y(_01135_),
    .A1(net7622),
    .A2(net8111));
 sg13g2_nand2_1 _26245_ (.Y(_04649_),
    .A(net3546),
    .B(net8110));
 sg13g2_o21ai_1 _26246_ (.B1(_04649_),
    .Y(_01136_),
    .A1(net7633),
    .A2(net8110));
 sg13g2_nor2_1 _26247_ (.A(_10596_),
    .B(_13283_),
    .Y(_04650_));
 sg13g2_o21ai_1 _26248_ (.B1(_10846_),
    .Y(_04651_),
    .A1(_10596_),
    .A2(_13283_));
 sg13g2_and4_1 _26249_ (.A(net9202),
    .B(net9203),
    .C(net8980),
    .D(net8974),
    .X(_04652_));
 sg13g2_nand2_1 _26250_ (.Y(_04653_),
    .A(net8977),
    .B(_03811_));
 sg13g2_o21ai_1 _26251_ (.B1(_10883_),
    .Y(_04654_),
    .A1(net9200),
    .A2(_10847_));
 sg13g2_o21ai_1 _26252_ (.B1(_11738_),
    .Y(_04655_),
    .A1(net9202),
    .A2(_10979_));
 sg13g2_a221oi_1 _26253_ (.B2(_04653_),
    .C1(_04652_),
    .B1(_04655_),
    .A1(_03810_),
    .Y(_04656_),
    .A2(_04654_));
 sg13g2_nand2b_1 _26254_ (.Y(_04657_),
    .B(_04656_),
    .A_N(_12465_));
 sg13g2_nor2_2 _26255_ (.A(_10876_),
    .B(_04657_),
    .Y(_04658_));
 sg13g2_and2_1 _26256_ (.A(_04651_),
    .B(_04658_),
    .X(_04659_));
 sg13g2_o21ai_1 _26257_ (.B1(net9381),
    .Y(_04660_),
    .A1(net2680),
    .A2(_04659_));
 sg13g2_a21oi_1 _26258_ (.A1(_10553_),
    .A2(_04659_),
    .Y(_01137_),
    .B1(_04660_));
 sg13g2_a21oi_2 _26259_ (.B1(_10553_),
    .Y(_04661_),
    .A2(_04658_),
    .A1(_04651_));
 sg13g2_nand2_1 _26260_ (.Y(_04662_),
    .A(net5071),
    .B(_04661_));
 sg13g2_o21ai_1 _26261_ (.B1(net9372),
    .Y(_04663_),
    .A1(net5071),
    .A2(_04661_));
 sg13g2_nor2b_1 _26262_ (.A(net5072),
    .B_N(_04662_),
    .Y(_01138_));
 sg13g2_and2_1 _26263_ (.A(net4129),
    .B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[1] ),
    .X(_04664_));
 sg13g2_nand2_1 _26264_ (.Y(_04665_),
    .A(_04661_),
    .B(_04664_));
 sg13g2_a221oi_1 _26265_ (.B2(_04661_),
    .C1(net9036),
    .B1(_04664_),
    .A1(_10552_),
    .Y(_01139_),
    .A2(_04662_));
 sg13g2_nor2_1 _26266_ (.A(_10551_),
    .B(_04665_),
    .Y(_04666_));
 sg13g2_a21oi_1 _26267_ (.A1(_10551_),
    .A2(_04665_),
    .Y(_04667_),
    .B1(net9036));
 sg13g2_nor2b_1 _26268_ (.A(_04666_),
    .B_N(_04667_),
    .Y(_01140_));
 sg13g2_nand4_1 _26269_ (.B(net5366),
    .C(_04661_),
    .A(net4903),
    .Y(_04668_),
    .D(_04664_));
 sg13g2_o21ai_1 _26270_ (.B1(net9371),
    .Y(_04669_),
    .A1(net4903),
    .A2(_04666_));
 sg13g2_nor2b_1 _26271_ (.A(net4904),
    .B_N(_04668_),
    .Y(_01141_));
 sg13g2_xnor2_1 _26272_ (.Y(_04670_),
    .A(_10550_),
    .B(_04668_));
 sg13g2_nor2_1 _26273_ (.A(net9035),
    .B(_04670_),
    .Y(_01142_));
 sg13g2_o21ai_1 _26274_ (.B1(_10549_),
    .Y(_04671_),
    .A1(_10550_),
    .A2(_04668_));
 sg13g2_inv_1 _26275_ (.Y(_04672_),
    .A(net5496));
 sg13g2_nor3_1 _26276_ (.A(_10549_),
    .B(_10550_),
    .C(_04668_),
    .Y(_04673_));
 sg13g2_nor3_1 _26277_ (.A(net9035),
    .B(_04672_),
    .C(_04673_),
    .Y(_01143_));
 sg13g2_nor4_2 _26278_ (.A(_10548_),
    .B(_10549_),
    .C(_10550_),
    .Y(_04674_),
    .D(_04668_));
 sg13g2_o21ai_1 _26279_ (.B1(net9370),
    .Y(_04675_),
    .A1(net4920),
    .A2(_04673_));
 sg13g2_nor2_1 _26280_ (.A(_04674_),
    .B(_04675_),
    .Y(_01144_));
 sg13g2_xnor2_1 _26281_ (.Y(_04676_),
    .A(net5006),
    .B(_04674_));
 sg13g2_nor2_1 _26282_ (.A(net9023),
    .B(net5007),
    .Y(_01145_));
 sg13g2_a21oi_1 _26283_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[8] ),
    .A2(_04674_),
    .Y(_04677_),
    .B1(net4114));
 sg13g2_nand3_1 _26284_ (.B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[8] ),
    .C(_04674_),
    .A(net4114),
    .Y(_04678_));
 sg13g2_nand2_1 _26285_ (.Y(_04679_),
    .A(net9348),
    .B(_04678_));
 sg13g2_nor2_1 _26286_ (.A(net4115),
    .B(_04679_),
    .Y(_01146_));
 sg13g2_nand4_1 _26287_ (.B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[9] ),
    .C(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[8] ),
    .A(net3098),
    .Y(_04680_),
    .D(_04674_));
 sg13g2_nand2_1 _26288_ (.Y(_04681_),
    .A(net9346),
    .B(_04680_));
 sg13g2_a21oi_1 _26289_ (.A1(_10547_),
    .A2(_04678_),
    .Y(_01147_),
    .B1(_04681_));
 sg13g2_and2_1 _26290_ (.A(_10546_),
    .B(_04680_),
    .X(_04682_));
 sg13g2_nor2_1 _26291_ (.A(_10546_),
    .B(_04680_),
    .Y(_04683_));
 sg13g2_nor3_1 _26292_ (.A(net9022),
    .B(_04682_),
    .C(_04683_),
    .Y(_01148_));
 sg13g2_xnor2_1 _26293_ (.Y(_04684_),
    .A(net4697),
    .B(_04683_));
 sg13g2_nor2_1 _26294_ (.A(net9029),
    .B(net4698),
    .Y(_01149_));
 sg13g2_a21oi_1 _26295_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[12] ),
    .A2(_04683_),
    .Y(_04685_),
    .B1(net4483));
 sg13g2_nor4_2 _26296_ (.A(_10544_),
    .B(_10545_),
    .C(_10546_),
    .Y(_04686_),
    .D(_04680_));
 sg13g2_nor3_1 _26297_ (.A(net9029),
    .B(net4484),
    .C(_04686_),
    .Y(_01150_));
 sg13g2_o21ai_1 _26298_ (.B1(net9357),
    .Y(_04687_),
    .A1(net5278),
    .A2(_04686_));
 sg13g2_a21oi_1 _26299_ (.A1(net5278),
    .A2(_04686_),
    .Y(_01151_),
    .B1(_04687_));
 sg13g2_a21oi_1 _26300_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[14] ),
    .A2(_04686_),
    .Y(_04688_),
    .B1(net4387));
 sg13g2_and3_2 _26301_ (.X(_04689_),
    .A(net4387),
    .B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[14] ),
    .C(_04686_));
 sg13g2_nor3_1 _26302_ (.A(net9017),
    .B(net4388),
    .C(_04689_),
    .Y(_01152_));
 sg13g2_xnor2_1 _26303_ (.Y(_04690_),
    .A(net5438),
    .B(_04689_));
 sg13g2_nor2_1 _26304_ (.A(net9018),
    .B(_04690_),
    .Y(_01153_));
 sg13g2_a21oi_1 _26305_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[16] ),
    .A2(_04689_),
    .Y(_04691_),
    .B1(net4935));
 sg13g2_and3_1 _26306_ (.X(_04692_),
    .A(net4935),
    .B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[16] ),
    .C(_04689_));
 sg13g2_nor3_1 _26307_ (.A(net9018),
    .B(net4936),
    .C(_04692_),
    .Y(_01154_));
 sg13g2_nand3_1 _26308_ (.B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[17] ),
    .C(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[16] ),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[18] ),
    .Y(_04693_));
 sg13g2_nand2_1 _26309_ (.Y(_04694_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[18] ),
    .B(_04692_));
 sg13g2_xnor2_1 _26310_ (.Y(_04695_),
    .A(net5433),
    .B(_04692_));
 sg13g2_nor2_1 _26311_ (.A(net9016),
    .B(_04695_),
    .Y(_01155_));
 sg13g2_nand3_1 _26312_ (.B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[18] ),
    .C(_04692_),
    .A(net5387),
    .Y(_04696_));
 sg13g2_xor2_1 _26313_ (.B(_04694_),
    .A(net5387),
    .X(_04697_));
 sg13g2_nor2_1 _26314_ (.A(net9016),
    .B(net5388),
    .Y(_01156_));
 sg13g2_nor2_1 _26315_ (.A(_10543_),
    .B(_04696_),
    .Y(_04698_));
 sg13g2_xnor2_1 _26316_ (.Y(_04699_),
    .A(_10543_),
    .B(_04696_));
 sg13g2_nor2_1 _26317_ (.A(net9018),
    .B(net5525),
    .Y(_01157_));
 sg13g2_nand2_1 _26318_ (.Y(_04700_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[21] ),
    .B(_04698_));
 sg13g2_xnor2_1 _26319_ (.Y(_04701_),
    .A(net5299),
    .B(_04698_));
 sg13g2_nor2_1 _26320_ (.A(net9018),
    .B(_04701_),
    .Y(_01158_));
 sg13g2_nand4_1 _26321_ (.B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[21] ),
    .C(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[20] ),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[22] ),
    .Y(_04702_),
    .D(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[19] ));
 sg13g2_nand3_1 _26322_ (.B(net5299),
    .C(_04698_),
    .A(net5159),
    .Y(_04703_));
 sg13g2_xor2_1 _26323_ (.B(_04700_),
    .A(net5159),
    .X(_04704_));
 sg13g2_nor2_1 _26324_ (.A(net9018),
    .B(net5160),
    .Y(_01159_));
 sg13g2_nor2_1 _26325_ (.A(_10542_),
    .B(_04703_),
    .Y(_04705_));
 sg13g2_xnor2_1 _26326_ (.Y(_04706_),
    .A(_10542_),
    .B(_04703_));
 sg13g2_nor2_1 _26327_ (.A(net9019),
    .B(_04706_),
    .Y(_01160_));
 sg13g2_xnor2_1 _26328_ (.Y(_04707_),
    .A(net5529),
    .B(_04705_));
 sg13g2_nor2_1 _26329_ (.A(net9018),
    .B(_04707_),
    .Y(_01161_));
 sg13g2_a21o_1 _26330_ (.A2(_04705_),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[24] ),
    .B1(net5558),
    .X(_04708_));
 sg13g2_nand3_1 _26331_ (.B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[24] ),
    .C(_04705_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[25] ),
    .Y(_04709_));
 sg13g2_and3_1 _26332_ (.X(_01162_),
    .A(net9344),
    .B(_04708_),
    .C(_04709_));
 sg13g2_nor2b_1 _26333_ (.A(net5415),
    .B_N(_04709_),
    .Y(_04710_));
 sg13g2_nand3_1 _26334_ (.B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[21] ),
    .C(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[16] ),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[22] ),
    .Y(_04711_));
 sg13g2_nand4_1 _26335_ (.B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[23] ),
    .C(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[18] ),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[26] ),
    .Y(_04712_),
    .D(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[17] ));
 sg13g2_nand4_1 _26336_ (.B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[24] ),
    .C(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[20] ),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[25] ),
    .Y(_04713_),
    .D(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[19] ));
 sg13g2_nor3_1 _26337_ (.A(_04711_),
    .B(_04712_),
    .C(_04713_),
    .Y(_04714_));
 sg13g2_nand4_1 _26338_ (.B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[14] ),
    .C(_04686_),
    .A(net4387),
    .Y(_04715_),
    .D(_04714_));
 sg13g2_nand4_1 _26339_ (.B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[25] ),
    .C(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[24] ),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[26] ),
    .Y(_04716_),
    .D(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[23] ));
 sg13g2_nor3_1 _26340_ (.A(_04693_),
    .B(_04702_),
    .C(_04716_),
    .Y(_04717_));
 sg13g2_and4_1 _26341_ (.A(net4387),
    .B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[14] ),
    .C(_04686_),
    .D(_04717_),
    .X(_04718_));
 sg13g2_nor3_1 _26342_ (.A(net9017),
    .B(_04710_),
    .C(_04718_),
    .Y(_01163_));
 sg13g2_o21ai_1 _26343_ (.B1(net9357),
    .Y(_04719_),
    .A1(net5486),
    .A2(_04718_));
 sg13g2_and2_1 _26344_ (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[27] ),
    .B(_04718_),
    .X(_04720_));
 sg13g2_nor2_1 _26345_ (.A(_04719_),
    .B(_04720_),
    .Y(_01164_));
 sg13g2_nor2_1 _26346_ (.A(net5238),
    .B(_04720_),
    .Y(_04721_));
 sg13g2_a21oi_1 _26347_ (.A1(net5238),
    .A2(_04720_),
    .Y(_04722_),
    .B1(net9027));
 sg13g2_nor2b_1 _26348_ (.A(_04721_),
    .B_N(_04722_),
    .Y(_01165_));
 sg13g2_a21oi_1 _26349_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[28] ),
    .A2(_04720_),
    .Y(_04723_),
    .B1(net4474));
 sg13g2_and2_1 _26350_ (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[29] ),
    .B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[28] ),
    .X(_04724_));
 sg13g2_nand2_1 _26351_ (.Y(_04725_),
    .A(net4474),
    .B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[28] ));
 sg13g2_and2_1 _26352_ (.A(_04720_),
    .B(_04724_),
    .X(_04726_));
 sg13g2_nor3_1 _26353_ (.A(net9027),
    .B(net4475),
    .C(_04726_),
    .Y(_01166_));
 sg13g2_nor2_1 _26354_ (.A(net5219),
    .B(_04726_),
    .Y(_04727_));
 sg13g2_nor4_2 _26355_ (.A(_10540_),
    .B(_10541_),
    .C(_04715_),
    .Y(_04728_),
    .D(_04725_));
 sg13g2_nand4_1 _26356_ (.B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[27] ),
    .C(_04718_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[30] ),
    .Y(_04729_),
    .D(_04724_));
 sg13g2_nor3_1 _26357_ (.A(net9027),
    .B(_04727_),
    .C(_04728_),
    .Y(_01167_));
 sg13g2_nor2_2 _26358_ (.A(_10539_),
    .B(_04729_),
    .Y(_04730_));
 sg13g2_o21ai_1 _26359_ (.B1(net9355),
    .Y(_04731_),
    .A1(net5411),
    .A2(_04728_));
 sg13g2_nor2_1 _26360_ (.A(_04730_),
    .B(net5412),
    .Y(_01168_));
 sg13g2_nor2_1 _26361_ (.A(net5449),
    .B(_04730_),
    .Y(_04732_));
 sg13g2_nand2_1 _26362_ (.Y(_04733_),
    .A(net5449),
    .B(_04730_));
 sg13g2_nand2_1 _26363_ (.Y(_04734_),
    .A(net9355),
    .B(_04733_));
 sg13g2_nor2_1 _26364_ (.A(_04732_),
    .B(_04734_),
    .Y(_01169_));
 sg13g2_nand2b_1 _26365_ (.Y(_04735_),
    .B(_04733_),
    .A_N(net5555));
 sg13g2_nand3_1 _26366_ (.B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[32] ),
    .C(_04730_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[33] ),
    .Y(_04736_));
 sg13g2_and3_1 _26367_ (.X(_01170_),
    .A(net9355),
    .B(_04735_),
    .C(_04736_));
 sg13g2_and2_1 _26368_ (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[34] ),
    .B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[33] ),
    .X(_04737_));
 sg13g2_nand2_1 _26369_ (.Y(_04738_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[34] ),
    .B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[33] ));
 sg13g2_nand4_1 _26370_ (.B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[31] ),
    .C(_04728_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[32] ),
    .Y(_04739_),
    .D(_04737_));
 sg13g2_nand2_1 _26371_ (.Y(_04740_),
    .A(net9355),
    .B(_04739_));
 sg13g2_nor4_2 _26372_ (.A(_10538_),
    .B(_10539_),
    .C(_04729_),
    .Y(_04741_),
    .D(_04738_));
 sg13g2_a21oi_1 _26373_ (.A1(_10537_),
    .A2(_04736_),
    .Y(_01171_),
    .B1(_04740_));
 sg13g2_nor2_1 _26374_ (.A(net5314),
    .B(_04741_),
    .Y(_04742_));
 sg13g2_and2_1 _26375_ (.A(net5314),
    .B(_04741_),
    .X(_04743_));
 sg13g2_nor3_1 _26376_ (.A(net9022),
    .B(_04742_),
    .C(_04743_),
    .Y(_01172_));
 sg13g2_o21ai_1 _26377_ (.B1(net9347),
    .Y(_04744_),
    .A1(net5430),
    .A2(_04743_));
 sg13g2_a21oi_1 _26378_ (.A1(net5430),
    .A2(_04743_),
    .Y(_01173_),
    .B1(_04744_));
 sg13g2_a21oi_1 _26379_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[36] ),
    .A2(_04743_),
    .Y(_04745_),
    .B1(net5199));
 sg13g2_nor4_2 _26380_ (.A(_10534_),
    .B(_10535_),
    .C(_10536_),
    .Y(_04746_),
    .D(_04739_));
 sg13g2_and4_1 _26381_ (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[37] ),
    .B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[36] ),
    .C(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[35] ),
    .D(_04741_),
    .X(_04747_));
 sg13g2_nor3_1 _26382_ (.A(net9022),
    .B(net5200),
    .C(_04747_),
    .Y(_01174_));
 sg13g2_nor2_1 _26383_ (.A(net5424),
    .B(_04746_),
    .Y(_04748_));
 sg13g2_and2_1 _26384_ (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[38] ),
    .B(_04747_),
    .X(_04749_));
 sg13g2_nor3_1 _26385_ (.A(net9026),
    .B(_04748_),
    .C(_04749_),
    .Y(_01175_));
 sg13g2_o21ai_1 _26386_ (.B1(net9346),
    .Y(_04750_),
    .A1(net4755),
    .A2(_04749_));
 sg13g2_a21oi_1 _26387_ (.A1(net4755),
    .A2(_04749_),
    .Y(_01176_),
    .B1(_04750_));
 sg13g2_a21oi_1 _26388_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[39] ),
    .A2(_04749_),
    .Y(_04751_),
    .B1(net4439));
 sg13g2_nand4_1 _26389_ (.B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[39] ),
    .C(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[38] ),
    .A(net4439),
    .Y(_04752_),
    .D(_04746_));
 sg13g2_nand4_1 _26390_ (.B(net4755),
    .C(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[38] ),
    .A(net4439),
    .Y(_04753_),
    .D(_04747_));
 sg13g2_nand2_1 _26391_ (.Y(_04754_),
    .A(net9346),
    .B(_04752_));
 sg13g2_nor2_1 _26392_ (.A(net4440),
    .B(_04754_),
    .Y(_01177_));
 sg13g2_nor2_1 _26393_ (.A(_10533_),
    .B(_04753_),
    .Y(_04755_));
 sg13g2_a21oi_1 _26394_ (.A1(_10533_),
    .A2(_04753_),
    .Y(_04756_),
    .B1(net9026));
 sg13g2_nor2b_1 _26395_ (.A(_04755_),
    .B_N(_04756_),
    .Y(_01178_));
 sg13g2_o21ai_1 _26396_ (.B1(_10532_),
    .Y(_04757_),
    .A1(_10533_),
    .A2(_04752_));
 sg13g2_nand2_1 _26397_ (.Y(_04758_),
    .A(net5344),
    .B(_04755_));
 sg13g2_and3_1 _26398_ (.X(_01179_),
    .A(net9347),
    .B(_04757_),
    .C(_04758_));
 sg13g2_a21oi_1 _26399_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[42] ),
    .A2(_04755_),
    .Y(_04759_),
    .B1(net4058));
 sg13g2_nor4_2 _26400_ (.A(_10531_),
    .B(_10532_),
    .C(_10533_),
    .Y(_04760_),
    .D(_04752_));
 sg13g2_nor4_2 _26401_ (.A(_10531_),
    .B(_10532_),
    .C(_10533_),
    .Y(_04761_),
    .D(_04753_));
 sg13g2_nor3_1 _26402_ (.A(net9022),
    .B(net4059),
    .C(_04760_),
    .Y(_01180_));
 sg13g2_and2_1 _26403_ (.A(net5274),
    .B(_04761_),
    .X(_04762_));
 sg13g2_o21ai_1 _26404_ (.B1(net9354),
    .Y(_04763_),
    .A1(net5274),
    .A2(_04761_));
 sg13g2_nor2_1 _26405_ (.A(_04762_),
    .B(net5275),
    .Y(_01181_));
 sg13g2_and2_1 _26406_ (.A(net5179),
    .B(_04762_),
    .X(_04764_));
 sg13g2_o21ai_1 _26407_ (.B1(net9354),
    .Y(_04765_),
    .A1(net5179),
    .A2(_04762_));
 sg13g2_nor2_1 _26408_ (.A(_04764_),
    .B(_04765_),
    .Y(_01182_));
 sg13g2_or2_1 _26409_ (.X(_04766_),
    .B(_04764_),
    .A(net5506));
 sg13g2_nand4_1 _26410_ (.B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[45] ),
    .C(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[44] ),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[46] ),
    .Y(_04767_),
    .D(_04760_));
 sg13g2_nand4_1 _26411_ (.B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[45] ),
    .C(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[44] ),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[46] ),
    .Y(_04768_),
    .D(_04761_));
 sg13g2_and3_1 _26412_ (.X(_01183_),
    .A(net9354),
    .B(_04766_),
    .C(_04768_));
 sg13g2_nand2b_1 _26413_ (.Y(_04769_),
    .B(_04767_),
    .A_N(net5479));
 sg13g2_nand3_1 _26414_ (.B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[46] ),
    .C(_04764_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[47] ),
    .Y(_04770_));
 sg13g2_and3_1 _26415_ (.X(_01184_),
    .A(net9358),
    .B(_04769_),
    .C(_04770_));
 sg13g2_nand2_2 _26416_ (.Y(_04771_),
    .A(net3791),
    .B(net5479));
 sg13g2_o21ai_1 _26417_ (.B1(net9359),
    .Y(_04772_),
    .A1(_04767_),
    .A2(_04771_));
 sg13g2_a21oi_1 _26418_ (.A1(_10530_),
    .A2(_04770_),
    .Y(_01185_),
    .B1(_04772_));
 sg13g2_o21ai_1 _26419_ (.B1(_10529_),
    .Y(_04773_),
    .A1(_04767_),
    .A2(_04771_));
 sg13g2_or3_1 _26420_ (.A(_10529_),
    .B(_04768_),
    .C(_04771_),
    .X(_04774_));
 sg13g2_and3_1 _26421_ (.X(_01186_),
    .A(net9360),
    .B(_04773_),
    .C(_04774_));
 sg13g2_nor4_2 _26422_ (.A(_10528_),
    .B(_10529_),
    .C(_04767_),
    .Y(_04775_),
    .D(_04771_));
 sg13g2_nor4_2 _26423_ (.A(_10528_),
    .B(_10529_),
    .C(_04768_),
    .Y(_04776_),
    .D(_04771_));
 sg13g2_a21o_1 _26424_ (.A2(_04774_),
    .A1(_10528_),
    .B1(net9027),
    .X(_04777_));
 sg13g2_nor2_1 _26425_ (.A(_04776_),
    .B(_04777_),
    .Y(_01187_));
 sg13g2_or2_1 _26426_ (.X(_04778_),
    .B(_04775_),
    .A(net5507));
 sg13g2_nand2_1 _26427_ (.Y(_04779_),
    .A(net5507),
    .B(_04776_));
 sg13g2_and3_1 _26428_ (.X(_01188_),
    .A(net9360),
    .B(_04778_),
    .C(_04779_));
 sg13g2_o21ai_1 _26429_ (.B1(net9360),
    .Y(_04780_),
    .A1(_10527_),
    .A2(_04779_));
 sg13g2_a21oi_1 _26430_ (.A1(_10527_),
    .A2(_04779_),
    .Y(_01189_),
    .B1(_04780_));
 sg13g2_o21ai_1 _26431_ (.B1(_10526_),
    .Y(_04781_),
    .A1(_10527_),
    .A2(_04779_));
 sg13g2_and4_1 _26432_ (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[53] ),
    .B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[52] ),
    .C(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[51] ),
    .D(_04775_),
    .X(_04782_));
 sg13g2_nand4_1 _26433_ (.B(net5093),
    .C(net5507),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[53] ),
    .Y(_04783_),
    .D(_04775_));
 sg13g2_nand4_1 _26434_ (.B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[52] ),
    .C(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[51] ),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[53] ),
    .Y(_04784_),
    .D(_04776_));
 sg13g2_and3_1 _26435_ (.X(_01190_),
    .A(net9359),
    .B(_04781_),
    .C(_04783_));
 sg13g2_nor2_1 _26436_ (.A(net4647),
    .B(_04782_),
    .Y(_04785_));
 sg13g2_nor2_1 _26437_ (.A(_10525_),
    .B(_04783_),
    .Y(_04786_));
 sg13g2_nor3_1 _26438_ (.A(net9033),
    .B(net4648),
    .C(_04786_),
    .Y(_01191_));
 sg13g2_nor2_1 _26439_ (.A(net5075),
    .B(_04786_),
    .Y(_04787_));
 sg13g2_nand2_1 _26440_ (.Y(_04788_),
    .A(net5075),
    .B(_04786_));
 sg13g2_nand2_1 _26441_ (.Y(_04789_),
    .A(net9365),
    .B(_04788_));
 sg13g2_nor2_1 _26442_ (.A(net5076),
    .B(_04789_),
    .Y(_01192_));
 sg13g2_nand4_1 _26443_ (.B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[55] ),
    .C(net4647),
    .A(net4511),
    .Y(_04790_),
    .D(_04782_));
 sg13g2_nor4_1 _26444_ (.A(_10523_),
    .B(_10524_),
    .C(_10525_),
    .D(_04784_),
    .Y(_04791_));
 sg13g2_nand2_1 _26445_ (.Y(_04792_),
    .A(net9359),
    .B(_04790_));
 sg13g2_a21oi_1 _26446_ (.A1(_10523_),
    .A2(_04788_),
    .Y(_01193_),
    .B1(_04792_));
 sg13g2_nor2_1 _26447_ (.A(net5034),
    .B(_04791_),
    .Y(_04793_));
 sg13g2_nor2_2 _26448_ (.A(_10522_),
    .B(_04790_),
    .Y(_04794_));
 sg13g2_nor3_1 _26449_ (.A(net9030),
    .B(net5035),
    .C(_04794_),
    .Y(_01194_));
 sg13g2_nor2_1 _26450_ (.A(net5073),
    .B(_04794_),
    .Y(_04795_));
 sg13g2_a21oi_1 _26451_ (.A1(net5073),
    .A2(_04794_),
    .Y(_04796_),
    .B1(net9030));
 sg13g2_nor2b_1 _26452_ (.A(_04795_),
    .B_N(_04796_),
    .Y(_01195_));
 sg13g2_a21oi_1 _26453_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[58] ),
    .A2(_04794_),
    .Y(_04797_),
    .B1(net4958));
 sg13g2_nand3_1 _26454_ (.B(net5073),
    .C(_04794_),
    .A(net4958),
    .Y(_04798_));
 sg13g2_and4_1 _26455_ (.A(net4958),
    .B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[58] ),
    .C(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[57] ),
    .D(_04791_),
    .X(_04799_));
 sg13g2_nor3_1 _26456_ (.A(net9032),
    .B(net4959),
    .C(_04799_),
    .Y(_01196_));
 sg13g2_o21ai_1 _26457_ (.B1(net9365),
    .Y(_04800_),
    .A1(_10521_),
    .A2(_04798_));
 sg13g2_a21oi_1 _26458_ (.A1(_10521_),
    .A2(_04798_),
    .Y(_01197_),
    .B1(_04800_));
 sg13g2_o21ai_1 _26459_ (.B1(_10520_),
    .Y(_04801_),
    .A1(_10521_),
    .A2(_04798_));
 sg13g2_or3_1 _26460_ (.A(_10520_),
    .B(_10521_),
    .C(_04798_),
    .X(_04802_));
 sg13g2_and3_1 _26461_ (.X(_01198_),
    .A(net9367),
    .B(_04801_),
    .C(_04802_));
 sg13g2_nand4_1 _26462_ (.B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[61] ),
    .C(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[60] ),
    .A(net3193),
    .Y(_04803_),
    .D(_04799_));
 sg13g2_nand2_1 _26463_ (.Y(_04804_),
    .A(net9367),
    .B(_04803_));
 sg13g2_a21oi_1 _26464_ (.A1(_10519_),
    .A2(_04802_),
    .Y(_01199_),
    .B1(_04804_));
 sg13g2_o21ai_1 _26465_ (.B1(net9367),
    .Y(_04805_),
    .A1(_10518_),
    .A2(_04803_));
 sg13g2_a21oi_1 _26466_ (.A1(_10518_),
    .A2(_04803_),
    .Y(_01200_),
    .B1(_04805_));
 sg13g2_nor2_2 _26467_ (.A(net9706),
    .B(_13832_),
    .Y(_04806_));
 sg13g2_or2_2 _26468_ (.X(_04807_),
    .B(_13832_),
    .A(net9706));
 sg13g2_nand2_2 _26469_ (.Y(_04808_),
    .A(_11651_),
    .B(net8254));
 sg13g2_or2_2 _26470_ (.X(_04809_),
    .B(_04808_),
    .A(_11109_));
 sg13g2_nor2_2 _26471_ (.A(_11100_),
    .B(_04809_),
    .Y(_04810_));
 sg13g2_nor3_2 _26472_ (.A(_11090_),
    .B(_11100_),
    .C(_04809_),
    .Y(_04811_));
 sg13g2_nor2b_2 _26473_ (.A(_11212_),
    .B_N(_04811_),
    .Y(_04812_));
 sg13g2_nand2b_1 _26474_ (.Y(_04813_),
    .B(_04812_),
    .A_N(_11250_));
 sg13g2_or2_2 _26475_ (.X(_04814_),
    .B(_04813_),
    .A(_11225_));
 sg13g2_or2_2 _26476_ (.X(_04815_),
    .B(_04814_),
    .A(_11238_));
 sg13g2_nor2_2 _26477_ (.A(_11294_),
    .B(_04815_),
    .Y(_04816_));
 sg13g2_nand2_2 _26478_ (.Y(_04817_),
    .A(_11307_),
    .B(_04816_));
 sg13g2_nand3_1 _26479_ (.B(net8290),
    .C(_04816_),
    .A(_11273_),
    .Y(_04818_));
 sg13g2_or2_1 _26480_ (.X(_04819_),
    .B(_04818_),
    .A(_11282_));
 sg13g2_nand2b_1 _26481_ (.Y(_04820_),
    .B(_11383_),
    .A_N(_04819_));
 sg13g2_nand2b_1 _26482_ (.Y(_04821_),
    .B(_11416_),
    .A_N(_04820_));
 sg13g2_nor2_1 _26483_ (.A(_11394_),
    .B(_04821_),
    .Y(_04822_));
 sg13g2_nand2b_1 _26484_ (.Y(_04823_),
    .B(_04822_),
    .A_N(_11404_));
 sg13g2_nand2b_1 _26485_ (.Y(_04824_),
    .B(_11354_),
    .A_N(_04823_));
 sg13g2_nand2b_1 _26486_ (.Y(_04825_),
    .B(_11366_),
    .A_N(_04824_));
 sg13g2_nand2b_1 _26487_ (.Y(_04826_),
    .B(_11326_),
    .A_N(_04825_));
 sg13g2_nand2b_1 _26488_ (.Y(_04827_),
    .B(_11339_),
    .A_N(_04826_));
 sg13g2_nor2_1 _26489_ (.A(_11465_),
    .B(_04827_),
    .Y(_04828_));
 sg13g2_nand2_1 _26490_ (.Y(_04829_),
    .A(_11477_),
    .B(_04828_));
 sg13g2_or2_1 _26491_ (.X(_04830_),
    .B(_04829_),
    .A(_11442_));
 sg13g2_nand2b_1 _26492_ (.Y(_04831_),
    .B(_11453_),
    .A_N(_04830_));
 sg13g2_nand2b_1 _26493_ (.Y(_04832_),
    .B(_11495_),
    .A_N(_04831_));
 sg13g2_or2_1 _26494_ (.X(_04833_),
    .B(_04832_),
    .A(_11080_));
 sg13g2_nor2_2 _26495_ (.A(net8008),
    .B(_04833_),
    .Y(_04834_));
 sg13g2_o21ai_1 _26496_ (.B1(_11021_),
    .Y(_04835_),
    .A1(_04807_),
    .A2(_04834_));
 sg13g2_and3_2 _26497_ (.X(_04836_),
    .A(_11016_),
    .B(_11020_),
    .C(_04806_));
 sg13g2_nand3_1 _26498_ (.B(_11020_),
    .C(_04806_),
    .A(_11016_),
    .Y(_04837_));
 sg13g2_xnor2_1 _26499_ (.Y(_04838_),
    .A(net8007),
    .B(_04832_));
 sg13g2_nor2_1 _26500_ (.A(net8482),
    .B(_04838_),
    .Y(_04839_));
 sg13g2_a21oi_2 _26501_ (.B1(_04839_),
    .Y(_04840_),
    .A2(net8482),
    .A1(net8007));
 sg13g2_xnor2_1 _26502_ (.Y(_04841_),
    .A(_11453_),
    .B(_04830_));
 sg13g2_nor2_1 _26503_ (.A(_11453_),
    .B(net8485),
    .Y(_04842_));
 sg13g2_a21oi_2 _26504_ (.B1(_04842_),
    .Y(_04843_),
    .A2(_04841_),
    .A1(net8485));
 sg13g2_xnor2_1 _26505_ (.Y(_04844_),
    .A(_11476_),
    .B(_04828_));
 sg13g2_nor2_1 _26506_ (.A(_11477_),
    .B(net8485),
    .Y(_04845_));
 sg13g2_a21oi_2 _26507_ (.B1(_04845_),
    .Y(_04846_),
    .A2(_04844_),
    .A1(net8485));
 sg13g2_xnor2_1 _26508_ (.Y(_04847_),
    .A(_11339_),
    .B(_04826_));
 sg13g2_nor2_1 _26509_ (.A(_11339_),
    .B(net8484),
    .Y(_04848_));
 sg13g2_a21oi_2 _26510_ (.B1(_04848_),
    .Y(_04849_),
    .A2(_04847_),
    .A1(net8484));
 sg13g2_xor2_1 _26511_ (.B(_04849_),
    .A(_00165_),
    .X(_04850_));
 sg13g2_xnor2_1 _26512_ (.Y(_04851_),
    .A(_11326_),
    .B(_04825_));
 sg13g2_nor2_1 _26513_ (.A(_11326_),
    .B(net8484),
    .Y(_04852_));
 sg13g2_a21oi_2 _26514_ (.B1(_04852_),
    .Y(_04853_),
    .A2(_04851_),
    .A1(net8483));
 sg13g2_nand2_1 _26515_ (.Y(_04854_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[21] ),
    .B(_04853_));
 sg13g2_xnor2_1 _26516_ (.Y(_04855_),
    .A(_11365_),
    .B(_04824_));
 sg13g2_nor2_1 _26517_ (.A(net8480),
    .B(_04855_),
    .Y(_04856_));
 sg13g2_a21oi_2 _26518_ (.B1(_04856_),
    .Y(_04857_),
    .A2(net8480),
    .A1(_11365_));
 sg13g2_nand2_1 _26519_ (.Y(_04858_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[20] ),
    .B(_04857_));
 sg13g2_xnor2_1 _26520_ (.Y(_04859_),
    .A(_00167_),
    .B(_04857_));
 sg13g2_xnor2_1 _26521_ (.Y(_04860_),
    .A(_11354_),
    .B(_04823_));
 sg13g2_nor2_1 _26522_ (.A(_11354_),
    .B(net8483),
    .Y(_04861_));
 sg13g2_a21oi_2 _26523_ (.B1(_04861_),
    .Y(_04862_),
    .A2(_04860_),
    .A1(net8483));
 sg13g2_xnor2_1 _26524_ (.Y(_04863_),
    .A(net8381),
    .B(_04818_));
 sg13g2_nor2_1 _26525_ (.A(net8481),
    .B(_04863_),
    .Y(_04864_));
 sg13g2_a21oi_2 _26526_ (.B1(_04864_),
    .Y(_04865_),
    .A2(net8480),
    .A1(net8381));
 sg13g2_and2_1 _26527_ (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[14] ),
    .B(_04865_),
    .X(_04866_));
 sg13g2_xor2_1 _26528_ (.B(_04810_),
    .A(net8522),
    .X(_04867_));
 sg13g2_nor2_1 _26529_ (.A(net8522),
    .B(net8483),
    .Y(_04868_));
 sg13g2_a21oi_2 _26530_ (.B1(_04868_),
    .Y(_04869_),
    .A2(_04867_),
    .A1(net8483));
 sg13g2_nand2b_1 _26531_ (.Y(_04870_),
    .B(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[6] ),
    .A_N(_04869_));
 sg13g2_nor2_1 _26532_ (.A(net8521),
    .B(net8483),
    .Y(_04871_));
 sg13g2_xnor2_1 _26533_ (.Y(_04872_),
    .A(net8521),
    .B(_04809_));
 sg13g2_a21oi_2 _26534_ (.B1(_04871_),
    .Y(_04873_),
    .A2(_04872_),
    .A1(net8483));
 sg13g2_nor2b_1 _26535_ (.A(_04873_),
    .B_N(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[5] ),
    .Y(_04874_));
 sg13g2_xnor2_1 _26536_ (.Y(_04875_),
    .A(net8520),
    .B(_04808_));
 sg13g2_nor2_1 _26537_ (.A(net8520),
    .B(net8484),
    .Y(_04876_));
 sg13g2_a21o_1 _26538_ (.A2(_04875_),
    .A1(net8484),
    .B1(_04876_),
    .X(_04877_));
 sg13g2_nand2_1 _26539_ (.Y(_04878_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[4] ),
    .B(_04877_));
 sg13g2_a21oi_1 _26540_ (.A1(net8437),
    .A2(_11651_),
    .Y(_04879_),
    .B1(net8477));
 sg13g2_xnor2_1 _26541_ (.Y(_04880_),
    .A(net8451),
    .B(_04879_));
 sg13g2_and2_1 _26542_ (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[3] ),
    .B(_04880_),
    .X(_04881_));
 sg13g2_a21oi_1 _26543_ (.A1(net8430),
    .A2(_11649_),
    .Y(_04882_),
    .B1(net8476));
 sg13g2_xnor2_1 _26544_ (.Y(_04883_),
    .A(net8441),
    .B(_04882_));
 sg13g2_nand2_1 _26545_ (.Y(_04884_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[2] ),
    .B(_04883_));
 sg13g2_a21oi_1 _26546_ (.A1(_11650_),
    .A2(net8484),
    .Y(_04885_),
    .B1(net8430));
 sg13g2_o21ai_1 _26547_ (.B1(net8424),
    .Y(_04886_),
    .A1(_11649_),
    .A2(net8476));
 sg13g2_nor3_1 _26548_ (.A(net8424),
    .B(_11649_),
    .C(net8476),
    .Y(_04887_));
 sg13g2_nand3_1 _26549_ (.B(_11650_),
    .C(net8484),
    .A(net8430),
    .Y(_04888_));
 sg13g2_nor3_1 _26550_ (.A(_10516_),
    .B(_04885_),
    .C(_04887_),
    .Y(_04889_));
 sg13g2_a221oi_1 _26551_ (.B2(_11177_),
    .C1(net8482),
    .B1(_11176_),
    .A1(_11165_),
    .Y(_04890_),
    .A2(_11166_));
 sg13g2_a221oi_1 _26552_ (.B2(_04836_),
    .C1(_11167_),
    .B1(_11180_),
    .A1(net8642),
    .Y(_04891_),
    .A2(_11163_));
 sg13g2_nor3_1 _26553_ (.A(_10517_),
    .B(_04890_),
    .C(_04891_),
    .Y(_04892_));
 sg13g2_nand2b_2 _26554_ (.Y(_04893_),
    .B(net8516),
    .A_N(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[31] ));
 sg13g2_o21ai_1 _26555_ (.B1(_10517_),
    .Y(_04894_),
    .A1(_04890_),
    .A2(_04891_));
 sg13g2_nor2b_1 _26556_ (.A(_04892_),
    .B_N(_04894_),
    .Y(_04895_));
 sg13g2_a21oi_1 _26557_ (.A1(_04893_),
    .A2(_04894_),
    .Y(_04896_),
    .B1(_04892_));
 sg13g2_nor3_1 _26558_ (.A(_00183_),
    .B(_04885_),
    .C(_04887_),
    .Y(_04897_));
 sg13g2_a21oi_1 _26559_ (.A1(_04886_),
    .A2(_04888_),
    .Y(_04898_),
    .B1(_10831_));
 sg13g2_nor3_1 _26560_ (.A(_04896_),
    .B(_04897_),
    .C(_04898_),
    .Y(_04899_));
 sg13g2_nor2_1 _26561_ (.A(_04889_),
    .B(_04899_),
    .Y(_04900_));
 sg13g2_xor2_1 _26562_ (.B(_04883_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[2] ),
    .X(_04901_));
 sg13g2_o21ai_1 _26563_ (.B1(_04901_),
    .Y(_04902_),
    .A1(_04889_),
    .A2(_04899_));
 sg13g2_xnor2_1 _26564_ (.Y(_04903_),
    .A(_10830_),
    .B(_04880_));
 sg13g2_a21oi_1 _26565_ (.A1(_04884_),
    .A2(_04902_),
    .Y(_04904_),
    .B1(_04903_));
 sg13g2_xnor2_1 _26566_ (.Y(_04905_),
    .A(_00181_),
    .B(_04877_));
 sg13g2_o21ai_1 _26567_ (.B1(_04905_),
    .Y(_04906_),
    .A1(_04881_),
    .A2(_04904_));
 sg13g2_xnor2_1 _26568_ (.Y(_04907_),
    .A(_00180_),
    .B(_04873_));
 sg13g2_a21oi_1 _26569_ (.A1(_04878_),
    .A2(_04906_),
    .Y(_04908_),
    .B1(_04907_));
 sg13g2_xnor2_1 _26570_ (.Y(_04909_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[6] ),
    .B(_04869_));
 sg13g2_o21ai_1 _26571_ (.B1(_04909_),
    .Y(_04910_),
    .A1(_04874_),
    .A2(_04908_));
 sg13g2_xor2_1 _26572_ (.B(_04811_),
    .A(net8507),
    .X(_04911_));
 sg13g2_nand2_1 _26573_ (.Y(_04912_),
    .A(net8507),
    .B(net8479));
 sg13g2_o21ai_1 _26574_ (.B1(_04912_),
    .Y(_04913_),
    .A1(net8479),
    .A2(_04911_));
 sg13g2_xnor2_1 _26575_ (.Y(_04914_),
    .A(_00179_),
    .B(_04913_));
 sg13g2_a21o_1 _26576_ (.A2(_04910_),
    .A1(_04870_),
    .B1(_04914_),
    .X(_04915_));
 sg13g2_or2_1 _26577_ (.X(_04916_),
    .B(_04913_),
    .A(_10515_));
 sg13g2_xor2_1 _26578_ (.B(_04812_),
    .A(net8505),
    .X(_04917_));
 sg13g2_nor2_1 _26579_ (.A(net8479),
    .B(_04917_),
    .Y(_04918_));
 sg13g2_a21oi_2 _26580_ (.B1(_04918_),
    .Y(_04919_),
    .A2(net8479),
    .A1(net8505));
 sg13g2_xor2_1 _26581_ (.B(_04919_),
    .A(_00178_),
    .X(_04920_));
 sg13g2_a21oi_1 _26582_ (.A1(_04915_),
    .A2(_04916_),
    .Y(_04921_),
    .B1(_04920_));
 sg13g2_a21oi_1 _26583_ (.A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[8] ),
    .A2(_04919_),
    .Y(_04922_),
    .B1(_04921_));
 sg13g2_xnor2_1 _26584_ (.Y(_04923_),
    .A(_11225_),
    .B(_04813_));
 sg13g2_nor2_1 _26585_ (.A(net8478),
    .B(_04923_),
    .Y(_04924_));
 sg13g2_a21oi_2 _26586_ (.B1(_04924_),
    .Y(_04925_),
    .A2(net8478),
    .A1(net8506));
 sg13g2_xnor2_1 _26587_ (.Y(_04926_),
    .A(_00177_),
    .B(_04925_));
 sg13g2_nand2b_1 _26588_ (.Y(_04927_),
    .B(_04926_),
    .A_N(_04922_));
 sg13g2_nand2_1 _26589_ (.Y(_04928_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[9] ),
    .B(_04925_));
 sg13g2_xnor2_1 _26590_ (.Y(_04929_),
    .A(net8382),
    .B(_04814_));
 sg13g2_nor2_1 _26591_ (.A(net8478),
    .B(_04929_),
    .Y(_04930_));
 sg13g2_a21oi_2 _26592_ (.B1(_04930_),
    .Y(_04931_),
    .A2(net8478),
    .A1(net8382));
 sg13g2_xnor2_1 _26593_ (.Y(_04932_),
    .A(_10825_),
    .B(_04931_));
 sg13g2_a21o_1 _26594_ (.A2(_04928_),
    .A1(_04927_),
    .B1(_04932_),
    .X(_04933_));
 sg13g2_nand2_1 _26595_ (.Y(_04934_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[10] ),
    .B(_04931_));
 sg13g2_xnor2_1 _26596_ (.Y(_04935_),
    .A(net8380),
    .B(_04815_));
 sg13g2_nor2_1 _26597_ (.A(net8478),
    .B(_04935_),
    .Y(_04936_));
 sg13g2_a21oi_2 _26598_ (.B1(_04936_),
    .Y(_04937_),
    .A2(net8478),
    .A1(net8380));
 sg13g2_xnor2_1 _26599_ (.Y(_04938_),
    .A(_00175_),
    .B(_04937_));
 sg13g2_inv_1 _26600_ (.Y(_04939_),
    .A(_04938_));
 sg13g2_a21oi_1 _26601_ (.A1(_04933_),
    .A2(_04934_),
    .Y(_04940_),
    .B1(_04939_));
 sg13g2_a21o_1 _26602_ (.A2(_04937_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[11] ),
    .B1(_04940_),
    .X(_04941_));
 sg13g2_xnor2_1 _26603_ (.Y(_04942_),
    .A(_11308_),
    .B(_04816_));
 sg13g2_nand2_1 _26604_ (.Y(_04943_),
    .A(net8290),
    .B(net8478));
 sg13g2_o21ai_1 _26605_ (.B1(_04943_),
    .Y(_04944_),
    .A1(net8478),
    .A2(_04942_));
 sg13g2_xnor2_1 _26606_ (.Y(_04945_),
    .A(_00174_),
    .B(_04944_));
 sg13g2_a22oi_1 _26607_ (.Y(_04946_),
    .B1(_04945_),
    .B2(_04941_),
    .A2(_04944_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[12] ));
 sg13g2_xnor2_1 _26608_ (.Y(_04947_),
    .A(_11273_),
    .B(_04817_));
 sg13g2_nand2_1 _26609_ (.Y(_04948_),
    .A(_11273_),
    .B(net8479));
 sg13g2_o21ai_1 _26610_ (.B1(_04948_),
    .Y(_04949_),
    .A1(net8480),
    .A2(_04947_));
 sg13g2_xnor2_1 _26611_ (.Y(_04950_),
    .A(_10823_),
    .B(_04949_));
 sg13g2_nand2_1 _26612_ (.Y(_04951_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[13] ),
    .B(_04949_));
 sg13g2_o21ai_1 _26613_ (.B1(_04951_),
    .Y(_04952_),
    .A1(_04946_),
    .A2(_04950_));
 sg13g2_xnor2_1 _26614_ (.Y(_04953_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[14] ),
    .B(_04865_));
 sg13g2_nor2b_1 _26615_ (.A(_04953_),
    .B_N(_04952_),
    .Y(_04954_));
 sg13g2_xnor2_1 _26616_ (.Y(_04955_),
    .A(_11383_),
    .B(_04819_));
 sg13g2_nand2_1 _26617_ (.Y(_04956_),
    .A(_11383_),
    .B(net8480));
 sg13g2_o21ai_1 _26618_ (.B1(_04956_),
    .Y(_04957_),
    .A1(net8480),
    .A2(_04955_));
 sg13g2_xnor2_1 _26619_ (.Y(_04958_),
    .A(_00172_),
    .B(_04957_));
 sg13g2_o21ai_1 _26620_ (.B1(_04958_),
    .Y(_04959_),
    .A1(_04866_),
    .A2(_04954_));
 sg13g2_nand2_1 _26621_ (.Y(_04960_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[15] ),
    .B(_04957_));
 sg13g2_xnor2_1 _26622_ (.Y(_04961_),
    .A(_11416_),
    .B(_04820_));
 sg13g2_nand2_1 _26623_ (.Y(_04962_),
    .A(_11416_),
    .B(net8480));
 sg13g2_o21ai_1 _26624_ (.B1(_04962_),
    .Y(_04963_),
    .A1(net8480),
    .A2(_04961_));
 sg13g2_xnor2_1 _26625_ (.Y(_04964_),
    .A(_00171_),
    .B(_04963_));
 sg13g2_inv_1 _26626_ (.Y(_04965_),
    .A(_04964_));
 sg13g2_a21oi_1 _26627_ (.A1(_04959_),
    .A2(_04960_),
    .Y(_04966_),
    .B1(_04965_));
 sg13g2_a21oi_1 _26628_ (.A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[16] ),
    .A2(_04963_),
    .Y(_04967_),
    .B1(_04966_));
 sg13g2_xor2_1 _26629_ (.B(_04821_),
    .A(net8379),
    .X(_04968_));
 sg13g2_and2_1 _26630_ (.A(net8379),
    .B(net8476),
    .X(_04969_));
 sg13g2_a21oi_2 _26631_ (.B1(_04969_),
    .Y(_04970_),
    .A2(_04968_),
    .A1(net8483));
 sg13g2_xnor2_1 _26632_ (.Y(_04971_),
    .A(_00170_),
    .B(_04970_));
 sg13g2_nor2b_1 _26633_ (.A(_04967_),
    .B_N(_04971_),
    .Y(_04972_));
 sg13g2_a21o_1 _26634_ (.A2(_04970_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[17] ),
    .B1(_04972_),
    .X(_04973_));
 sg13g2_xor2_1 _26635_ (.B(_04822_),
    .A(_11404_),
    .X(_04974_));
 sg13g2_nor2_1 _26636_ (.A(net8477),
    .B(_04974_),
    .Y(_04975_));
 sg13g2_a21oi_2 _26637_ (.B1(_04975_),
    .Y(_04976_),
    .A2(net8477),
    .A1(_11404_));
 sg13g2_xnor2_1 _26638_ (.Y(_04977_),
    .A(_00169_),
    .B(_04976_));
 sg13g2_a22oi_1 _26639_ (.Y(_04978_),
    .B1(_04977_),
    .B2(_04973_),
    .A2(_04976_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[18] ));
 sg13g2_xnor2_1 _26640_ (.Y(_04979_),
    .A(_00168_),
    .B(_04862_));
 sg13g2_nor2b_1 _26641_ (.A(_04978_),
    .B_N(_04979_),
    .Y(_04980_));
 sg13g2_a21o_1 _26642_ (.A2(_04862_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[19] ),
    .B1(_04980_),
    .X(_04981_));
 sg13g2_nand2_1 _26643_ (.Y(_04982_),
    .A(_04859_),
    .B(_04981_));
 sg13g2_xor2_1 _26644_ (.B(_04853_),
    .A(_00166_),
    .X(_04983_));
 sg13g2_a21o_1 _26645_ (.A2(_04982_),
    .A1(_04858_),
    .B1(_04983_),
    .X(_04984_));
 sg13g2_a21oi_1 _26646_ (.A1(_04854_),
    .A2(_04984_),
    .Y(_04985_),
    .B1(_04850_));
 sg13g2_a21o_1 _26647_ (.A2(_04849_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[22] ),
    .B1(_04985_),
    .X(_04986_));
 sg13g2_xnor2_1 _26648_ (.Y(_04987_),
    .A(_11465_),
    .B(_04827_));
 sg13g2_nor2_1 _26649_ (.A(net8476),
    .B(_04987_),
    .Y(_04988_));
 sg13g2_a21oi_2 _26650_ (.B1(_04988_),
    .Y(_04989_),
    .A2(net8476),
    .A1(_11465_));
 sg13g2_xnor2_1 _26651_ (.Y(_04990_),
    .A(_00164_),
    .B(_04989_));
 sg13g2_a22oi_1 _26652_ (.Y(_04991_),
    .B1(_04990_),
    .B2(_04986_),
    .A2(_04989_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[23] ));
 sg13g2_xnor2_1 _26653_ (.Y(_04992_),
    .A(_00163_),
    .B(_04846_));
 sg13g2_nor2b_1 _26654_ (.A(_04991_),
    .B_N(_04992_),
    .Y(_04993_));
 sg13g2_a21o_1 _26655_ (.A2(_04846_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[24] ),
    .B1(_04993_),
    .X(_04994_));
 sg13g2_xnor2_1 _26656_ (.Y(_04995_),
    .A(net8006),
    .B(_04829_));
 sg13g2_nor2_1 _26657_ (.A(net8476),
    .B(_04995_),
    .Y(_04996_));
 sg13g2_a21oi_2 _26658_ (.B1(_04996_),
    .Y(_04997_),
    .A2(net8476),
    .A1(net8006));
 sg13g2_xnor2_1 _26659_ (.Y(_04998_),
    .A(_00162_),
    .B(_04997_));
 sg13g2_a22oi_1 _26660_ (.Y(_04999_),
    .B1(_04998_),
    .B2(_04994_),
    .A2(_04997_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[25] ));
 sg13g2_xnor2_1 _26661_ (.Y(_05000_),
    .A(_00161_),
    .B(_04843_));
 sg13g2_nor2b_1 _26662_ (.A(_04999_),
    .B_N(_05000_),
    .Y(_05001_));
 sg13g2_a21o_1 _26663_ (.A2(_04843_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[26] ),
    .B1(_05001_),
    .X(_05002_));
 sg13g2_xnor2_1 _26664_ (.Y(_05003_),
    .A(_11495_),
    .B(_04831_));
 sg13g2_nor2_1 _26665_ (.A(_11495_),
    .B(net8485),
    .Y(_05004_));
 sg13g2_a21oi_2 _26666_ (.B1(_05004_),
    .Y(_05005_),
    .A2(_05003_),
    .A1(net8485));
 sg13g2_xnor2_1 _26667_ (.Y(_05006_),
    .A(_00160_),
    .B(_05005_));
 sg13g2_nand2_1 _26668_ (.Y(_05007_),
    .A(_05002_),
    .B(_05006_));
 sg13g2_nand2_1 _26669_ (.Y(_05008_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[27] ),
    .B(_05005_));
 sg13g2_xor2_1 _26670_ (.B(_04840_),
    .A(_00159_),
    .X(_05009_));
 sg13g2_a21oi_1 _26671_ (.A1(_05007_),
    .A2(_05008_),
    .Y(_05010_),
    .B1(_05009_));
 sg13g2_a21oi_1 _26672_ (.A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[28] ),
    .A2(_04840_),
    .Y(_05011_),
    .B1(_05010_));
 sg13g2_xnor2_1 _26673_ (.Y(_05012_),
    .A(net8008),
    .B(_04833_));
 sg13g2_nor2_1 _26674_ (.A(net8482),
    .B(_05012_),
    .Y(_05013_));
 sg13g2_a21oi_2 _26675_ (.B1(_05013_),
    .Y(_05014_),
    .A2(net8482),
    .A1(net8008));
 sg13g2_xor2_1 _26676_ (.B(_05014_),
    .A(_00158_),
    .X(_05015_));
 sg13g2_nand2_1 _26677_ (.Y(_05016_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[29] ),
    .B(_05014_));
 sg13g2_o21ai_1 _26678_ (.B1(_05016_),
    .Y(_05017_),
    .A1(_05011_),
    .A2(_05015_));
 sg13g2_a21o_1 _26679_ (.A2(_04835_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[30] ),
    .B1(_05017_),
    .X(_05018_));
 sg13g2_nand2b_1 _26680_ (.Y(_05019_),
    .B(_10514_),
    .A_N(_04835_));
 sg13g2_and2_2 _26681_ (.A(_05018_),
    .B(_05019_),
    .X(_05020_));
 sg13g2_and2_1 _26682_ (.A(net9229),
    .B(_05020_),
    .X(_05021_));
 sg13g2_nand2_2 _26683_ (.Y(_05022_),
    .A(net9229),
    .B(_05020_));
 sg13g2_nand3b_1 _26684_ (.B(_13831_),
    .C(net9698),
    .Y(_05023_),
    .A_N(\soc_I.kianv_I.control_unit_I.div_ready ));
 sg13g2_nand2_2 _26685_ (.Y(_05024_),
    .A(net5490),
    .B(_05023_));
 sg13g2_nor2_1 _26686_ (.A(net9238),
    .B(net9228),
    .Y(_05025_));
 sg13g2_or2_1 _26687_ (.X(_05026_),
    .B(net9228),
    .A(net9238));
 sg13g2_nor2_1 _26688_ (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_state[0] ),
    .B(net9226),
    .Y(_05027_));
 sg13g2_o21ai_1 _26689_ (.B1(_05024_),
    .Y(_05028_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_state[0] ),
    .A2(net8939));
 sg13g2_nand2_1 _26690_ (.Y(_05029_),
    .A(_11022_),
    .B(_04834_));
 sg13g2_nand3_1 _26691_ (.B(_04806_),
    .C(_05029_),
    .A(_11600_),
    .Y(_05030_));
 sg13g2_a21oi_1 _26692_ (.A1(net9237),
    .A2(_05030_),
    .Y(_05031_),
    .B1(_05028_));
 sg13g2_a22oi_1 _26693_ (.Y(_05032_),
    .B1(_11186_),
    .B2(net8940),
    .A2(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[0] ),
    .A1(net9239));
 sg13g2_nand3_1 _26694_ (.B(net7387),
    .C(_05032_),
    .A(net7330),
    .Y(_05033_));
 sg13g2_o21ai_1 _26695_ (.B1(net9418),
    .Y(_05034_),
    .A1(net5560),
    .A2(net7387));
 sg13g2_nor2b_1 _26696_ (.A(_05034_),
    .B_N(_05033_),
    .Y(_01201_));
 sg13g2_o21ai_1 _26697_ (.B1(net9239),
    .Y(_05035_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[1] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[0] ));
 sg13g2_a21oi_1 _26698_ (.A1(net5414),
    .A2(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[0] ),
    .Y(_05036_),
    .B1(_05035_));
 sg13g2_nor2_2 _26699_ (.A(net8315),
    .B(_04807_),
    .Y(_05037_));
 sg13g2_nand2_1 _26700_ (.Y(_05038_),
    .A(_10993_),
    .B(_04806_));
 sg13g2_nor2_1 _26701_ (.A(net8299),
    .B(_11186_),
    .Y(_05039_));
 sg13g2_xnor2_1 _26702_ (.Y(_05040_),
    .A(net8299),
    .B(net8298));
 sg13g2_nor2_1 _26703_ (.A(net7982),
    .B(_05040_),
    .Y(_05041_));
 sg13g2_a21oi_1 _26704_ (.A1(_11160_),
    .A2(net7982),
    .Y(_05042_),
    .B1(_05041_));
 sg13g2_a221oi_1 _26705_ (.B2(_05042_),
    .C1(_05036_),
    .B1(net8940),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[0] ),
    .Y(_05043_),
    .A2(net9225));
 sg13g2_o21ai_1 _26706_ (.B1(net9414),
    .Y(_05044_),
    .A1(net5414),
    .A2(net7388));
 sg13g2_a21oi_1 _26707_ (.A1(net7388),
    .A2(_05043_),
    .Y(_01202_),
    .B1(_05044_));
 sg13g2_nand2_1 _26708_ (.Y(_05045_),
    .A(_11143_),
    .B(_05039_));
 sg13g2_xnor2_1 _26709_ (.Y(_05046_),
    .A(_11143_),
    .B(_05039_));
 sg13g2_o21ai_1 _26710_ (.B1(net8940),
    .Y(_05047_),
    .A1(_11144_),
    .A2(net7986));
 sg13g2_a21oi_1 _26711_ (.A1(net7983),
    .A2(_05046_),
    .Y(_05048_),
    .B1(_05047_));
 sg13g2_or3_1 _26712_ (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[2] ),
    .B(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[1] ),
    .C(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[0] ),
    .X(_05049_));
 sg13g2_o21ai_1 _26713_ (.B1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[2] ),
    .Y(_05050_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[1] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[0] ));
 sg13g2_and2_1 _26714_ (.A(net9239),
    .B(_05050_),
    .X(_05051_));
 sg13g2_a221oi_1 _26715_ (.B2(_05051_),
    .C1(_05048_),
    .B1(_05049_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[1] ),
    .Y(_05052_),
    .A2(net9224));
 sg13g2_o21ai_1 _26716_ (.B1(net9414),
    .Y(_05053_),
    .A1(net5402),
    .A2(net7379));
 sg13g2_a21oi_1 _26717_ (.A1(net7379),
    .A2(_05052_),
    .Y(_01203_),
    .B1(_05053_));
 sg13g2_or2_1 _26718_ (.X(_05054_),
    .B(_05045_),
    .A(net8302));
 sg13g2_xnor2_1 _26719_ (.Y(_05055_),
    .A(net8301),
    .B(_05045_));
 sg13g2_o21ai_1 _26720_ (.B1(net8940),
    .Y(_05056_),
    .A1(net8301),
    .A2(net7983));
 sg13g2_a21oi_1 _26721_ (.A1(net7983),
    .A2(_05055_),
    .Y(_05057_),
    .B1(_05056_));
 sg13g2_or2_1 _26722_ (.X(_05058_),
    .B(_05049_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[3] ));
 sg13g2_a21oi_1 _26723_ (.A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[3] ),
    .A2(_05049_),
    .Y(_05059_),
    .B1(net9062));
 sg13g2_a221oi_1 _26724_ (.B2(_05059_),
    .C1(_05057_),
    .B1(_05058_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[2] ),
    .Y(_05060_),
    .A2(net9224));
 sg13g2_o21ai_1 _26725_ (.B1(net9414),
    .Y(_05061_),
    .A1(net5325),
    .A2(net7379));
 sg13g2_a21oi_1 _26726_ (.A1(net7379),
    .A2(_05060_),
    .Y(_01204_),
    .B1(_05061_));
 sg13g2_or2_1 _26727_ (.X(_05062_),
    .B(_05054_),
    .A(_11118_));
 sg13g2_xnor2_1 _26728_ (.Y(_05063_),
    .A(_11117_),
    .B(_05054_));
 sg13g2_o21ai_1 _26729_ (.B1(net8941),
    .Y(_05064_),
    .A1(net7982),
    .A2(_05063_));
 sg13g2_a21oi_1 _26730_ (.A1(net8303),
    .A2(net7982),
    .Y(_05065_),
    .B1(_05064_));
 sg13g2_or2_1 _26731_ (.X(_05066_),
    .B(_05058_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[4] ));
 sg13g2_a21oi_1 _26732_ (.A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[4] ),
    .A2(_05058_),
    .Y(_05067_),
    .B1(net9062));
 sg13g2_a221oi_1 _26733_ (.B2(_05067_),
    .C1(_05065_),
    .B1(_05066_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[3] ),
    .Y(_05068_),
    .A2(net9224));
 sg13g2_o21ai_1 _26734_ (.B1(net9415),
    .Y(_05069_),
    .A1(net5290),
    .A2(net7378));
 sg13g2_a21oi_1 _26735_ (.A1(net7378),
    .A2(_05068_),
    .Y(_01205_),
    .B1(_05069_));
 sg13g2_xnor2_1 _26736_ (.Y(_05070_),
    .A(net8305),
    .B(_05062_));
 sg13g2_nor2_1 _26737_ (.A(net8305),
    .B(net7984),
    .Y(_05071_));
 sg13g2_a21oi_1 _26738_ (.A1(net7984),
    .A2(_05070_),
    .Y(_05072_),
    .B1(_05071_));
 sg13g2_o21ai_1 _26739_ (.B1(net9239),
    .Y(_05073_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[5] ),
    .A2(_05066_));
 sg13g2_a21oi_1 _26740_ (.A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[5] ),
    .A2(_05066_),
    .Y(_05074_),
    .B1(_05073_));
 sg13g2_a221oi_1 _26741_ (.B2(_05072_),
    .C1(_05074_),
    .B1(net8940),
    .A1(net5290),
    .Y(_05075_),
    .A2(net9224));
 sg13g2_o21ai_1 _26742_ (.B1(net9415),
    .Y(_05076_),
    .A1(net5447),
    .A2(net7376));
 sg13g2_a21oi_1 _26743_ (.A1(net7376),
    .A2(_05075_),
    .Y(_01206_),
    .B1(_05076_));
 sg13g2_nor3_2 _26744_ (.A(_11096_),
    .B(net8305),
    .C(_05062_),
    .Y(_05077_));
 sg13g2_o21ai_1 _26745_ (.B1(_11096_),
    .Y(_05078_),
    .A1(net8304),
    .A2(_05062_));
 sg13g2_nand2b_1 _26746_ (.Y(_05079_),
    .B(_05078_),
    .A_N(_05077_));
 sg13g2_o21ai_1 _26747_ (.B1(net8940),
    .Y(_05080_),
    .A1(_11096_),
    .A2(net7983));
 sg13g2_a21oi_1 _26748_ (.A1(net7983),
    .A2(_05079_),
    .Y(_05081_),
    .B1(_05080_));
 sg13g2_nor3_1 _26749_ (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[6] ),
    .B(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[5] ),
    .C(_05066_),
    .Y(_05082_));
 sg13g2_o21ai_1 _26750_ (.B1(net5256),
    .Y(_05083_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[5] ),
    .A2(_05066_));
 sg13g2_nor2_1 _26751_ (.A(net9062),
    .B(_05082_),
    .Y(_05084_));
 sg13g2_a221oi_1 _26752_ (.B2(_05084_),
    .C1(_05081_),
    .B1(_05083_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[5] ),
    .Y(_05085_),
    .A2(net9224));
 sg13g2_o21ai_1 _26753_ (.B1(net9415),
    .Y(_05086_),
    .A1(net5256),
    .A2(net7376));
 sg13g2_a21oi_1 _26754_ (.A1(net7376),
    .A2(_05085_),
    .Y(_01207_),
    .B1(_05086_));
 sg13g2_and2_1 _26755_ (.A(_11087_),
    .B(_05077_),
    .X(_05087_));
 sg13g2_xnor2_1 _26756_ (.Y(_05088_),
    .A(_11087_),
    .B(_05077_));
 sg13g2_o21ai_1 _26757_ (.B1(net8942),
    .Y(_05089_),
    .A1(_11086_),
    .A2(net7986));
 sg13g2_a21oi_1 _26758_ (.A1(net7986),
    .A2(_05088_),
    .Y(_05090_),
    .B1(_05089_));
 sg13g2_nand2b_1 _26759_ (.Y(_05091_),
    .B(_05082_),
    .A_N(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[7] ));
 sg13g2_nor2b_1 _26760_ (.A(_05082_),
    .B_N(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[7] ),
    .Y(_05092_));
 sg13g2_nor2_1 _26761_ (.A(net9062),
    .B(_05092_),
    .Y(_05093_));
 sg13g2_a221oi_1 _26762_ (.B2(_05093_),
    .C1(_05090_),
    .B1(_05091_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[6] ),
    .Y(_05094_),
    .A2(net9225));
 sg13g2_o21ai_1 _26763_ (.B1(net9414),
    .Y(_05095_),
    .A1(net5283),
    .A2(net7376));
 sg13g2_a21oi_1 _26764_ (.A1(net7376),
    .A2(_05094_),
    .Y(_01208_),
    .B1(_05095_));
 sg13g2_nand2_1 _26765_ (.Y(_05096_),
    .A(_11207_),
    .B(_05087_));
 sg13g2_xnor2_1 _26766_ (.Y(_05097_),
    .A(_11207_),
    .B(_05087_));
 sg13g2_o21ai_1 _26767_ (.B1(net8942),
    .Y(_05098_),
    .A1(_11208_),
    .A2(net7986));
 sg13g2_a21oi_1 _26768_ (.A1(net7986),
    .A2(_05097_),
    .Y(_05099_),
    .B1(_05098_));
 sg13g2_or2_1 _26769_ (.X(_05100_),
    .B(_05091_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[8] ));
 sg13g2_a21oi_1 _26770_ (.A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[8] ),
    .A2(_05091_),
    .Y(_05101_),
    .B1(net9062));
 sg13g2_a221oi_1 _26771_ (.B2(_05101_),
    .C1(_05099_),
    .B1(_05100_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[7] ),
    .Y(_05102_),
    .A2(net9225));
 sg13g2_o21ai_1 _26772_ (.B1(net9414),
    .Y(_05103_),
    .A1(net5230),
    .A2(net7376));
 sg13g2_a21oi_1 _26773_ (.A1(net7376),
    .A2(_05102_),
    .Y(_01209_),
    .B1(_05103_));
 sg13g2_nand3_1 _26774_ (.B(_11246_),
    .C(_05087_),
    .A(_11207_),
    .Y(_05104_));
 sg13g2_xnor2_1 _26775_ (.Y(_05105_),
    .A(_11247_),
    .B(_05096_));
 sg13g2_nor2_1 _26776_ (.A(_11247_),
    .B(net7984),
    .Y(_05106_));
 sg13g2_a21oi_1 _26777_ (.A1(net7983),
    .A2(_05105_),
    .Y(_05107_),
    .B1(_05106_));
 sg13g2_nor2_2 _26778_ (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[9] ),
    .B(_05100_),
    .Y(_05108_));
 sg13g2_a21oi_1 _26779_ (.A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[9] ),
    .A2(_05100_),
    .Y(_05109_),
    .B1(net9062));
 sg13g2_nor2b_1 _26780_ (.A(_05108_),
    .B_N(_05109_),
    .Y(_05110_));
 sg13g2_a221oi_1 _26781_ (.B2(_05107_),
    .C1(_05110_),
    .B1(net8940),
    .A1(net5230),
    .Y(_05111_),
    .A2(net9224));
 sg13g2_o21ai_1 _26782_ (.B1(net9414),
    .Y(_05112_),
    .A1(net5301),
    .A2(net7377));
 sg13g2_a21oi_1 _26783_ (.A1(net7377),
    .A2(_05111_),
    .Y(_01210_),
    .B1(_05112_));
 sg13g2_or2_1 _26784_ (.X(_05113_),
    .B(_05104_),
    .A(_11222_));
 sg13g2_xnor2_1 _26785_ (.Y(_05114_),
    .A(_11222_),
    .B(_05104_));
 sg13g2_o21ai_1 _26786_ (.B1(net8940),
    .Y(_05115_),
    .A1(_11222_),
    .A2(net7984));
 sg13g2_a21oi_1 _26787_ (.A1(net7983),
    .A2(_05114_),
    .Y(_05116_),
    .B1(_05115_));
 sg13g2_nand2b_2 _26788_ (.Y(_05117_),
    .B(_05108_),
    .A_N(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[10] ));
 sg13g2_nor2b_1 _26789_ (.A(_05108_),
    .B_N(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[10] ),
    .Y(_05118_));
 sg13g2_nor2_1 _26790_ (.A(net9062),
    .B(_05118_),
    .Y(_05119_));
 sg13g2_a221oi_1 _26791_ (.B2(_05119_),
    .C1(_05116_),
    .B1(_05117_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[9] ),
    .Y(_05120_),
    .A2(net9224));
 sg13g2_o21ai_1 _26792_ (.B1(net9414),
    .Y(_05121_),
    .A1(net5224),
    .A2(net7377));
 sg13g2_a21oi_1 _26793_ (.A1(net7377),
    .A2(_05120_),
    .Y(_01211_),
    .B1(_05121_));
 sg13g2_nor2_1 _26794_ (.A(net8297),
    .B(_05113_),
    .Y(_05122_));
 sg13g2_xnor2_1 _26795_ (.Y(_05123_),
    .A(net8297),
    .B(_05113_));
 sg13g2_nor2_1 _26796_ (.A(net8297),
    .B(net7984),
    .Y(_05124_));
 sg13g2_a21oi_1 _26797_ (.A1(net7983),
    .A2(_05123_),
    .Y(_05125_),
    .B1(_05124_));
 sg13g2_o21ai_1 _26798_ (.B1(net9239),
    .Y(_05126_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[11] ),
    .A2(_05117_));
 sg13g2_a21oi_1 _26799_ (.A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[11] ),
    .A2(_05117_),
    .Y(_05127_),
    .B1(_05126_));
 sg13g2_a221oi_1 _26800_ (.B2(_05125_),
    .C1(_05127_),
    .B1(net8941),
    .A1(net5224),
    .Y(_05128_),
    .A2(net9224));
 sg13g2_o21ai_1 _26801_ (.B1(net9414),
    .Y(_05129_),
    .A1(net5502),
    .A2(net7377));
 sg13g2_a21oi_1 _26802_ (.A1(net7377),
    .A2(_05128_),
    .Y(_01212_),
    .B1(_05129_));
 sg13g2_nor3_2 _26803_ (.A(net8296),
    .B(net8292),
    .C(_05113_),
    .Y(_05130_));
 sg13g2_xnor2_1 _26804_ (.Y(_05131_),
    .A(_11292_),
    .B(_05122_));
 sg13g2_o21ai_1 _26805_ (.B1(net8941),
    .Y(_05132_),
    .A1(net8292),
    .A2(net7985));
 sg13g2_a21oi_1 _26806_ (.A1(net7985),
    .A2(_05131_),
    .Y(_05133_),
    .B1(_05132_));
 sg13g2_nor3_2 _26807_ (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[12] ),
    .B(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[11] ),
    .C(_05117_),
    .Y(_05134_));
 sg13g2_o21ai_1 _26808_ (.B1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[12] ),
    .Y(_05135_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[11] ),
    .A2(_05117_));
 sg13g2_nor2_1 _26809_ (.A(net9064),
    .B(_05134_),
    .Y(_05136_));
 sg13g2_a221oi_1 _26810_ (.B2(_05136_),
    .C1(_05133_),
    .B1(_05135_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[11] ),
    .Y(_05137_),
    .A2(net9231));
 sg13g2_o21ai_1 _26811_ (.B1(net9418),
    .Y(_05138_),
    .A1(net5473),
    .A2(net7380));
 sg13g2_a21oi_1 _26812_ (.A1(net7380),
    .A2(_05137_),
    .Y(_01213_),
    .B1(_05138_));
 sg13g2_nand2_1 _26813_ (.Y(_05139_),
    .A(net8291),
    .B(_05130_));
 sg13g2_xnor2_1 _26814_ (.Y(_05140_),
    .A(net8291),
    .B(_05130_));
 sg13g2_o21ai_1 _26815_ (.B1(net8942),
    .Y(_05141_),
    .A1(_11304_),
    .A2(net7986));
 sg13g2_a21oi_1 _26816_ (.A1(net7985),
    .A2(_05140_),
    .Y(_05142_),
    .B1(_05141_));
 sg13g2_nand2b_2 _26817_ (.Y(_05143_),
    .B(_05134_),
    .A_N(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[13] ));
 sg13g2_nor2b_1 _26818_ (.A(_05134_),
    .B_N(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[13] ),
    .Y(_05144_));
 sg13g2_nor2_1 _26819_ (.A(net9062),
    .B(_05144_),
    .Y(_05145_));
 sg13g2_a221oi_1 _26820_ (.B2(_05145_),
    .C1(_05142_),
    .B1(_05143_),
    .A1(net5473),
    .Y(_05146_),
    .A2(net9231));
 sg13g2_o21ai_1 _26821_ (.B1(net9418),
    .Y(_05147_),
    .A1(net5520),
    .A2(net7380));
 sg13g2_a21oi_1 _26822_ (.A1(net7380),
    .A2(_05146_),
    .Y(_01214_),
    .B1(_05147_));
 sg13g2_nand3_1 _26823_ (.B(net8291),
    .C(_05130_),
    .A(net8295),
    .Y(_05148_));
 sg13g2_xnor2_1 _26824_ (.Y(_05149_),
    .A(_11268_),
    .B(_05139_));
 sg13g2_nand2_1 _26825_ (.Y(_05150_),
    .A(net8295),
    .B(net7981));
 sg13g2_a21oi_1 _26826_ (.A1(net7988),
    .A2(_05149_),
    .Y(_05151_),
    .B1(net8939));
 sg13g2_o21ai_1 _26827_ (.B1(net9238),
    .Y(_05152_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[14] ),
    .A2(_05143_));
 sg13g2_a21oi_1 _26828_ (.A1(net5580),
    .A2(_05143_),
    .Y(_05153_),
    .B1(_05152_));
 sg13g2_a221oi_1 _26829_ (.B2(_05151_),
    .C1(_05153_),
    .B1(_05150_),
    .A1(net5567),
    .Y(_05154_),
    .A2(net9230));
 sg13g2_o21ai_1 _26830_ (.B1(net9418),
    .Y(_05155_),
    .A1(net5437),
    .A2(net7386));
 sg13g2_a21oi_1 _26831_ (.A1(net7386),
    .A2(_05154_),
    .Y(_01215_),
    .B1(_05155_));
 sg13g2_or2_1 _26832_ (.X(_05156_),
    .B(_05148_),
    .A(net8294));
 sg13g2_xnor2_1 _26833_ (.Y(_05157_),
    .A(net8293),
    .B(_05148_));
 sg13g2_o21ai_1 _26834_ (.B1(net8944),
    .Y(_05158_),
    .A1(net8293),
    .A2(net7988));
 sg13g2_a21oi_1 _26835_ (.A1(net7988),
    .A2(_05157_),
    .Y(_05159_),
    .B1(_05158_));
 sg13g2_nor3_2 _26836_ (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[15] ),
    .B(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[14] ),
    .C(_05143_),
    .Y(_05160_));
 sg13g2_o21ai_1 _26837_ (.B1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[15] ),
    .Y(_05161_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[14] ),
    .A2(_05143_));
 sg13g2_nor2_1 _26838_ (.A(net9064),
    .B(_05160_),
    .Y(_05162_));
 sg13g2_a221oi_1 _26839_ (.B2(_05162_),
    .C1(_05159_),
    .B1(_05161_),
    .A1(net5437),
    .Y(_05163_),
    .A2(net9228));
 sg13g2_o21ai_1 _26840_ (.B1(net9418),
    .Y(_05164_),
    .A1(net5446),
    .A2(net7384));
 sg13g2_a21oi_1 _26841_ (.A1(net7384),
    .A2(_05163_),
    .Y(_01216_),
    .B1(_05164_));
 sg13g2_or2_1 _26842_ (.X(_05165_),
    .B(_05156_),
    .A(_11379_));
 sg13g2_xnor2_1 _26843_ (.Y(_05166_),
    .A(_11379_),
    .B(_05156_));
 sg13g2_nand2_1 _26844_ (.Y(_05167_),
    .A(net8283),
    .B(net7981));
 sg13g2_a21oi_1 _26845_ (.A1(net7988),
    .A2(_05166_),
    .Y(_05168_),
    .B1(net8939));
 sg13g2_nand2b_2 _26846_ (.Y(_05169_),
    .B(_05160_),
    .A_N(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[16] ));
 sg13g2_nand2b_1 _26847_ (.Y(_05170_),
    .B(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[16] ),
    .A_N(_05160_));
 sg13g2_and3_1 _26848_ (.X(_05171_),
    .A(net9238),
    .B(_05169_),
    .C(_05170_));
 sg13g2_a221oi_1 _26849_ (.B2(_05168_),
    .C1(_05171_),
    .B1(_05167_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[15] ),
    .Y(_05172_),
    .A2(net9228));
 sg13g2_o21ai_1 _26850_ (.B1(net9417),
    .Y(_05173_),
    .A1(net5305),
    .A2(net7386));
 sg13g2_a21oi_1 _26851_ (.A1(net7385),
    .A2(_05172_),
    .Y(_01217_),
    .B1(_05173_));
 sg13g2_nor2_2 _26852_ (.A(net8276),
    .B(_05165_),
    .Y(_05174_));
 sg13g2_xnor2_1 _26853_ (.Y(_05175_),
    .A(net8276),
    .B(_05165_));
 sg13g2_nor2_1 _26854_ (.A(net8276),
    .B(net7987),
    .Y(_05176_));
 sg13g2_a21oi_1 _26855_ (.A1(net7988),
    .A2(_05175_),
    .Y(_05177_),
    .B1(_05176_));
 sg13g2_nor2_1 _26856_ (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[17] ),
    .B(_05169_),
    .Y(_05178_));
 sg13g2_a21oi_1 _26857_ (.A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[17] ),
    .A2(_05169_),
    .Y(_05179_),
    .B1(net9063));
 sg13g2_nor2b_1 _26858_ (.A(_05178_),
    .B_N(_05179_),
    .Y(_05180_));
 sg13g2_a221oi_1 _26859_ (.B2(_05177_),
    .C1(_05180_),
    .B1(net8943),
    .A1(net5305),
    .Y(_05181_),
    .A2(net9228));
 sg13g2_o21ai_1 _26860_ (.B1(net9418),
    .Y(_05182_),
    .A1(net5478),
    .A2(net7384));
 sg13g2_a21oi_1 _26861_ (.A1(net7384),
    .A2(_05181_),
    .Y(_01218_),
    .B1(_05182_));
 sg13g2_nand2_1 _26862_ (.Y(_05183_),
    .A(net8282),
    .B(_05174_));
 sg13g2_xnor2_1 _26863_ (.Y(_05184_),
    .A(net8281),
    .B(_05174_));
 sg13g2_nand2_1 _26864_ (.Y(_05185_),
    .A(net8281),
    .B(net7981));
 sg13g2_a21oi_1 _26865_ (.A1(net7987),
    .A2(_05184_),
    .Y(_05186_),
    .B1(_05026_));
 sg13g2_nor3_2 _26866_ (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[18] ),
    .B(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[17] ),
    .C(_05169_),
    .Y(_05187_));
 sg13g2_nor2b_1 _26867_ (.A(_05178_),
    .B_N(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[18] ),
    .Y(_05188_));
 sg13g2_nor3_1 _26868_ (.A(net9064),
    .B(_05187_),
    .C(_05188_),
    .Y(_05189_));
 sg13g2_a221oi_1 _26869_ (.B2(_05186_),
    .C1(_05189_),
    .B1(_05185_),
    .A1(net5488),
    .Y(_05190_),
    .A2(net9228));
 sg13g2_o21ai_1 _26870_ (.B1(net9417),
    .Y(_05191_),
    .A1(net5360),
    .A2(net7384));
 sg13g2_a21oi_1 _26871_ (.A1(net7384),
    .A2(_05190_),
    .Y(_01219_),
    .B1(_05191_));
 sg13g2_nand3_1 _26872_ (.B(_11402_),
    .C(_05174_),
    .A(net8281),
    .Y(_05192_));
 sg13g2_xnor2_1 _26873_ (.Y(_05193_),
    .A(net8279),
    .B(_05183_));
 sg13g2_o21ai_1 _26874_ (.B1(net8944),
    .Y(_05194_),
    .A1(net8279),
    .A2(net7987));
 sg13g2_a21oi_1 _26875_ (.A1(net7988),
    .A2(_05193_),
    .Y(_05195_),
    .B1(_05194_));
 sg13g2_nand2b_2 _26876_ (.Y(_05196_),
    .B(_05187_),
    .A_N(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[19] ));
 sg13g2_nor2b_1 _26877_ (.A(_05187_),
    .B_N(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[19] ),
    .Y(_05197_));
 sg13g2_nor2_1 _26878_ (.A(net9064),
    .B(_05197_),
    .Y(_05198_));
 sg13g2_a221oi_1 _26879_ (.B2(_05198_),
    .C1(_05195_),
    .B1(_05196_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[18] ),
    .Y(_05199_),
    .A2(net9228));
 sg13g2_o21ai_1 _26880_ (.B1(net9417),
    .Y(_05200_),
    .A1(net5212),
    .A2(net7384));
 sg13g2_a21oi_1 _26881_ (.A1(net7384),
    .A2(_05199_),
    .Y(_01220_),
    .B1(_05200_));
 sg13g2_or2_1 _26882_ (.X(_05201_),
    .B(_05192_),
    .A(_11350_));
 sg13g2_xnor2_1 _26883_ (.Y(_05202_),
    .A(_11350_),
    .B(_05192_));
 sg13g2_nand2_1 _26884_ (.Y(_05203_),
    .A(net8286),
    .B(net7981));
 sg13g2_a21oi_1 _26885_ (.A1(net7987),
    .A2(_05202_),
    .Y(_05204_),
    .B1(net8939));
 sg13g2_o21ai_1 _26886_ (.B1(net9238),
    .Y(_05205_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[20] ),
    .A2(_05196_));
 sg13g2_a21oi_1 _26887_ (.A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[20] ),
    .A2(_05196_),
    .Y(_05206_),
    .B1(_05205_));
 sg13g2_a221oi_1 _26888_ (.B2(_05204_),
    .C1(_05206_),
    .B1(_05203_),
    .A1(net5212),
    .Y(_05207_),
    .A2(net9228));
 sg13g2_o21ai_1 _26889_ (.B1(net9417),
    .Y(_05208_),
    .A1(net5463),
    .A2(net7385));
 sg13g2_a21oi_1 _26890_ (.A1(net7385),
    .A2(_05207_),
    .Y(_01221_),
    .B1(_05208_));
 sg13g2_or2_1 _26891_ (.X(_05209_),
    .B(_05201_),
    .A(net8284));
 sg13g2_xnor2_1 _26892_ (.Y(_05210_),
    .A(net8284),
    .B(_05201_));
 sg13g2_o21ai_1 _26893_ (.B1(net8944),
    .Y(_05211_),
    .A1(net8285),
    .A2(net7987));
 sg13g2_a21oi_1 _26894_ (.A1(net7987),
    .A2(_05210_),
    .Y(_05212_),
    .B1(_05211_));
 sg13g2_nor3_2 _26895_ (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[21] ),
    .B(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[20] ),
    .C(_05196_),
    .Y(_05213_));
 sg13g2_o21ai_1 _26896_ (.B1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[21] ),
    .Y(_05214_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[20] ),
    .A2(_05196_));
 sg13g2_nor2_1 _26897_ (.A(net9063),
    .B(_05213_),
    .Y(_05215_));
 sg13g2_a221oi_1 _26898_ (.B2(_05215_),
    .C1(_05212_),
    .B1(_05214_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[20] ),
    .Y(_05216_),
    .A2(net9230));
 sg13g2_o21ai_1 _26899_ (.B1(net9417),
    .Y(_05217_),
    .A1(net5392),
    .A2(net7385));
 sg13g2_a21oi_1 _26900_ (.A1(net7385),
    .A2(_05216_),
    .Y(_01222_),
    .B1(_05217_));
 sg13g2_or2_1 _26901_ (.X(_05218_),
    .B(_05209_),
    .A(_11323_));
 sg13g2_xnor2_1 _26902_ (.Y(_05219_),
    .A(_11323_),
    .B(_05209_));
 sg13g2_nand2_1 _26903_ (.Y(_05220_),
    .A(net8288),
    .B(net7981));
 sg13g2_a21oi_1 _26904_ (.A1(net7987),
    .A2(_05219_),
    .Y(_05221_),
    .B1(net8939));
 sg13g2_nand2b_2 _26905_ (.Y(_05222_),
    .B(_05213_),
    .A_N(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[22] ));
 sg13g2_nand2b_1 _26906_ (.Y(_05223_),
    .B(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[22] ),
    .A_N(_05213_));
 sg13g2_and3_1 _26907_ (.X(_05224_),
    .A(net9238),
    .B(_05222_),
    .C(_05223_));
 sg13g2_a221oi_1 _26908_ (.B2(_05221_),
    .C1(_05224_),
    .B1(_05220_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[21] ),
    .Y(_05225_),
    .A2(net9229));
 sg13g2_o21ai_1 _26909_ (.B1(net9417),
    .Y(_05226_),
    .A1(net5248),
    .A2(net7385));
 sg13g2_a21oi_1 _26910_ (.A1(net7385),
    .A2(_05225_),
    .Y(_01223_),
    .B1(_05226_));
 sg13g2_nor2_1 _26911_ (.A(_11335_),
    .B(_05218_),
    .Y(_05227_));
 sg13g2_xnor2_1 _26912_ (.Y(_05228_),
    .A(net8287),
    .B(_05218_));
 sg13g2_nor2_1 _26913_ (.A(net8287),
    .B(net7989),
    .Y(_05229_));
 sg13g2_a21oi_1 _26914_ (.A1(net7987),
    .A2(_05228_),
    .Y(_05230_),
    .B1(_05229_));
 sg13g2_nor2_1 _26915_ (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[23] ),
    .B(_05222_),
    .Y(_05231_));
 sg13g2_a21oi_1 _26916_ (.A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[23] ),
    .A2(_05222_),
    .Y(_05232_),
    .B1(net9063));
 sg13g2_nor2b_1 _26917_ (.A(_05231_),
    .B_N(_05232_),
    .Y(_05233_));
 sg13g2_a221oi_1 _26918_ (.B2(_05230_),
    .C1(_05233_),
    .B1(net8943),
    .A1(net5248),
    .Y(_05234_),
    .A2(net9229));
 sg13g2_o21ai_1 _26919_ (.B1(net9417),
    .Y(_05235_),
    .A1(net5400),
    .A2(net7383));
 sg13g2_a21oi_1 _26920_ (.A1(net7383),
    .A2(_05234_),
    .Y(_01224_),
    .B1(_05235_));
 sg13g2_xnor2_1 _26921_ (.Y(_05236_),
    .A(net8272),
    .B(_05227_));
 sg13g2_nand2_1 _26922_ (.Y(_05237_),
    .A(net8272),
    .B(net7981));
 sg13g2_a21oi_1 _26923_ (.A1(net7989),
    .A2(_05236_),
    .Y(_05238_),
    .B1(_05026_));
 sg13g2_nor3_2 _26924_ (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[24] ),
    .B(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[23] ),
    .C(_05222_),
    .Y(_05239_));
 sg13g2_nor2b_1 _26925_ (.A(_05231_),
    .B_N(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[24] ),
    .Y(_05240_));
 sg13g2_nor3_1 _26926_ (.A(net9063),
    .B(_05239_),
    .C(_05240_),
    .Y(_05241_));
 sg13g2_a221oi_1 _26927_ (.B2(_05238_),
    .C1(_05241_),
    .B1(_05237_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[23] ),
    .Y(_05242_),
    .A2(net9229));
 sg13g2_o21ai_1 _26928_ (.B1(net9417),
    .Y(_05243_),
    .A1(net5373),
    .A2(net7383));
 sg13g2_a21oi_1 _26929_ (.A1(net7383),
    .A2(_05242_),
    .Y(_01225_),
    .B1(_05243_));
 sg13g2_nand3_1 _26930_ (.B(net8270),
    .C(_05227_),
    .A(net8271),
    .Y(_05244_));
 sg13g2_a21o_1 _26931_ (.A2(_05227_),
    .A1(net8271),
    .B1(net8270),
    .X(_05245_));
 sg13g2_nand2_1 _26932_ (.Y(_05246_),
    .A(_05244_),
    .B(_05245_));
 sg13g2_nand2_1 _26933_ (.Y(_05247_),
    .A(net8270),
    .B(net7980));
 sg13g2_a21oi_1 _26934_ (.A1(net7989),
    .A2(_05246_),
    .Y(_05248_),
    .B1(net8939));
 sg13g2_nand2b_2 _26935_ (.Y(_05249_),
    .B(_05239_),
    .A_N(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[25] ));
 sg13g2_nand2b_1 _26936_ (.Y(_05250_),
    .B(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[25] ),
    .A_N(_05239_));
 sg13g2_and3_1 _26937_ (.X(_05251_),
    .A(net9238),
    .B(_05249_),
    .C(_05250_));
 sg13g2_a221oi_1 _26938_ (.B2(_05248_),
    .C1(_05251_),
    .B1(_05247_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[24] ),
    .Y(_05252_),
    .A2(net9229));
 sg13g2_o21ai_1 _26939_ (.B1(net9412),
    .Y(_05253_),
    .A1(net5315),
    .A2(net7383));
 sg13g2_a21oi_1 _26940_ (.A1(net7383),
    .A2(_05252_),
    .Y(_01226_),
    .B1(_05253_));
 sg13g2_nor2_1 _26941_ (.A(_11440_),
    .B(_05244_),
    .Y(_05254_));
 sg13g2_xnor2_1 _26942_ (.Y(_05255_),
    .A(net8275),
    .B(_05244_));
 sg13g2_nor2_1 _26943_ (.A(net7980),
    .B(_05255_),
    .Y(_05256_));
 sg13g2_a21oi_1 _26944_ (.A1(net8275),
    .A2(net7980),
    .Y(_05257_),
    .B1(_05256_));
 sg13g2_o21ai_1 _26945_ (.B1(net9237),
    .Y(_05258_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[26] ),
    .A2(_05249_));
 sg13g2_a21oi_1 _26946_ (.A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[26] ),
    .A2(_05249_),
    .Y(_05259_),
    .B1(_05258_));
 sg13g2_a221oi_1 _26947_ (.B2(_05257_),
    .C1(_05259_),
    .B1(net8943),
    .A1(net5315),
    .Y(_05260_),
    .A2(net9227));
 sg13g2_o21ai_1 _26948_ (.B1(net9412),
    .Y(_05261_),
    .A1(net5504),
    .A2(net7381));
 sg13g2_a21oi_1 _26949_ (.A1(net7381),
    .A2(_05260_),
    .Y(_01227_),
    .B1(_05261_));
 sg13g2_nor3_2 _26950_ (.A(_11440_),
    .B(net8273),
    .C(_05244_),
    .Y(_05262_));
 sg13g2_xor2_1 _26951_ (.B(_05254_),
    .A(net8274),
    .X(_05263_));
 sg13g2_o21ai_1 _26952_ (.B1(net8943),
    .Y(_05264_),
    .A1(net8273),
    .A2(net7989));
 sg13g2_a21oi_1 _26953_ (.A1(net7989),
    .A2(_05263_),
    .Y(_05265_),
    .B1(_05264_));
 sg13g2_nor3_2 _26954_ (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[27] ),
    .B(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[26] ),
    .C(_05249_),
    .Y(_05266_));
 sg13g2_o21ai_1 _26955_ (.B1(net5245),
    .Y(_05267_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[26] ),
    .A2(_05249_));
 sg13g2_nor2_1 _26956_ (.A(net9063),
    .B(_05266_),
    .Y(_05268_));
 sg13g2_a221oi_1 _26957_ (.B2(_05268_),
    .C1(_05265_),
    .B1(_05267_),
    .A1(net5566),
    .Y(_05269_),
    .A2(net9227));
 sg13g2_o21ai_1 _26958_ (.B1(net9412),
    .Y(_05270_),
    .A1(net5245),
    .A2(net7381));
 sg13g2_a21oi_1 _26959_ (.A1(net7381),
    .A2(_05269_),
    .Y(_01228_),
    .B1(_05270_));
 sg13g2_nand2_1 _26960_ (.Y(_05271_),
    .A(net8268),
    .B(_05262_));
 sg13g2_xnor2_1 _26961_ (.Y(_05272_),
    .A(net8268),
    .B(_05262_));
 sg13g2_nand2_1 _26962_ (.Y(_05273_),
    .A(net8268),
    .B(net7980));
 sg13g2_a21oi_1 _26963_ (.A1(net7989),
    .A2(_05272_),
    .Y(_05274_),
    .B1(net8939));
 sg13g2_nand2b_2 _26964_ (.Y(_05275_),
    .B(_05266_),
    .A_N(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[28] ));
 sg13g2_nand2b_1 _26965_ (.Y(_05276_),
    .B(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[28] ),
    .A_N(_05266_));
 sg13g2_and3_1 _26966_ (.X(_05277_),
    .A(net9237),
    .B(_05275_),
    .C(_05276_));
 sg13g2_a221oi_1 _26967_ (.B2(_05274_),
    .C1(_05277_),
    .B1(_05273_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[27] ),
    .Y(_05278_),
    .A2(net9227));
 sg13g2_o21ai_1 _26968_ (.B1(net9412),
    .Y(_05279_),
    .A1(net5222),
    .A2(net7381));
 sg13g2_a21oi_1 _26969_ (.A1(net7381),
    .A2(_05278_),
    .Y(_01229_),
    .B1(_05279_));
 sg13g2_nand3_1 _26970_ (.B(net8268),
    .C(_05262_),
    .A(net8307),
    .Y(_05280_));
 sg13g2_xnor2_1 _26971_ (.Y(_05281_),
    .A(net8307),
    .B(_05271_));
 sg13g2_nor2_1 _26972_ (.A(net7981),
    .B(_05281_),
    .Y(_05282_));
 sg13g2_a21oi_1 _26973_ (.A1(net8308),
    .A2(net7980),
    .Y(_05283_),
    .B1(_05282_));
 sg13g2_o21ai_1 _26974_ (.B1(net9237),
    .Y(_05284_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[29] ),
    .A2(_05275_));
 sg13g2_a21oi_1 _26975_ (.A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[29] ),
    .A2(_05275_),
    .Y(_05285_),
    .B1(_05284_));
 sg13g2_a221oi_1 _26976_ (.B2(_05283_),
    .C1(_05285_),
    .B1(net8943),
    .A1(net5222),
    .Y(_05286_),
    .A2(net9227));
 sg13g2_o21ai_1 _26977_ (.B1(net9412),
    .Y(_05287_),
    .A1(net5409),
    .A2(net7381));
 sg13g2_a21oi_1 _26978_ (.A1(net7381),
    .A2(_05286_),
    .Y(_01230_),
    .B1(_05287_));
 sg13g2_nor2_1 _26979_ (.A(_11053_),
    .B(_05280_),
    .Y(_05288_));
 sg13g2_xnor2_1 _26980_ (.Y(_05289_),
    .A(_11052_),
    .B(_05280_));
 sg13g2_o21ai_1 _26981_ (.B1(net8943),
    .Y(_05290_),
    .A1(net7980),
    .A2(_05289_));
 sg13g2_a21oi_1 _26982_ (.A1(_11052_),
    .A2(net7980),
    .Y(_05291_),
    .B1(_05290_));
 sg13g2_nor3_1 _26983_ (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[30] ),
    .B(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[29] ),
    .C(_05275_),
    .Y(_05292_));
 sg13g2_o21ai_1 _26984_ (.B1(net5261),
    .Y(_05293_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[29] ),
    .A2(_05275_));
 sg13g2_nor2_1 _26985_ (.A(net9063),
    .B(_05292_),
    .Y(_05294_));
 sg13g2_a221oi_1 _26986_ (.B2(_05294_),
    .C1(_05291_),
    .B1(_05293_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[29] ),
    .Y(_05295_),
    .A2(net9227));
 sg13g2_o21ai_1 _26987_ (.B1(net9412),
    .Y(_05296_),
    .A1(net5261),
    .A2(net7382));
 sg13g2_a21oi_1 _26988_ (.A1(net7382),
    .A2(_05295_),
    .Y(_01231_),
    .B1(_05296_));
 sg13g2_nor2_1 _26989_ (.A(_04807_),
    .B(_05288_),
    .Y(_05297_));
 sg13g2_nor3_1 _26990_ (.A(net8314),
    .B(net8939),
    .C(_05297_),
    .Y(_05298_));
 sg13g2_xnor2_1 _26991_ (.Y(_05299_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[31] ),
    .B(_05292_));
 sg13g2_a221oi_1 _26992_ (.B2(net9237),
    .C1(_05298_),
    .B1(_05299_),
    .A1(net5261),
    .Y(_05300_),
    .A2(net9227));
 sg13g2_o21ai_1 _26993_ (.B1(net9412),
    .Y(_05301_),
    .A1(net5477),
    .A2(net7382));
 sg13g2_a21oi_1 _26994_ (.A1(net7382),
    .A2(_05300_),
    .Y(_01232_),
    .B1(_05301_));
 sg13g2_a21o_2 _26995_ (.A2(net7980),
    .A1(net9237),
    .B1(_05028_),
    .X(_05302_));
 sg13g2_nor2_1 _26996_ (.A(net8943),
    .B(net7879),
    .Y(_05303_));
 sg13g2_a21o_1 _26997_ (.A2(_05020_),
    .A1(net8516),
    .B1(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[31] ),
    .X(_05304_));
 sg13g2_nand3_1 _26998_ (.B(net8516),
    .C(_05020_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[31] ),
    .Y(_05305_));
 sg13g2_nand3_1 _26999_ (.B(_05304_),
    .C(_05305_),
    .A(net9230),
    .Y(_05306_));
 sg13g2_o21ai_1 _27000_ (.B1(_05306_),
    .Y(_05307_),
    .A1(net9063),
    .A2(_10517_));
 sg13g2_a22oi_1 _27001_ (.Y(_05308_),
    .B1(net7757),
    .B2(_05307_),
    .A2(net7879),
    .A1(net4684));
 sg13g2_nor2_1 _27002_ (.A(net9056),
    .B(_05308_),
    .Y(_01233_));
 sg13g2_xnor2_1 _27003_ (.Y(_05309_),
    .A(_04893_),
    .B(_04895_));
 sg13g2_nand2_1 _27004_ (.Y(_05310_),
    .A(_10516_),
    .B(_10517_));
 sg13g2_a21oi_1 _27005_ (.A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[1] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[0] ),
    .Y(_05311_),
    .B1(net9232));
 sg13g2_nor2b_1 _27006_ (.A(_05020_),
    .B_N(net9229),
    .Y(_05312_));
 sg13g2_inv_2 _27007_ (.Y(_05313_),
    .A(net7328));
 sg13g2_a22oi_1 _27008_ (.Y(_05314_),
    .B1(net7329),
    .B2(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[0] ),
    .A2(_05311_),
    .A1(_05310_));
 sg13g2_o21ai_1 _27009_ (.B1(_05314_),
    .Y(_05315_),
    .A1(net7330),
    .A2(_05309_));
 sg13g2_a22oi_1 _27010_ (.Y(_05316_),
    .B1(net7757),
    .B2(_05315_),
    .A2(net7879),
    .A1(net4362));
 sg13g2_nor2_1 _27011_ (.A(net9056),
    .B(net4363),
    .Y(_01234_));
 sg13g2_o21ai_1 _27012_ (.B1(_04896_),
    .Y(_05317_),
    .A1(_04897_),
    .A2(_04898_));
 sg13g2_nand2b_1 _27013_ (.Y(_05318_),
    .B(_05317_),
    .A_N(_04899_));
 sg13g2_or2_1 _27014_ (.X(_05319_),
    .B(_05310_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[2] ));
 sg13g2_a21oi_1 _27015_ (.A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[2] ),
    .A2(_05310_),
    .Y(_05320_),
    .B1(net9232));
 sg13g2_a22oi_1 _27016_ (.Y(_05321_),
    .B1(_05319_),
    .B2(_05320_),
    .A2(net7329),
    .A1(_10831_));
 sg13g2_o21ai_1 _27017_ (.B1(_05321_),
    .Y(_05322_),
    .A1(net7330),
    .A2(_05318_));
 sg13g2_a22oi_1 _27018_ (.Y(_05323_),
    .B1(net7759),
    .B2(_05322_),
    .A2(net7881),
    .A1(net5239));
 sg13g2_nor2_1 _27019_ (.A(net9056),
    .B(net5240),
    .Y(_01235_));
 sg13g2_xor2_1 _27020_ (.B(_04901_),
    .A(_04900_),
    .X(_05324_));
 sg13g2_or2_1 _27021_ (.X(_05325_),
    .B(_05319_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[3] ));
 sg13g2_a21oi_1 _27022_ (.A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[3] ),
    .A2(_05319_),
    .Y(_05326_),
    .B1(net9234));
 sg13g2_a22oi_1 _27023_ (.Y(_05327_),
    .B1(_05325_),
    .B2(_05326_),
    .A2(net7329),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[2] ));
 sg13g2_o21ai_1 _27024_ (.B1(_05327_),
    .Y(_05328_),
    .A1(net7330),
    .A2(_05324_));
 sg13g2_a22oi_1 _27025_ (.Y(_05329_),
    .B1(net7759),
    .B2(_05328_),
    .A2(net7881),
    .A1(net5154));
 sg13g2_nor2_1 _27026_ (.A(net9056),
    .B(net5155),
    .Y(_01236_));
 sg13g2_nand3_1 _27027_ (.B(_04902_),
    .C(_04903_),
    .A(_04884_),
    .Y(_05330_));
 sg13g2_nand2b_1 _27028_ (.Y(_05331_),
    .B(_05330_),
    .A_N(_04904_));
 sg13g2_nand2_1 _27029_ (.Y(_05332_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[4] ),
    .B(_05325_));
 sg13g2_or2_1 _27030_ (.X(_05333_),
    .B(_05325_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[4] ));
 sg13g2_nor2b_1 _27031_ (.A(net9234),
    .B_N(_05333_),
    .Y(_05334_));
 sg13g2_a22oi_1 _27032_ (.Y(_05335_),
    .B1(_05332_),
    .B2(_05334_),
    .A2(net7327),
    .A1(_10830_));
 sg13g2_o21ai_1 _27033_ (.B1(_05335_),
    .Y(_05336_),
    .A1(_05022_),
    .A2(_05331_));
 sg13g2_a22oi_1 _27034_ (.Y(_05337_),
    .B1(net7759),
    .B2(_05336_),
    .A2(net7881),
    .A1(net5052));
 sg13g2_nor2_1 _27035_ (.A(net9056),
    .B(net5053),
    .Y(_01237_));
 sg13g2_or3_1 _27036_ (.A(_04881_),
    .B(_04904_),
    .C(_04905_),
    .X(_05338_));
 sg13g2_nand2_1 _27037_ (.Y(_05339_),
    .A(_04906_),
    .B(_05338_));
 sg13g2_nand2_1 _27038_ (.Y(_05340_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[5] ),
    .B(_05333_));
 sg13g2_nor2_1 _27039_ (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[5] ),
    .B(_05333_),
    .Y(_05341_));
 sg13g2_nor2_1 _27040_ (.A(net9234),
    .B(_05341_),
    .Y(_05342_));
 sg13g2_a22oi_1 _27041_ (.Y(_05343_),
    .B1(_05340_),
    .B2(_05342_),
    .A2(net7327),
    .A1(_10829_));
 sg13g2_o21ai_1 _27042_ (.B1(_05343_),
    .Y(_05344_),
    .A1(net7330),
    .A2(_05339_));
 sg13g2_a22oi_1 _27043_ (.Y(_05345_),
    .B1(net7759),
    .B2(_05344_),
    .A2(net7881),
    .A1(net5280));
 sg13g2_nor2_1 _27044_ (.A(net9057),
    .B(net5281),
    .Y(_01238_));
 sg13g2_nand3_1 _27045_ (.B(_04906_),
    .C(_04907_),
    .A(_04878_),
    .Y(_05346_));
 sg13g2_nor2b_1 _27046_ (.A(_04908_),
    .B_N(_05346_),
    .Y(_05347_));
 sg13g2_nor3_2 _27047_ (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[6] ),
    .B(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[5] ),
    .C(_05333_),
    .Y(_05348_));
 sg13g2_xor2_1 _27048_ (.B(_05341_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[6] ),
    .X(_05349_));
 sg13g2_a22oi_1 _27049_ (.Y(_05350_),
    .B1(_05347_),
    .B2(net7331),
    .A2(net7327),
    .A1(_10828_));
 sg13g2_o21ai_1 _27050_ (.B1(_05350_),
    .Y(_05351_),
    .A1(net9233),
    .A2(_05349_));
 sg13g2_a22oi_1 _27051_ (.Y(_05352_),
    .B1(net7758),
    .B2(_05351_),
    .A2(net7880),
    .A1(net5376));
 sg13g2_nor2_1 _27052_ (.A(net9057),
    .B(net5377),
    .Y(_01239_));
 sg13g2_or3_1 _27053_ (.A(_04874_),
    .B(_04908_),
    .C(_04909_),
    .X(_05353_));
 sg13g2_and2_1 _27054_ (.A(_04910_),
    .B(_05353_),
    .X(_05354_));
 sg13g2_nand2_2 _27055_ (.Y(_05355_),
    .A(_10515_),
    .B(_05348_));
 sg13g2_xnor2_1 _27056_ (.Y(_05356_),
    .A(_10515_),
    .B(_05348_));
 sg13g2_a22oi_1 _27057_ (.Y(_05357_),
    .B1(_05354_),
    .B2(net7331),
    .A2(net7327),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[6] ));
 sg13g2_o21ai_1 _27058_ (.B1(_05357_),
    .Y(_05358_),
    .A1(net9233),
    .A2(_05356_));
 sg13g2_a22oi_1 _27059_ (.Y(_05359_),
    .B1(net7758),
    .B2(_05358_),
    .A2(net7880),
    .A1(net3964));
 sg13g2_nor2_1 _27060_ (.A(net9057),
    .B(_05359_),
    .Y(_01240_));
 sg13g2_nand3_1 _27061_ (.B(_04910_),
    .C(_04914_),
    .A(_04870_),
    .Y(_05360_));
 sg13g2_and2_1 _27062_ (.A(_04915_),
    .B(_05360_),
    .X(_05361_));
 sg13g2_xnor2_1 _27063_ (.Y(_05362_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[8] ),
    .B(_05355_));
 sg13g2_a22oi_1 _27064_ (.Y(_05363_),
    .B1(_05361_),
    .B2(net7331),
    .A2(net7327),
    .A1(_10827_));
 sg13g2_o21ai_1 _27065_ (.B1(_05363_),
    .Y(_05364_),
    .A1(net9233),
    .A2(_05362_));
 sg13g2_a22oi_1 _27066_ (.Y(_05365_),
    .B1(net7758),
    .B2(net5362),
    .A2(net7880),
    .A1(net5310));
 sg13g2_nor2_1 _27067_ (.A(net9057),
    .B(_05365_),
    .Y(_01241_));
 sg13g2_nand3_1 _27068_ (.B(_04916_),
    .C(_04920_),
    .A(_04915_),
    .Y(_05366_));
 sg13g2_nor2b_1 _27069_ (.A(_04921_),
    .B_N(_05366_),
    .Y(_05367_));
 sg13g2_o21ai_1 _27070_ (.B1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[9] ),
    .Y(_05368_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[8] ),
    .A2(_05355_));
 sg13g2_nor3_2 _27071_ (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[9] ),
    .B(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[8] ),
    .C(_05355_),
    .Y(_05369_));
 sg13g2_nor2_1 _27072_ (.A(net9233),
    .B(_05369_),
    .Y(_05370_));
 sg13g2_a22oi_1 _27073_ (.Y(_05371_),
    .B1(_05368_),
    .B2(_05370_),
    .A2(_05367_),
    .A1(net7331));
 sg13g2_o21ai_1 _27074_ (.B1(_05371_),
    .Y(_05372_),
    .A1(net4080),
    .A2(net7326));
 sg13g2_a22oi_1 _27075_ (.Y(_05373_),
    .B1(net7758),
    .B2(_05372_),
    .A2(net7880),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[9] ));
 sg13g2_nor2_1 _27076_ (.A(net9057),
    .B(net4081),
    .Y(_01242_));
 sg13g2_xnor2_1 _27077_ (.Y(_05374_),
    .A(_04922_),
    .B(_04926_));
 sg13g2_nand2b_2 _27078_ (.Y(_05375_),
    .B(_05369_),
    .A_N(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[10] ));
 sg13g2_xor2_1 _27079_ (.B(_05369_),
    .A(net5020),
    .X(_05376_));
 sg13g2_a22oi_1 _27080_ (.Y(_05377_),
    .B1(_05374_),
    .B2(net7331),
    .A2(net7327),
    .A1(_10826_));
 sg13g2_o21ai_1 _27081_ (.B1(_05377_),
    .Y(_05378_),
    .A1(net9233),
    .A2(_05376_));
 sg13g2_a22oi_1 _27082_ (.Y(_05379_),
    .B1(net7758),
    .B2(_05378_),
    .A2(net7880),
    .A1(net5020));
 sg13g2_nor2_1 _27083_ (.A(net9057),
    .B(net5021),
    .Y(_01243_));
 sg13g2_nand3_1 _27084_ (.B(_04928_),
    .C(_04932_),
    .A(_04927_),
    .Y(_05380_));
 sg13g2_and2_1 _27085_ (.A(net7331),
    .B(_05380_),
    .X(_05381_));
 sg13g2_xnor2_1 _27086_ (.Y(_05382_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[11] ),
    .B(_05375_));
 sg13g2_a22oi_1 _27087_ (.Y(_05383_),
    .B1(_05381_),
    .B2(_04933_),
    .A2(net7328),
    .A1(_10825_));
 sg13g2_o21ai_1 _27088_ (.B1(_05383_),
    .Y(_05384_),
    .A1(net9233),
    .A2(_05382_));
 sg13g2_a22oi_1 _27089_ (.Y(_05385_),
    .B1(net7758),
    .B2(_05384_),
    .A2(net7880),
    .A1(net5332));
 sg13g2_nor2_1 _27090_ (.A(net9057),
    .B(net5333),
    .Y(_01244_));
 sg13g2_nand3_1 _27091_ (.B(_04934_),
    .C(_04939_),
    .A(_04933_),
    .Y(_05386_));
 sg13g2_nor2b_1 _27092_ (.A(_04940_),
    .B_N(_05386_),
    .Y(_05387_));
 sg13g2_o21ai_1 _27093_ (.B1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[12] ),
    .Y(_05388_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[11] ),
    .A2(_05375_));
 sg13g2_nor3_2 _27094_ (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[12] ),
    .B(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[11] ),
    .C(_05375_),
    .Y(_05389_));
 sg13g2_nor2_1 _27095_ (.A(net9233),
    .B(_05389_),
    .Y(_05390_));
 sg13g2_a22oi_1 _27096_ (.Y(_05391_),
    .B1(_05388_),
    .B2(_05390_),
    .A2(_05387_),
    .A1(net7331));
 sg13g2_o21ai_1 _27097_ (.B1(_05391_),
    .Y(_05392_),
    .A1(net4802),
    .A2(net7326));
 sg13g2_a22oi_1 _27098_ (.Y(_05393_),
    .B1(net7758),
    .B2(_05392_),
    .A2(net7880),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[12] ));
 sg13g2_nor2_1 _27099_ (.A(net9057),
    .B(net4803),
    .Y(_01245_));
 sg13g2_xor2_1 _27100_ (.B(_04945_),
    .A(_04941_),
    .X(_05394_));
 sg13g2_nand2b_2 _27101_ (.Y(_05395_),
    .B(_05389_),
    .A_N(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[13] ));
 sg13g2_xor2_1 _27102_ (.B(_05389_),
    .A(net4914),
    .X(_05396_));
 sg13g2_a22oi_1 _27103_ (.Y(_05397_),
    .B1(_05394_),
    .B2(net7331),
    .A2(net7328),
    .A1(_10824_));
 sg13g2_o21ai_1 _27104_ (.B1(_05397_),
    .Y(_05398_),
    .A1(net9233),
    .A2(_05396_));
 sg13g2_a22oi_1 _27105_ (.Y(_05399_),
    .B1(net7758),
    .B2(_05398_),
    .A2(net7880),
    .A1(net4914));
 sg13g2_nor2_1 _27106_ (.A(net9058),
    .B(net4915),
    .Y(_01246_));
 sg13g2_xnor2_1 _27107_ (.Y(_05400_),
    .A(_04946_),
    .B(_04950_));
 sg13g2_nand2_1 _27108_ (.Y(_05401_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[14] ),
    .B(_05395_));
 sg13g2_nor2_1 _27109_ (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[14] ),
    .B(_05395_),
    .Y(_05402_));
 sg13g2_nor2_1 _27110_ (.A(net9234),
    .B(_05402_),
    .Y(_05403_));
 sg13g2_a22oi_1 _27111_ (.Y(_05404_),
    .B1(_05401_),
    .B2(_05403_),
    .A2(net7327),
    .A1(_10823_));
 sg13g2_o21ai_1 _27112_ (.B1(_05404_),
    .Y(_05405_),
    .A1(net7330),
    .A2(_05400_));
 sg13g2_a22oi_1 _27113_ (.Y(_05406_),
    .B1(net7759),
    .B2(_05405_),
    .A2(net7881),
    .A1(net5337));
 sg13g2_nor2_1 _27114_ (.A(net9058),
    .B(net5338),
    .Y(_01247_));
 sg13g2_xnor2_1 _27115_ (.Y(_05407_),
    .A(_04952_),
    .B(_04953_));
 sg13g2_nor3_2 _27116_ (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[15] ),
    .B(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[14] ),
    .C(_05395_),
    .Y(_05408_));
 sg13g2_xor2_1 _27117_ (.B(_05402_),
    .A(net4937),
    .X(_05409_));
 sg13g2_a22oi_1 _27118_ (.Y(_05410_),
    .B1(_05407_),
    .B2(net7332),
    .A2(net7327),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[14] ));
 sg13g2_o21ai_1 _27119_ (.B1(_05410_),
    .Y(_05411_),
    .A1(net9234),
    .A2(_05409_));
 sg13g2_a22oi_1 _27120_ (.Y(_05412_),
    .B1(net7759),
    .B2(_05411_),
    .A2(net7881),
    .A1(net4937));
 sg13g2_nor2_1 _27121_ (.A(net9059),
    .B(_05412_),
    .Y(_01248_));
 sg13g2_or3_1 _27122_ (.A(_04866_),
    .B(_04954_),
    .C(_04958_),
    .X(_05413_));
 sg13g2_and2_1 _27123_ (.A(_04959_),
    .B(_05413_),
    .X(_05414_));
 sg13g2_nand2b_2 _27124_ (.Y(_05415_),
    .B(_05408_),
    .A_N(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[16] ));
 sg13g2_xor2_1 _27125_ (.B(_05408_),
    .A(net4911),
    .X(_05416_));
 sg13g2_a22oi_1 _27126_ (.Y(_05417_),
    .B1(_05414_),
    .B2(net7332),
    .A2(net7328),
    .A1(_10822_));
 sg13g2_o21ai_1 _27127_ (.B1(_05417_),
    .Y(_05418_),
    .A1(net9236),
    .A2(_05416_));
 sg13g2_a22oi_1 _27128_ (.Y(_05419_),
    .B1(net7761),
    .B2(_05418_),
    .A2(_05302_),
    .A1(net4911));
 sg13g2_nor2_1 _27129_ (.A(net9058),
    .B(net4912),
    .Y(_01249_));
 sg13g2_nand3_1 _27130_ (.B(_04960_),
    .C(_04965_),
    .A(_04959_),
    .Y(_05420_));
 sg13g2_nor2b_1 _27131_ (.A(_04966_),
    .B_N(_05420_),
    .Y(_05421_));
 sg13g2_xnor2_1 _27132_ (.Y(_05422_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[17] ),
    .B(_05415_));
 sg13g2_a22oi_1 _27133_ (.Y(_05423_),
    .B1(_05421_),
    .B2(net7332),
    .A2(net7328),
    .A1(_10821_));
 sg13g2_o21ai_1 _27134_ (.B1(_05423_),
    .Y(_05424_),
    .A1(net9235),
    .A2(_05422_));
 sg13g2_a22oi_1 _27135_ (.Y(_05425_),
    .B1(net7760),
    .B2(_05424_),
    .A2(net7882),
    .A1(net5138));
 sg13g2_nor2_1 _27136_ (.A(net9058),
    .B(net5139),
    .Y(_01250_));
 sg13g2_xor2_1 _27137_ (.B(_04971_),
    .A(_04967_),
    .X(_05426_));
 sg13g2_o21ai_1 _27138_ (.B1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[18] ),
    .Y(_05427_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[17] ),
    .A2(_05415_));
 sg13g2_nor3_2 _27139_ (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[18] ),
    .B(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[17] ),
    .C(_05415_),
    .Y(_05428_));
 sg13g2_nor2_1 _27140_ (.A(net9235),
    .B(_05428_),
    .Y(_05429_));
 sg13g2_a22oi_1 _27141_ (.Y(_05430_),
    .B1(_05427_),
    .B2(_05429_),
    .A2(net7329),
    .A1(_10820_));
 sg13g2_o21ai_1 _27142_ (.B1(_05430_),
    .Y(_05431_),
    .A1(net7330),
    .A2(_05426_));
 sg13g2_a22oi_1 _27143_ (.Y(_05432_),
    .B1(net7760),
    .B2(_05431_),
    .A2(net7882),
    .A1(net4999));
 sg13g2_nor2_1 _27144_ (.A(net9059),
    .B(net5000),
    .Y(_01251_));
 sg13g2_xor2_1 _27145_ (.B(_04977_),
    .A(_04973_),
    .X(_05433_));
 sg13g2_nand2b_2 _27146_ (.Y(_05434_),
    .B(_05428_),
    .A_N(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[19] ));
 sg13g2_xor2_1 _27147_ (.B(_05428_),
    .A(net5057),
    .X(_05435_));
 sg13g2_a22oi_1 _27148_ (.Y(_05436_),
    .B1(_05433_),
    .B2(net7332),
    .A2(net7328),
    .A1(_10819_));
 sg13g2_o21ai_1 _27149_ (.B1(_05436_),
    .Y(_05437_),
    .A1(net9235),
    .A2(_05435_));
 sg13g2_a22oi_1 _27150_ (.Y(_05438_),
    .B1(net7760),
    .B2(_05437_),
    .A2(net7882),
    .A1(net5057));
 sg13g2_nor2_1 _27151_ (.A(net9058),
    .B(net5058),
    .Y(_01252_));
 sg13g2_xnor2_1 _27152_ (.Y(_05439_),
    .A(_04978_),
    .B(_04979_));
 sg13g2_xnor2_1 _27153_ (.Y(_05440_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[20] ),
    .B(_05434_));
 sg13g2_a22oi_1 _27154_ (.Y(_05441_),
    .B1(_05439_),
    .B2(net7332),
    .A2(net7328),
    .A1(_10818_));
 sg13g2_o21ai_1 _27155_ (.B1(_05441_),
    .Y(_05442_),
    .A1(net9235),
    .A2(_05440_));
 sg13g2_a22oi_1 _27156_ (.Y(_05443_),
    .B1(net7760),
    .B2(_05442_),
    .A2(net7882),
    .A1(net5171));
 sg13g2_nor2_1 _27157_ (.A(net9058),
    .B(net5172),
    .Y(_01253_));
 sg13g2_xor2_1 _27158_ (.B(_04981_),
    .A(_04859_),
    .X(_05444_));
 sg13g2_nor3_1 _27159_ (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[21] ),
    .B(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[20] ),
    .C(_05434_),
    .Y(_05445_));
 sg13g2_o21ai_1 _27160_ (.B1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[21] ),
    .Y(_05446_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[20] ),
    .A2(_05434_));
 sg13g2_nor2_1 _27161_ (.A(net9235),
    .B(_05445_),
    .Y(_05447_));
 sg13g2_a22oi_1 _27162_ (.Y(_05448_),
    .B1(_05446_),
    .B2(_05447_),
    .A2(_05444_),
    .A1(net7333));
 sg13g2_o21ai_1 _27163_ (.B1(_05448_),
    .Y(_05449_),
    .A1(net4896),
    .A2(_05313_));
 sg13g2_a22oi_1 _27164_ (.Y(_05450_),
    .B1(net7760),
    .B2(_05449_),
    .A2(net7882),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[21] ));
 sg13g2_nor2_1 _27165_ (.A(net9058),
    .B(net4897),
    .Y(_01254_));
 sg13g2_nand3_1 _27166_ (.B(_04982_),
    .C(_04983_),
    .A(_04858_),
    .Y(_05451_));
 sg13g2_and2_1 _27167_ (.A(net7332),
    .B(_05451_),
    .X(_05452_));
 sg13g2_nand2b_1 _27168_ (.Y(_05453_),
    .B(_05445_),
    .A_N(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[22] ));
 sg13g2_nand2b_1 _27169_ (.Y(_05454_),
    .B(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[22] ),
    .A_N(_05445_));
 sg13g2_nand3b_1 _27170_ (.B(_05453_),
    .C(_05454_),
    .Y(_05455_),
    .A_N(net9235));
 sg13g2_o21ai_1 _27171_ (.B1(_05455_),
    .Y(_05456_),
    .A1(_00166_),
    .A2(_05313_));
 sg13g2_a21o_1 _27172_ (.A2(_05452_),
    .A1(_04984_),
    .B1(_05456_),
    .X(_05457_));
 sg13g2_a22oi_1 _27173_ (.Y(_05458_),
    .B1(net7760),
    .B2(_05457_),
    .A2(net7882),
    .A1(net5081));
 sg13g2_nor2_1 _27174_ (.A(net9056),
    .B(net5082),
    .Y(_01255_));
 sg13g2_nand3_1 _27175_ (.B(_04854_),
    .C(_04984_),
    .A(_04850_),
    .Y(_05459_));
 sg13g2_nor2b_1 _27176_ (.A(_04985_),
    .B_N(_05459_),
    .Y(_05460_));
 sg13g2_or2_2 _27177_ (.X(_05461_),
    .B(_05453_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[23] ));
 sg13g2_a21oi_1 _27178_ (.A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[23] ),
    .A2(_05453_),
    .Y(_05462_),
    .B1(net9235));
 sg13g2_a22oi_1 _27179_ (.Y(_05463_),
    .B1(_05461_),
    .B2(_05462_),
    .A2(_05460_),
    .A1(net7332));
 sg13g2_o21ai_1 _27180_ (.B1(_05463_),
    .Y(_05464_),
    .A1(_00165_),
    .A2(_05313_));
 sg13g2_a22oi_1 _27181_ (.Y(_05465_),
    .B1(net7760),
    .B2(_05464_),
    .A2(net7882),
    .A1(net4408));
 sg13g2_nor2_1 _27182_ (.A(net9059),
    .B(net4409),
    .Y(_01256_));
 sg13g2_nand2_1 _27183_ (.Y(_05466_),
    .A(net5186),
    .B(net7878));
 sg13g2_xnor2_1 _27184_ (.Y(_05467_),
    .A(_04986_),
    .B(_04990_));
 sg13g2_nor2_1 _27185_ (.A(_00164_),
    .B(net7326),
    .Y(_05468_));
 sg13g2_a21oi_1 _27186_ (.A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[24] ),
    .A2(_05461_),
    .Y(_05469_),
    .B1(net9232));
 sg13g2_o21ai_1 _27187_ (.B1(_05469_),
    .Y(_05470_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[24] ),
    .A2(_05461_));
 sg13g2_o21ai_1 _27188_ (.B1(_05470_),
    .Y(_05471_),
    .A1(net7330),
    .A2(_05467_));
 sg13g2_o21ai_1 _27189_ (.B1(net7757),
    .Y(_05472_),
    .A1(_05468_),
    .A2(_05471_));
 sg13g2_a21oi_1 _27190_ (.A1(_05466_),
    .A2(_05472_),
    .Y(_01257_),
    .B1(net9059));
 sg13g2_xnor2_1 _27191_ (.Y(_05473_),
    .A(_04991_),
    .B(_04992_));
 sg13g2_o21ai_1 _27192_ (.B1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[25] ),
    .Y(_05474_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[24] ),
    .A2(_05461_));
 sg13g2_or3_2 _27193_ (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[25] ),
    .B(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[24] ),
    .C(_05461_),
    .X(_05475_));
 sg13g2_nor2b_1 _27194_ (.A(net9232),
    .B_N(_05474_),
    .Y(_05476_));
 sg13g2_a22oi_1 _27195_ (.Y(_05477_),
    .B1(_05475_),
    .B2(_05476_),
    .A2(_05473_),
    .A1(net7333));
 sg13g2_o21ai_1 _27196_ (.B1(_05477_),
    .Y(_05478_),
    .A1(_00163_),
    .A2(net7326));
 sg13g2_a22oi_1 _27197_ (.Y(_05479_),
    .B1(net7757),
    .B2(_05478_),
    .A2(net7878),
    .A1(net4768));
 sg13g2_nor2_1 _27198_ (.A(net9056),
    .B(net4769),
    .Y(_01258_));
 sg13g2_xor2_1 _27199_ (.B(_04998_),
    .A(_04994_),
    .X(_05480_));
 sg13g2_nand2_1 _27200_ (.Y(_05481_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[26] ),
    .B(_05475_));
 sg13g2_nor2_1 _27201_ (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[26] ),
    .B(_05475_),
    .Y(_05482_));
 sg13g2_nor2_1 _27202_ (.A(net9232),
    .B(_05482_),
    .Y(_05483_));
 sg13g2_a22oi_1 _27203_ (.Y(_05484_),
    .B1(_05481_),
    .B2(_05483_),
    .A2(_05480_),
    .A1(net7333));
 sg13g2_o21ai_1 _27204_ (.B1(_05484_),
    .Y(_05485_),
    .A1(net4821),
    .A2(net7326));
 sg13g2_a22oi_1 _27205_ (.Y(_05486_),
    .B1(net7757),
    .B2(_05485_),
    .A2(net7878),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[26] ));
 sg13g2_nor2_1 _27206_ (.A(net9056),
    .B(net4822),
    .Y(_01259_));
 sg13g2_xnor2_1 _27207_ (.Y(_05487_),
    .A(_04999_),
    .B(_05000_));
 sg13g2_nor2b_1 _27208_ (.A(_05482_),
    .B_N(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[27] ),
    .Y(_05488_));
 sg13g2_nor3_2 _27209_ (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[27] ),
    .B(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[26] ),
    .C(_05475_),
    .Y(_05489_));
 sg13g2_inv_1 _27210_ (.Y(_05490_),
    .A(_05489_));
 sg13g2_nor2_1 _27211_ (.A(net9232),
    .B(_05488_),
    .Y(_05491_));
 sg13g2_a22oi_1 _27212_ (.Y(_05492_),
    .B1(_05490_),
    .B2(_05491_),
    .A2(_05487_),
    .A1(net7333));
 sg13g2_o21ai_1 _27213_ (.B1(_05492_),
    .Y(_05493_),
    .A1(net5022),
    .A2(net7326));
 sg13g2_a22oi_1 _27214_ (.Y(_05494_),
    .B1(net7757),
    .B2(_05493_),
    .A2(net7878),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[27] ));
 sg13g2_nor2_1 _27215_ (.A(net9054),
    .B(net5023),
    .Y(_01260_));
 sg13g2_nand2b_2 _27216_ (.Y(_05495_),
    .B(_05489_),
    .A_N(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[28] ));
 sg13g2_a21oi_1 _27217_ (.A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[28] ),
    .A2(_05490_),
    .Y(_05496_),
    .B1(net9232));
 sg13g2_xor2_1 _27218_ (.B(_05006_),
    .A(_05002_),
    .X(_05497_));
 sg13g2_a22oi_1 _27219_ (.Y(_05498_),
    .B1(_05497_),
    .B2(net7333),
    .A2(_05496_),
    .A1(_05495_));
 sg13g2_o21ai_1 _27220_ (.B1(_05498_),
    .Y(_05499_),
    .A1(_00160_),
    .A2(net7326));
 sg13g2_a22oi_1 _27221_ (.Y(_05500_),
    .B1(net7761),
    .B2(_05499_),
    .A2(net7878),
    .A1(net4872));
 sg13g2_nor2_1 _27222_ (.A(net9054),
    .B(net4873),
    .Y(_01261_));
 sg13g2_nand3_1 _27223_ (.B(_05008_),
    .C(_05009_),
    .A(_05007_),
    .Y(_05501_));
 sg13g2_nor2b_1 _27224_ (.A(_05010_),
    .B_N(_05501_),
    .Y(_05502_));
 sg13g2_nand2b_1 _27225_ (.Y(_05503_),
    .B(net7329),
    .A_N(_00159_));
 sg13g2_xnor2_1 _27226_ (.Y(_05504_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[29] ),
    .B(_05495_));
 sg13g2_o21ai_1 _27227_ (.B1(_05503_),
    .Y(_05505_),
    .A1(net9232),
    .A2(_05504_));
 sg13g2_a21o_1 _27228_ (.A2(_05502_),
    .A1(net7333),
    .B1(_05505_),
    .X(_05506_));
 sg13g2_a22oi_1 _27229_ (.Y(_05507_),
    .B1(net7757),
    .B2(_05506_),
    .A2(net7878),
    .A1(net5217));
 sg13g2_nor2_1 _27230_ (.A(net9055),
    .B(_05507_),
    .Y(_01262_));
 sg13g2_xor2_1 _27231_ (.B(_05015_),
    .A(_05011_),
    .X(_05508_));
 sg13g2_nor3_1 _27232_ (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[30] ),
    .B(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[29] ),
    .C(_05495_),
    .Y(_05509_));
 sg13g2_o21ai_1 _27233_ (.B1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[30] ),
    .Y(_05510_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[29] ),
    .A2(_05495_));
 sg13g2_nor2_1 _27234_ (.A(net9236),
    .B(_05509_),
    .Y(_05511_));
 sg13g2_a22oi_1 _27235_ (.Y(_05512_),
    .B1(_05510_),
    .B2(_05511_),
    .A2(_05508_),
    .A1(net7333));
 sg13g2_o21ai_1 _27236_ (.B1(_05512_),
    .Y(_05513_),
    .A1(net4917),
    .A2(net7326));
 sg13g2_a22oi_1 _27237_ (.Y(_05514_),
    .B1(net7757),
    .B2(_05513_),
    .A2(net7878),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[30] ));
 sg13g2_nor2_1 _27238_ (.A(net9055),
    .B(net4918),
    .Y(_01263_));
 sg13g2_nand3_1 _27239_ (.B(_04835_),
    .C(_05017_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[30] ),
    .Y(_05515_));
 sg13g2_o21ai_1 _27240_ (.B1(_05515_),
    .Y(_05516_),
    .A1(_10514_),
    .A2(_05018_));
 sg13g2_nand2_1 _27241_ (.Y(_05517_),
    .A(net9229),
    .B(_05516_));
 sg13g2_xor2_1 _27242_ (.B(_05509_),
    .A(net4668),
    .X(_05518_));
 sg13g2_o21ai_1 _27243_ (.B1(_05517_),
    .Y(_05519_),
    .A1(net9236),
    .A2(_05518_));
 sg13g2_a22oi_1 _27244_ (.Y(_05520_),
    .B1(net7761),
    .B2(_05519_),
    .A2(net7878),
    .A1(net4668));
 sg13g2_nor2_1 _27245_ (.A(net9055),
    .B(net4669),
    .Y(_01264_));
 sg13g2_and2_1 _27246_ (.A(net9370),
    .B(net2600),
    .X(_01265_));
 sg13g2_o21ai_1 _27247_ (.B1(net9371),
    .Y(_05521_),
    .A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[0] ),
    .A2(net4284));
 sg13g2_a21oi_1 _27248_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[0] ),
    .A2(net4284),
    .Y(_01266_),
    .B1(_05521_));
 sg13g2_a21oi_1 _27249_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[0] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[1] ),
    .Y(_05522_),
    .B1(net3459));
 sg13g2_nand3_1 _27250_ (.B(net4284),
    .C(net3459),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[0] ),
    .Y(_05523_));
 sg13g2_nand2_1 _27251_ (.Y(_05524_),
    .A(net9371),
    .B(_05523_));
 sg13g2_nor2_1 _27252_ (.A(net3460),
    .B(_05524_),
    .Y(_01267_));
 sg13g2_and2_1 _27253_ (.A(_10651_),
    .B(_05523_),
    .X(_05525_));
 sg13g2_nor2_1 _27254_ (.A(_10651_),
    .B(_05523_),
    .Y(_05526_));
 sg13g2_nor3_1 _27255_ (.A(net9036),
    .B(net5294),
    .C(_05526_),
    .Y(_01268_));
 sg13g2_and2_1 _27256_ (.A(net5013),
    .B(_05526_),
    .X(_05527_));
 sg13g2_o21ai_1 _27257_ (.B1(net9371),
    .Y(_05528_),
    .A1(net5013),
    .A2(_05526_));
 sg13g2_nor2_1 _27258_ (.A(_05527_),
    .B(net5014),
    .Y(_01269_));
 sg13g2_xnor2_1 _27259_ (.Y(_05529_),
    .A(net4986),
    .B(_05527_));
 sg13g2_nor2_1 _27260_ (.A(net9036),
    .B(net4987),
    .Y(_01270_));
 sg13g2_a21oi_1 _27261_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[5] ),
    .A2(_05527_),
    .Y(_05530_),
    .B1(net3817));
 sg13g2_nand3_1 _27262_ (.B(net3817),
    .C(_05527_),
    .A(net4986),
    .Y(_05531_));
 sg13g2_nand2_1 _27263_ (.Y(_05532_),
    .A(net9370),
    .B(_05531_));
 sg13g2_nor2_1 _27264_ (.A(net3818),
    .B(_05532_),
    .Y(_01271_));
 sg13g2_and2_1 _27265_ (.A(_10652_),
    .B(_05531_),
    .X(_05533_));
 sg13g2_nor2_1 _27266_ (.A(_10652_),
    .B(_05531_),
    .Y(_05534_));
 sg13g2_nor3_1 _27267_ (.A(net9024),
    .B(_05533_),
    .C(_05534_),
    .Y(_01272_));
 sg13g2_and2_2 _27268_ (.A(net4717),
    .B(_05534_),
    .X(_05535_));
 sg13g2_o21ai_1 _27269_ (.B1(net9349),
    .Y(_05536_),
    .A1(net4717),
    .A2(_05534_));
 sg13g2_nor2_1 _27270_ (.A(_05535_),
    .B(net4718),
    .Y(_01273_));
 sg13g2_xnor2_1 _27271_ (.Y(_05537_),
    .A(net4734),
    .B(_05535_));
 sg13g2_nor2_1 _27272_ (.A(net9022),
    .B(_05537_),
    .Y(_01274_));
 sg13g2_a21oi_1 _27273_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[9] ),
    .A2(_05535_),
    .Y(_05538_),
    .B1(net3364));
 sg13g2_and3_2 _27274_ (.X(_05539_),
    .A(net4734),
    .B(net3364),
    .C(_05535_));
 sg13g2_nor3_1 _27275_ (.A(net9022),
    .B(net3365),
    .C(_05539_),
    .Y(_01275_));
 sg13g2_xnor2_1 _27276_ (.Y(_05540_),
    .A(net4921),
    .B(_05539_));
 sg13g2_nor2_1 _27277_ (.A(net9022),
    .B(_05540_),
    .Y(_01276_));
 sg13g2_a21oi_1 _27278_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[11] ),
    .A2(_05539_),
    .Y(_05541_),
    .B1(net3795));
 sg13g2_and3_1 _27279_ (.X(_05542_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[11] ),
    .B(net3795),
    .C(_05539_));
 sg13g2_nor3_1 _27280_ (.A(net9026),
    .B(net3796),
    .C(_05542_),
    .Y(_01277_));
 sg13g2_nor2_1 _27281_ (.A(net4499),
    .B(_05542_),
    .Y(_05543_));
 sg13g2_and2_1 _27282_ (.A(net4499),
    .B(_05542_),
    .X(_05544_));
 sg13g2_nor3_1 _27283_ (.A(net9029),
    .B(net4500),
    .C(_05544_),
    .Y(_01278_));
 sg13g2_and2_2 _27284_ (.A(net4689),
    .B(_05544_),
    .X(_05545_));
 sg13g2_o21ai_1 _27285_ (.B1(net9357),
    .Y(_05546_),
    .A1(net4689),
    .A2(_05544_));
 sg13g2_nor2_1 _27286_ (.A(_05545_),
    .B(_05546_),
    .Y(_01279_));
 sg13g2_xnor2_1 _27287_ (.Y(_05547_),
    .A(net4761),
    .B(_05545_));
 sg13g2_nor2_1 _27288_ (.A(net9028),
    .B(_05547_),
    .Y(_01280_));
 sg13g2_a21oi_1 _27289_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[15] ),
    .A2(_05545_),
    .Y(_05548_),
    .B1(net3419));
 sg13g2_and3_1 _27290_ (.X(_05549_),
    .A(net4761),
    .B(net3419),
    .C(_05545_));
 sg13g2_nor3_1 _27291_ (.A(net9028),
    .B(net3420),
    .C(_05549_),
    .Y(_01281_));
 sg13g2_xnor2_1 _27292_ (.Y(_05550_),
    .A(net4858),
    .B(_05549_));
 sg13g2_nor2_1 _27293_ (.A(net9028),
    .B(_05550_),
    .Y(_01282_));
 sg13g2_a21oi_1 _27294_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[17] ),
    .A2(_05549_),
    .Y(_05551_),
    .B1(net3933));
 sg13g2_and3_1 _27295_ (.X(_05552_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[17] ),
    .B(net3933),
    .C(_05549_));
 sg13g2_nor3_1 _27296_ (.A(net9028),
    .B(net3934),
    .C(_05552_),
    .Y(_01283_));
 sg13g2_nor2_1 _27297_ (.A(net4364),
    .B(_05552_),
    .Y(_05553_));
 sg13g2_and2_1 _27298_ (.A(net4364),
    .B(_05552_),
    .X(_05554_));
 sg13g2_nor3_1 _27299_ (.A(net9028),
    .B(net4365),
    .C(_05554_),
    .Y(_01284_));
 sg13g2_and2_1 _27300_ (.A(net5321),
    .B(_05554_),
    .X(_05555_));
 sg13g2_o21ai_1 _27301_ (.B1(net9343),
    .Y(_05556_),
    .A1(net5321),
    .A2(_05554_));
 sg13g2_nor2_1 _27302_ (.A(_05555_),
    .B(_05556_),
    .Y(_01285_));
 sg13g2_xnor2_1 _27303_ (.Y(_05557_),
    .A(net4927),
    .B(_05555_));
 sg13g2_nor2_1 _27304_ (.A(net9017),
    .B(_05557_),
    .Y(_01286_));
 sg13g2_a21oi_1 _27305_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[21] ),
    .A2(_05555_),
    .Y(_05558_),
    .B1(net3780));
 sg13g2_and3_2 _27306_ (.X(_05559_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[21] ),
    .B(net3780),
    .C(_05555_));
 sg13g2_nor3_1 _27307_ (.A(net9017),
    .B(net3781),
    .C(_05559_),
    .Y(_01287_));
 sg13g2_xnor2_1 _27308_ (.Y(_05560_),
    .A(net4961),
    .B(_05559_));
 sg13g2_nor2_1 _27309_ (.A(net9042),
    .B(net4962),
    .Y(_01288_));
 sg13g2_a21oi_1 _27310_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[23] ),
    .A2(_05559_),
    .Y(_05561_),
    .B1(net3760));
 sg13g2_and3_1 _27311_ (.X(_05562_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[23] ),
    .B(net3760),
    .C(_05559_));
 sg13g2_nor3_1 _27312_ (.A(net9042),
    .B(net3761),
    .C(_05562_),
    .Y(_01289_));
 sg13g2_nor2_1 _27313_ (.A(net4374),
    .B(_05562_),
    .Y(_05563_));
 sg13g2_and2_1 _27314_ (.A(net4374),
    .B(_05562_),
    .X(_05564_));
 sg13g2_nor3_1 _27315_ (.A(net9042),
    .B(net4375),
    .C(_05564_),
    .Y(_01290_));
 sg13g2_and2_1 _27316_ (.A(net4806),
    .B(_05564_),
    .X(_05565_));
 sg13g2_o21ai_1 _27317_ (.B1(net9383),
    .Y(_05566_),
    .A1(net4806),
    .A2(_05564_));
 sg13g2_nor2_1 _27318_ (.A(_05565_),
    .B(_05566_),
    .Y(_01291_));
 sg13g2_xnor2_1 _27319_ (.Y(_05567_),
    .A(net4714),
    .B(_05565_));
 sg13g2_nor2_1 _27320_ (.A(net9041),
    .B(net4715),
    .Y(_01292_));
 sg13g2_a21oi_1 _27321_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[27] ),
    .A2(_05565_),
    .Y(_05568_),
    .B1(net2828));
 sg13g2_and3_1 _27322_ (.X(_05569_),
    .A(net4714),
    .B(net2828),
    .C(_05565_));
 sg13g2_nor3_1 _27323_ (.A(net9041),
    .B(net2829),
    .C(_05569_),
    .Y(_01293_));
 sg13g2_xnor2_1 _27324_ (.Y(_05570_),
    .A(net4748),
    .B(_05569_));
 sg13g2_nor2_1 _27325_ (.A(net9041),
    .B(_05570_),
    .Y(_01294_));
 sg13g2_a21oi_1 _27326_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[29] ),
    .A2(_05569_),
    .Y(_05571_),
    .B1(net3254));
 sg13g2_and3_2 _27327_ (.X(_05572_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[29] ),
    .B(net3254),
    .C(_05569_));
 sg13g2_nor3_1 _27328_ (.A(net9041),
    .B(net3255),
    .C(_05572_),
    .Y(_01295_));
 sg13g2_nor2_1 _27329_ (.A(net4201),
    .B(_05572_),
    .Y(_05573_));
 sg13g2_and2_1 _27330_ (.A(net4201),
    .B(_05572_),
    .X(_05574_));
 sg13g2_nor3_1 _27331_ (.A(net9040),
    .B(net4202),
    .C(_05574_),
    .Y(_01296_));
 sg13g2_and2_2 _27332_ (.A(net4843),
    .B(_05574_),
    .X(_05575_));
 sg13g2_o21ai_1 _27333_ (.B1(net9382),
    .Y(_05576_),
    .A1(net4843),
    .A2(_05574_));
 sg13g2_nor2_1 _27334_ (.A(_05575_),
    .B(_05576_),
    .Y(_01297_));
 sg13g2_xnor2_1 _27335_ (.Y(_05577_),
    .A(net4879),
    .B(_05575_));
 sg13g2_nor2_1 _27336_ (.A(net9035),
    .B(_05577_),
    .Y(_01298_));
 sg13g2_a21oi_1 _27337_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[33] ),
    .A2(_05575_),
    .Y(_05578_),
    .B1(net3688));
 sg13g2_and3_1 _27338_ (.X(_05579_),
    .A(net4879),
    .B(net3688),
    .C(_05575_));
 sg13g2_nor3_1 _27339_ (.A(net9035),
    .B(net3689),
    .C(_05579_),
    .Y(_01299_));
 sg13g2_xnor2_1 _27340_ (.Y(_05580_),
    .A(net4953),
    .B(_05579_));
 sg13g2_nor2_1 _27341_ (.A(net9035),
    .B(_05580_),
    .Y(_01300_));
 sg13g2_a21oi_1 _27342_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[35] ),
    .A2(_05579_),
    .Y(_05581_),
    .B1(net4343));
 sg13g2_and3_1 _27343_ (.X(_05582_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[35] ),
    .B(net4343),
    .C(_05579_));
 sg13g2_nor3_1 _27344_ (.A(net9035),
    .B(net4344),
    .C(_05582_),
    .Y(_01301_));
 sg13g2_nor2_1 _27345_ (.A(net4723),
    .B(_05582_),
    .Y(_05583_));
 sg13g2_and2_1 _27346_ (.A(net4723),
    .B(_05582_),
    .X(_05584_));
 sg13g2_nor3_1 _27347_ (.A(net9035),
    .B(net4724),
    .C(_05584_),
    .Y(_01302_));
 sg13g2_and2_1 _27348_ (.A(net5080),
    .B(_05584_),
    .X(_05585_));
 sg13g2_o21ai_1 _27349_ (.B1(net9370),
    .Y(_05586_),
    .A1(net5080),
    .A2(_05584_));
 sg13g2_nor2_1 _27350_ (.A(_05585_),
    .B(_05586_),
    .Y(_01303_));
 sg13g2_xnor2_1 _27351_ (.Y(_05587_),
    .A(net4940),
    .B(_05585_));
 sg13g2_nor2_1 _27352_ (.A(net9024),
    .B(net4941),
    .Y(_01304_));
 sg13g2_a21oi_1 _27353_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[39] ),
    .A2(_05585_),
    .Y(_05588_),
    .B1(net3737));
 sg13g2_and3_2 _27354_ (.X(_05589_),
    .A(net5569),
    .B(net3737),
    .C(_05585_));
 sg13g2_nor3_1 _27355_ (.A(net9024),
    .B(net3738),
    .C(_05589_),
    .Y(_01305_));
 sg13g2_xnor2_1 _27356_ (.Y(_05590_),
    .A(net4809),
    .B(_05589_));
 sg13g2_nor2_1 _27357_ (.A(net9023),
    .B(net4810),
    .Y(_01306_));
 sg13g2_a21oi_1 _27358_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[41] ),
    .A2(_05589_),
    .Y(_05591_),
    .B1(net3710));
 sg13g2_and3_1 _27359_ (.X(_05592_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[41] ),
    .B(net3710),
    .C(_05589_));
 sg13g2_nor3_1 _27360_ (.A(net9023),
    .B(net3711),
    .C(_05592_),
    .Y(_01307_));
 sg13g2_nor2_1 _27361_ (.A(net4168),
    .B(_05592_),
    .Y(_05593_));
 sg13g2_and2_2 _27362_ (.A(net4168),
    .B(_05592_),
    .X(_05594_));
 sg13g2_nor3_1 _27363_ (.A(net9023),
    .B(net4169),
    .C(_05594_),
    .Y(_01308_));
 sg13g2_and2_2 _27364_ (.A(net5045),
    .B(_05594_),
    .X(_05595_));
 sg13g2_o21ai_1 _27365_ (.B1(net9362),
    .Y(_05596_),
    .A1(net5045),
    .A2(_05594_));
 sg13g2_nor2_1 _27366_ (.A(_05595_),
    .B(_05596_),
    .Y(_01309_));
 sg13g2_xnor2_1 _27367_ (.Y(_05597_),
    .A(net4893),
    .B(_05595_));
 sg13g2_nor2_1 _27368_ (.A(net9029),
    .B(net4894),
    .Y(_01310_));
 sg13g2_a21oi_1 _27369_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[45] ),
    .A2(_05595_),
    .Y(_05598_),
    .B1(net3309));
 sg13g2_and3_2 _27370_ (.X(_05599_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[45] ),
    .B(net3309),
    .C(_05595_));
 sg13g2_nor3_1 _27371_ (.A(net9019),
    .B(net3310),
    .C(_05599_),
    .Y(_01311_));
 sg13g2_xnor2_1 _27372_ (.Y(_05600_),
    .A(net4813),
    .B(_05599_));
 sg13g2_nor2_1 _27373_ (.A(net9017),
    .B(net4814),
    .Y(_01312_));
 sg13g2_a21oi_1 _27374_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[47] ),
    .A2(_05599_),
    .Y(_05601_),
    .B1(net3774));
 sg13g2_and3_1 _27375_ (.X(_05602_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[47] ),
    .B(net3774),
    .C(_05599_));
 sg13g2_nor3_1 _27376_ (.A(net9017),
    .B(net3775),
    .C(_05602_),
    .Y(_01313_));
 sg13g2_nor2_1 _27377_ (.A(net4389),
    .B(_05602_),
    .Y(_05603_));
 sg13g2_and2_1 _27378_ (.A(net4389),
    .B(_05602_),
    .X(_05604_));
 sg13g2_nor3_1 _27379_ (.A(net9017),
    .B(net4390),
    .C(_05604_),
    .Y(_01314_));
 sg13g2_and2_1 _27380_ (.A(net4926),
    .B(_05604_),
    .X(_05605_));
 sg13g2_o21ai_1 _27381_ (.B1(net9358),
    .Y(_05606_),
    .A1(net4926),
    .A2(_05604_));
 sg13g2_nor2_1 _27382_ (.A(_05605_),
    .B(_05606_),
    .Y(_01315_));
 sg13g2_xnor2_1 _27383_ (.Y(_05607_),
    .A(net5011),
    .B(_05605_));
 sg13g2_nor2_1 _27384_ (.A(net9028),
    .B(_05607_),
    .Y(_01316_));
 sg13g2_a21oi_1 _27385_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[51] ),
    .A2(_05605_),
    .Y(_05608_),
    .B1(net3484));
 sg13g2_and3_1 _27386_ (.X(_05609_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[51] ),
    .B(net3484),
    .C(_05605_));
 sg13g2_nor3_1 _27387_ (.A(net9028),
    .B(net3485),
    .C(_05609_),
    .Y(_01317_));
 sg13g2_xnor2_1 _27388_ (.Y(_05610_),
    .A(net4636),
    .B(_05609_));
 sg13g2_nor2_1 _27389_ (.A(net9028),
    .B(net4637),
    .Y(_01318_));
 sg13g2_a21oi_1 _27390_ (.A1(net4636),
    .A2(_05609_),
    .Y(_05611_),
    .B1(net4942));
 sg13g2_and3_2 _27391_ (.X(_05612_),
    .A(net4636),
    .B(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[54] ),
    .C(_05609_));
 sg13g2_nor3_1 _27392_ (.A(net9017),
    .B(net4943),
    .C(_05612_),
    .Y(_01319_));
 sg13g2_nor2_1 _27393_ (.A(net4148),
    .B(_05612_),
    .Y(_05613_));
 sg13g2_and2_1 _27394_ (.A(net4148),
    .B(_05612_),
    .X(_05614_));
 sg13g2_nor3_1 _27395_ (.A(net9030),
    .B(net4149),
    .C(_05614_),
    .Y(_01320_));
 sg13g2_and2_1 _27396_ (.A(net4763),
    .B(_05614_),
    .X(_05615_));
 sg13g2_o21ai_1 _27397_ (.B1(net9384),
    .Y(_05616_),
    .A1(net4763),
    .A2(_05614_));
 sg13g2_nor2_1 _27398_ (.A(_05615_),
    .B(_05616_),
    .Y(_01321_));
 sg13g2_xnor2_1 _27399_ (.Y(_05617_),
    .A(net4594),
    .B(_05615_));
 sg13g2_nor2_1 _27400_ (.A(net9042),
    .B(net4595),
    .Y(_01322_));
 sg13g2_a21oi_1 _27401_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[57] ),
    .A2(_05615_),
    .Y(_05618_),
    .B1(net3205));
 sg13g2_and3_1 _27402_ (.X(_05619_),
    .A(net4594),
    .B(net3205),
    .C(_05615_));
 sg13g2_nor3_1 _27403_ (.A(net9032),
    .B(net3206),
    .C(_05619_),
    .Y(_01323_));
 sg13g2_xnor2_1 _27404_ (.Y(_05620_),
    .A(net5176),
    .B(_05619_));
 sg13g2_nor2_1 _27405_ (.A(net9030),
    .B(_05620_),
    .Y(_01324_));
 sg13g2_a21oi_1 _27406_ (.A1(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[59] ),
    .A2(_05619_),
    .Y(_05621_),
    .B1(net3471));
 sg13g2_and3_1 _27407_ (.X(_05622_),
    .A(net5570),
    .B(net3471),
    .C(_05619_));
 sg13g2_nor3_1 _27408_ (.A(net9032),
    .B(net3472),
    .C(_05622_),
    .Y(_01325_));
 sg13g2_nor2_1 _27409_ (.A(net4301),
    .B(_05622_),
    .Y(_05623_));
 sg13g2_and2_1 _27410_ (.A(net4301),
    .B(_05622_),
    .X(_05624_));
 sg13g2_nor3_1 _27411_ (.A(net9030),
    .B(net4302),
    .C(_05624_),
    .Y(_01326_));
 sg13g2_nand2_1 _27412_ (.Y(_05625_),
    .A(net4793),
    .B(_05624_));
 sg13g2_o21ai_1 _27413_ (.B1(net9364),
    .Y(_05626_),
    .A1(net4793),
    .A2(_05624_));
 sg13g2_nor2b_1 _27414_ (.A(_05626_),
    .B_N(_05625_),
    .Y(_01327_));
 sg13g2_o21ai_1 _27415_ (.B1(net9362),
    .Y(_05627_),
    .A1(_10653_),
    .A2(_05625_));
 sg13g2_a21oi_1 _27416_ (.A1(_10653_),
    .A2(_05625_),
    .Y(_01328_),
    .B1(_05627_));
 sg13g2_a21oi_1 _27417_ (.A1(net9226),
    .A2(_05024_),
    .Y(_05628_),
    .B1(net3757));
 sg13g2_a21oi_2 _27418_ (.B1(_05027_),
    .Y(_05629_),
    .A2(_05023_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_state[0] ));
 sg13g2_o21ai_1 _27419_ (.B1(_05024_),
    .Y(_05630_),
    .A1(\soc_I.kianv_I.datapath_unit_I.div_I.div_state[0] ),
    .A2(net9226));
 sg13g2_a21oi_1 _27420_ (.A1(net3757),
    .A2(_05629_),
    .Y(_05631_),
    .B1(net9054));
 sg13g2_nor2b_1 _27421_ (.A(net3758),
    .B_N(_05631_),
    .Y(_01329_));
 sg13g2_a21oi_1 _27422_ (.A1(\soc_I.kianv_I.datapath_unit_I.div_I.bit_idx[0] ),
    .A2(_05629_),
    .Y(_05632_),
    .B1(net2869));
 sg13g2_and2_1 _27423_ (.A(net2869),
    .B(net3757),
    .X(_05633_));
 sg13g2_nor2b_1 _27424_ (.A(_05633_),
    .B_N(net9226),
    .Y(_05634_));
 sg13g2_o21ai_1 _27425_ (.B1(net9411),
    .Y(_05635_),
    .A1(_05630_),
    .A2(_05634_));
 sg13g2_nor2_1 _27426_ (.A(net2870),
    .B(_05635_),
    .Y(_01330_));
 sg13g2_a21oi_1 _27427_ (.A1(_05629_),
    .A2(_05633_),
    .Y(_05636_),
    .B1(net3978));
 sg13g2_nand2_1 _27428_ (.Y(_05637_),
    .A(net3978),
    .B(_05633_));
 sg13g2_a21oi_1 _27429_ (.A1(net9226),
    .A2(_05637_),
    .Y(_05638_),
    .B1(_05630_));
 sg13g2_nor3_1 _27430_ (.A(net9054),
    .B(_05636_),
    .C(_05638_),
    .Y(_01331_));
 sg13g2_nand4_1 _27431_ (.B(net9226),
    .C(_05024_),
    .A(net3978),
    .Y(_05639_),
    .D(_05633_));
 sg13g2_mux2_1 _27432_ (.A0(_05639_),
    .A1(_05638_),
    .S(net4931),
    .X(_05640_));
 sg13g2_nor2_1 _27433_ (.A(net9054),
    .B(_05640_),
    .Y(_01332_));
 sg13g2_nand3_1 _27434_ (.B(net3978),
    .C(_05633_),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.bit_idx[3] ),
    .Y(_05641_));
 sg13g2_o21ai_1 _27435_ (.B1(net9226),
    .Y(_05642_),
    .A1(net2601),
    .A2(_05641_));
 sg13g2_a21o_1 _27436_ (.A2(_05641_),
    .A1(net2601),
    .B1(_05642_),
    .X(_05643_));
 sg13g2_o21ai_1 _27437_ (.B1(net9411),
    .Y(_05644_),
    .A1(net4298),
    .A2(_05629_));
 sg13g2_a21oi_1 _27438_ (.A1(_05629_),
    .A2(_05643_),
    .Y(_01333_),
    .B1(_05644_));
 sg13g2_a21oi_1 _27439_ (.A1(net5302),
    .A2(_10592_),
    .Y(_05645_),
    .B1(net9237));
 sg13g2_nor2_1 _27440_ (.A(net9054),
    .B(net5303),
    .Y(_01334_));
 sg13g2_nor3_2 _27441_ (.A(\soc_I.kianv_I.control_unit_I.mul_ready ),
    .B(net4610),
    .C(net8617),
    .Y(_05646_));
 sg13g2_and2_1 _27442_ (.A(net9001),
    .B(_05646_),
    .X(_05647_));
 sg13g2_nand2_1 _27443_ (.Y(_05648_),
    .A(net9001),
    .B(_05646_));
 sg13g2_nor2_1 _27444_ (.A(net4880),
    .B(net8466),
    .Y(_05649_));
 sg13g2_a21oi_1 _27445_ (.A1(net8298),
    .A2(net8466),
    .Y(_01335_),
    .B1(_05649_));
 sg13g2_nand2_1 _27446_ (.Y(_05650_),
    .A(net5096),
    .B(net8456));
 sg13g2_xnor2_1 _27447_ (.Y(_05651_),
    .A(_10924_),
    .B(_13289_));
 sg13g2_nor2_2 _27448_ (.A(net8315),
    .B(_05651_),
    .Y(_05652_));
 sg13g2_or2_1 _27449_ (.X(_05653_),
    .B(_05651_),
    .A(net8315));
 sg13g2_nor2_1 _27450_ (.A(_05040_),
    .B(net7972),
    .Y(_05654_));
 sg13g2_o21ai_1 _27451_ (.B1(net8466),
    .Y(_05655_),
    .A1(net8299),
    .A2(net7973));
 sg13g2_o21ai_1 _27452_ (.B1(_05650_),
    .Y(_01336_),
    .A1(_05654_),
    .A2(_05655_));
 sg13g2_o21ai_1 _27453_ (.B1(net8467),
    .Y(_05656_),
    .A1(_11144_),
    .A2(net7976));
 sg13g2_a21oi_2 _27454_ (.B1(_05656_),
    .Y(_05657_),
    .A2(net7973),
    .A1(_05046_));
 sg13g2_a21o_1 _27455_ (.A2(net8462),
    .A1(net4414),
    .B1(_05657_),
    .X(_01337_));
 sg13g2_o21ai_1 _27456_ (.B1(net8466),
    .Y(_05658_),
    .A1(net8301),
    .A2(net7973));
 sg13g2_a21oi_2 _27457_ (.B1(_05658_),
    .Y(_05659_),
    .A2(net7973),
    .A1(_05055_));
 sg13g2_a21o_1 _27458_ (.A2(net8459),
    .A1(net5002),
    .B1(_05659_),
    .X(_01338_));
 sg13g2_a21oi_1 _27459_ (.A1(net8303),
    .A2(net7972),
    .Y(_05660_),
    .B1(net8456));
 sg13g2_o21ai_1 _27460_ (.B1(_05660_),
    .Y(_05661_),
    .A1(_05063_),
    .A2(net7972));
 sg13g2_o21ai_1 _27461_ (.B1(_05661_),
    .Y(_01339_),
    .A1(_10623_),
    .A2(net8475));
 sg13g2_o21ai_1 _27462_ (.B1(net8466),
    .Y(_05662_),
    .A1(net8304),
    .A2(net7974));
 sg13g2_a21oi_2 _27463_ (.B1(_05662_),
    .Y(_05663_),
    .A2(net7974),
    .A1(_05070_));
 sg13g2_a21o_1 _27464_ (.A2(net8459),
    .A1(net4427),
    .B1(_05663_),
    .X(_01340_));
 sg13g2_o21ai_1 _27465_ (.B1(net8466),
    .Y(_05664_),
    .A1(_11096_),
    .A2(net7973));
 sg13g2_a21o_2 _27466_ (.A2(net7973),
    .A1(_05079_),
    .B1(_05664_),
    .X(_05665_));
 sg13g2_o21ai_1 _27467_ (.B1(_05665_),
    .Y(_01341_),
    .A1(_10624_),
    .A2(net8475));
 sg13g2_o21ai_1 _27468_ (.B1(net8467),
    .Y(_05666_),
    .A1(_11086_),
    .A2(net7976));
 sg13g2_a21oi_2 _27469_ (.B1(_05666_),
    .Y(_05667_),
    .A2(net7976),
    .A1(_05088_));
 sg13g2_a21o_1 _27470_ (.A2(net8463),
    .A1(net4376),
    .B1(_05667_),
    .X(_01342_));
 sg13g2_nand2_1 _27471_ (.Y(_05668_),
    .A(_05097_),
    .B(net7973));
 sg13g2_a21oi_1 _27472_ (.A1(_11207_),
    .A2(net7972),
    .Y(_05669_),
    .B1(net8456));
 sg13g2_a22oi_1 _27473_ (.Y(_05670_),
    .B1(_05668_),
    .B2(_05669_),
    .A2(net8456),
    .A1(net5008));
 sg13g2_inv_1 _27474_ (.Y(_01343_),
    .A(_05670_));
 sg13g2_o21ai_1 _27475_ (.B1(net8469),
    .Y(_05671_),
    .A1(_11247_),
    .A2(net7974));
 sg13g2_a21oi_2 _27476_ (.B1(_05671_),
    .Y(_05672_),
    .A2(net7974),
    .A1(_05105_));
 sg13g2_a21o_1 _27477_ (.A2(net8462),
    .A1(net4455),
    .B1(_05672_),
    .X(_01344_));
 sg13g2_nand2_1 _27478_ (.Y(_05673_),
    .A(_05114_),
    .B(net7973));
 sg13g2_a21oi_1 _27479_ (.A1(_11221_),
    .A2(net7972),
    .Y(_05674_),
    .B1(net8456));
 sg13g2_a22oi_1 _27480_ (.Y(_05675_),
    .B1(_05673_),
    .B2(_05674_),
    .A2(net8458),
    .A1(net5036));
 sg13g2_inv_1 _27481_ (.Y(_01345_),
    .A(_05675_));
 sg13g2_o21ai_1 _27482_ (.B1(net8467),
    .Y(_05676_),
    .A1(net8296),
    .A2(net7974));
 sg13g2_a21oi_2 _27483_ (.B1(_05676_),
    .Y(_05677_),
    .A2(net7974),
    .A1(_05123_));
 sg13g2_a21o_1 _27484_ (.A2(net8462),
    .A1(net4833),
    .B1(_05677_),
    .X(_01346_));
 sg13g2_o21ai_1 _27485_ (.B1(net8468),
    .Y(_05678_),
    .A1(net8292),
    .A2(net7975));
 sg13g2_a21oi_2 _27486_ (.B1(_05678_),
    .Y(_05679_),
    .A2(net7975),
    .A1(_05131_));
 sg13g2_a21o_1 _27487_ (.A2(net8462),
    .A1(net4450),
    .B1(_05679_),
    .X(_01347_));
 sg13g2_nand2_2 _27488_ (.Y(_05680_),
    .A(_05140_),
    .B(net7975));
 sg13g2_a21oi_2 _27489_ (.B1(net8459),
    .Y(_05681_),
    .A2(net7972),
    .A1(net8291));
 sg13g2_a22oi_1 _27490_ (.Y(_05682_),
    .B1(_05680_),
    .B2(_05681_),
    .A2(net8463),
    .A1(net3604));
 sg13g2_inv_1 _27491_ (.Y(_01348_),
    .A(_05682_));
 sg13g2_nand2_1 _27492_ (.Y(_05683_),
    .A(_05149_),
    .B(net7978));
 sg13g2_a21oi_1 _27493_ (.A1(net8295),
    .A2(net7971),
    .Y(_05684_),
    .B1(net8460));
 sg13g2_a22oi_1 _27494_ (.Y(_05685_),
    .B1(_05683_),
    .B2(_05684_),
    .A2(net8460),
    .A1(net4702));
 sg13g2_inv_1 _27495_ (.Y(_01349_),
    .A(_05685_));
 sg13g2_o21ai_1 _27496_ (.B1(net8471),
    .Y(_05686_),
    .A1(net8293),
    .A2(net7978));
 sg13g2_a21oi_2 _27497_ (.B1(_05686_),
    .Y(_05687_),
    .A2(net7978),
    .A1(_05157_));
 sg13g2_a21o_1 _27498_ (.A2(net8464),
    .A1(net3674),
    .B1(_05687_),
    .X(_01350_));
 sg13g2_nand2_1 _27499_ (.Y(_05688_),
    .A(_05166_),
    .B(net7977));
 sg13g2_a21oi_1 _27500_ (.A1(net8283),
    .A2(net7971),
    .Y(_05689_),
    .B1(net8455));
 sg13g2_a22oi_1 _27501_ (.Y(_05690_),
    .B1(_05688_),
    .B2(_05689_),
    .A2(net8460),
    .A1(net4421));
 sg13g2_inv_1 _27502_ (.Y(_01351_),
    .A(_05690_));
 sg13g2_o21ai_1 _27503_ (.B1(net8470),
    .Y(_05691_),
    .A1(net8276),
    .A2(net7977));
 sg13g2_a21oi_2 _27504_ (.B1(_05691_),
    .Y(_05692_),
    .A2(net7978),
    .A1(_05175_));
 sg13g2_a21o_1 _27505_ (.A2(net8464),
    .A1(net4245),
    .B1(_05692_),
    .X(_01352_));
 sg13g2_nand2_1 _27506_ (.Y(_05693_),
    .A(_05184_),
    .B(net7977));
 sg13g2_a21oi_1 _27507_ (.A1(net8281),
    .A2(net7971),
    .Y(_05694_),
    .B1(net8460));
 sg13g2_a22oi_1 _27508_ (.Y(_05695_),
    .B1(_05693_),
    .B2(_05694_),
    .A2(net8460),
    .A1(net4399));
 sg13g2_inv_1 _27509_ (.Y(_01353_),
    .A(_05695_));
 sg13g2_o21ai_1 _27510_ (.B1(net8471),
    .Y(_05696_),
    .A1(net8279),
    .A2(net7978));
 sg13g2_a21oi_1 _27511_ (.A1(_05193_),
    .A2(net7978),
    .Y(_05697_),
    .B1(_05696_));
 sg13g2_a21o_1 _27512_ (.A2(net8460),
    .A1(net4360),
    .B1(_05697_),
    .X(_01354_));
 sg13g2_nand2_1 _27513_ (.Y(_05698_),
    .A(_05202_),
    .B(net7977));
 sg13g2_a21oi_1 _27514_ (.A1(net8286),
    .A2(net7971),
    .Y(_05699_),
    .B1(net8455));
 sg13g2_a22oi_1 _27515_ (.Y(_05700_),
    .B1(_05698_),
    .B2(_05699_),
    .A2(net8454),
    .A1(net4138));
 sg13g2_inv_1 _27516_ (.Y(_01355_),
    .A(_05700_));
 sg13g2_o21ai_1 _27517_ (.B1(net8470),
    .Y(_05701_),
    .A1(net8284),
    .A2(net7977));
 sg13g2_a21oi_2 _27518_ (.B1(_05701_),
    .Y(_05702_),
    .A2(net7977),
    .A1(_05210_));
 sg13g2_a21o_1 _27519_ (.A2(net8464),
    .A1(net4569),
    .B1(_05702_),
    .X(_01356_));
 sg13g2_nand2_1 _27520_ (.Y(_05703_),
    .A(_05219_),
    .B(net7977));
 sg13g2_a21oi_1 _27521_ (.A1(net8288),
    .A2(net7971),
    .Y(_05704_),
    .B1(net8455));
 sg13g2_a22oi_1 _27522_ (.Y(_05705_),
    .B1(_05703_),
    .B2(_05704_),
    .A2(net8460),
    .A1(net4261));
 sg13g2_inv_1 _27523_ (.Y(_01357_),
    .A(_05705_));
 sg13g2_o21ai_1 _27524_ (.B1(net8470),
    .Y(_05706_),
    .A1(net8287),
    .A2(net7979));
 sg13g2_a21oi_2 _27525_ (.B1(_05706_),
    .Y(_05707_),
    .A2(net7977),
    .A1(_05228_));
 sg13g2_a21o_1 _27526_ (.A2(net8464),
    .A1(net3962),
    .B1(_05707_),
    .X(_01358_));
 sg13g2_nand2_1 _27527_ (.Y(_05708_),
    .A(_05236_),
    .B(net7979));
 sg13g2_a21oi_1 _27528_ (.A1(net8271),
    .A2(net7970),
    .Y(_05709_),
    .B1(net8454));
 sg13g2_a22oi_1 _27529_ (.Y(_05710_),
    .B1(_05708_),
    .B2(_05709_),
    .A2(net8455),
    .A1(net4824));
 sg13g2_inv_1 _27530_ (.Y(_01359_),
    .A(_05710_));
 sg13g2_nand2_1 _27531_ (.Y(_05711_),
    .A(_05246_),
    .B(net7979));
 sg13g2_a21oi_1 _27532_ (.A1(net8270),
    .A2(net7971),
    .Y(_05712_),
    .B1(net8454));
 sg13g2_a22oi_1 _27533_ (.Y(_05713_),
    .B1(_05711_),
    .B2(_05712_),
    .A2(net8454),
    .A1(net5129));
 sg13g2_inv_1 _27534_ (.Y(_01360_),
    .A(_05713_));
 sg13g2_nand2_1 _27535_ (.Y(_05714_),
    .A(net8275),
    .B(net7970));
 sg13g2_o21ai_1 _27536_ (.B1(_05714_),
    .Y(_05715_),
    .A1(_05255_),
    .A2(net7970));
 sg13g2_nor2_2 _27537_ (.A(net8454),
    .B(_05715_),
    .Y(_05716_));
 sg13g2_a21oi_1 _27538_ (.A1(net3701),
    .A2(net8465),
    .Y(_05717_),
    .B1(_05716_));
 sg13g2_inv_1 _27539_ (.Y(_01361_),
    .A(_05717_));
 sg13g2_o21ai_1 _27540_ (.B1(net8470),
    .Y(_05718_),
    .A1(net8273),
    .A2(net7979));
 sg13g2_a21oi_2 _27541_ (.B1(_05718_),
    .Y(_05719_),
    .A2(net7979),
    .A1(_05263_));
 sg13g2_a21o_1 _27542_ (.A2(net8465),
    .A1(net3857),
    .B1(_05719_),
    .X(_01362_));
 sg13g2_nand2_1 _27543_ (.Y(_05720_),
    .A(_05272_),
    .B(net7979));
 sg13g2_a21oi_1 _27544_ (.A1(net8268),
    .A2(net7970),
    .Y(_05721_),
    .B1(net8457));
 sg13g2_a22oi_1 _27545_ (.Y(_05722_),
    .B1(_05720_),
    .B2(_05721_),
    .A2(net8457),
    .A1(net5116));
 sg13g2_inv_1 _27546_ (.Y(_01363_),
    .A(_05722_));
 sg13g2_nand2_1 _27547_ (.Y(_05723_),
    .A(net8307),
    .B(net7970));
 sg13g2_o21ai_1 _27548_ (.B1(_05723_),
    .Y(_05724_),
    .A1(_05281_),
    .A2(net7970));
 sg13g2_nor2_2 _27549_ (.A(net8454),
    .B(_05724_),
    .Y(_05725_));
 sg13g2_a21oi_1 _27550_ (.A1(net4126),
    .A2(net8454),
    .Y(_05726_),
    .B1(_05725_));
 sg13g2_inv_1 _27551_ (.Y(_01364_),
    .A(_05726_));
 sg13g2_a21oi_1 _27552_ (.A1(_11052_),
    .A2(net7970),
    .Y(_05727_),
    .B1(net8454));
 sg13g2_o21ai_1 _27553_ (.B1(_05727_),
    .Y(_05728_),
    .A1(_05289_),
    .A2(net7970));
 sg13g2_o21ai_1 _27554_ (.B1(_05728_),
    .Y(_01365_),
    .A1(_10633_),
    .A2(net8470));
 sg13g2_nor2_1 _27555_ (.A(_05288_),
    .B(_05651_),
    .Y(_05729_));
 sg13g2_nor3_2 _27556_ (.A(net8314),
    .B(net8457),
    .C(_05729_),
    .Y(_05730_));
 sg13g2_a21o_1 _27557_ (.A2(net8464),
    .A1(net4468),
    .B1(_05730_),
    .X(_01366_));
 sg13g2_o21ai_1 _27558_ (.B1(net5048),
    .Y(_05731_),
    .A1(\soc_I.kianv_I.control_unit_I.mul_ready ),
    .A2(net8617));
 sg13g2_a21oi_1 _27559_ (.A1(net8984),
    .A2(net4610),
    .Y(_05732_),
    .B1(_05731_));
 sg13g2_or3_1 _27560_ (.A(net9217),
    .B(net9060),
    .C(_05732_),
    .X(_01367_));
 sg13g2_or2_1 _27561_ (.X(_05733_),
    .B(net5471),
    .A(net9209));
 sg13g2_and2_2 _27562_ (.A(_05731_),
    .B(_05733_),
    .X(_05734_));
 sg13g2_nand2_1 _27563_ (.Y(_05735_),
    .A(_05731_),
    .B(_05733_));
 sg13g2_nor2_1 _27564_ (.A(net9060),
    .B(net8984),
    .Y(_05736_));
 sg13g2_a22oi_1 _27565_ (.Y(_05737_),
    .B1(_05731_),
    .B2(_05736_),
    .A2(net9416),
    .A1(net9759));
 sg13g2_a21oi_1 _27566_ (.A1(net9759),
    .A2(_05734_),
    .Y(_01368_),
    .B1(_05737_));
 sg13g2_a21oi_1 _27567_ (.A1(net9759),
    .A2(_05734_),
    .Y(_05738_),
    .B1(net9752));
 sg13g2_and2_1 _27568_ (.A(net9752),
    .B(net9759),
    .X(_05739_));
 sg13g2_nand2_1 _27569_ (.Y(_05740_),
    .A(net9752),
    .B(net9759));
 sg13g2_a22oi_1 _27570_ (.Y(_05741_),
    .B1(_05736_),
    .B2(_05740_),
    .A2(_05735_),
    .A1(net9416));
 sg13g2_nor2_1 _27571_ (.A(_05738_),
    .B(_05741_),
    .Y(_01369_));
 sg13g2_nand2b_1 _27572_ (.Y(_05742_),
    .B(_05739_),
    .A_N(_00255_));
 sg13g2_a21oi_1 _27573_ (.A1(_00255_),
    .A2(_05740_),
    .Y(_05743_),
    .B1(net8984));
 sg13g2_nand2_1 _27574_ (.Y(_05744_),
    .A(_05742_),
    .B(_05743_));
 sg13g2_o21ai_1 _27575_ (.B1(net9416),
    .Y(_05745_),
    .A1(net9744),
    .A2(_05734_));
 sg13g2_a21oi_1 _27576_ (.A1(_05734_),
    .A2(_05744_),
    .Y(_01370_),
    .B1(_05745_));
 sg13g2_a21oi_1 _27577_ (.A1(net9732),
    .A2(_05742_),
    .Y(_05746_),
    .B1(net8984));
 sg13g2_o21ai_1 _27578_ (.B1(_05746_),
    .Y(_05747_),
    .A1(net9732),
    .A2(_05742_));
 sg13g2_o21ai_1 _27579_ (.B1(net9416),
    .Y(_05748_),
    .A1(net9740),
    .A2(_05734_));
 sg13g2_a21oi_1 _27580_ (.A1(_05734_),
    .A2(_05747_),
    .Y(_01371_),
    .B1(_05748_));
 sg13g2_nand2_1 _27581_ (.Y(_05749_),
    .A(net9740),
    .B(net9744));
 sg13g2_or2_1 _27582_ (.X(_05750_),
    .B(_05749_),
    .A(_05740_));
 sg13g2_o21ai_1 _27583_ (.B1(net9209),
    .Y(_05751_),
    .A1(net9718),
    .A2(_05750_));
 sg13g2_a21oi_1 _27584_ (.A1(net9718),
    .A2(_05750_),
    .Y(_05752_),
    .B1(_05751_));
 sg13g2_nand2_1 _27585_ (.Y(_05753_),
    .A(_05734_),
    .B(_05752_));
 sg13g2_nand2_1 _27586_ (.Y(_05754_),
    .A(net9719),
    .B(_05735_));
 sg13g2_a21oi_1 _27587_ (.A1(_05753_),
    .A2(_05754_),
    .Y(_01372_),
    .B1(net9060));
 sg13g2_nand3_1 _27588_ (.B(net9411),
    .C(_05024_),
    .A(net9063),
    .Y(_01373_));
 sg13g2_nand2b_1 _27589_ (.Y(_05755_),
    .B(\soc_I.kianv_I.control_unit_I.mul_ready ),
    .A_N(net5048));
 sg13g2_a21oi_1 _27590_ (.A1(net9078),
    .A2(net5049),
    .Y(_01374_),
    .B1(net9060));
 sg13g2_nor2_1 _27591_ (.A(net8857),
    .B(net8728),
    .Y(_05756_));
 sg13g2_a22oi_1 _27592_ (.Y(_05757_),
    .B1(net8586),
    .B2(net5565),
    .A2(\soc_I.kianv_I.datapath_unit_I.Data[0] ),
    .A1(net8854));
 sg13g2_o21ai_1 _27593_ (.B1(_05757_),
    .Y(_05758_),
    .A1(_10865_),
    .A2(_11729_));
 sg13g2_and2_1 _27594_ (.A(net9386),
    .B(_05758_),
    .X(_01375_));
 sg13g2_nor2_1 _27595_ (.A(_10865_),
    .B(_11837_),
    .Y(_05759_));
 sg13g2_a221oi_1 _27596_ (.B2(net5068),
    .C1(_05759_),
    .B1(net8590),
    .A1(net8859),
    .Y(_05760_),
    .A2(\soc_I.kianv_I.datapath_unit_I.Data[1] ));
 sg13g2_nor2_1 _27597_ (.A(net9049),
    .B(_05760_),
    .Y(_01376_));
 sg13g2_nand2b_1 _27598_ (.Y(_05761_),
    .B(net8725),
    .A_N(_11936_));
 sg13g2_a22oi_1 _27599_ (.Y(_05762_),
    .B1(net8588),
    .B2(net4619),
    .A2(\soc_I.kianv_I.datapath_unit_I.Data[2] ),
    .A1(net8857));
 sg13g2_a21oi_1 _27600_ (.A1(_05761_),
    .A2(_05762_),
    .Y(_01377_),
    .B1(net9047));
 sg13g2_nand2b_1 _27601_ (.Y(_05763_),
    .B(net8725),
    .A_N(_12376_));
 sg13g2_a22oi_1 _27602_ (.Y(_05764_),
    .B1(net8588),
    .B2(net4599),
    .A2(\soc_I.kianv_I.datapath_unit_I.Data[3] ),
    .A1(net8857));
 sg13g2_a21oi_1 _27603_ (.A1(_05763_),
    .A2(_05764_),
    .Y(_01378_),
    .B1(net9047));
 sg13g2_nand2_1 _27604_ (.Y(_05765_),
    .A(net8725),
    .B(_12417_));
 sg13g2_a22oi_1 _27605_ (.Y(_05766_),
    .B1(net8587),
    .B2(net4391),
    .A2(\soc_I.kianv_I.datapath_unit_I.Data[4] ),
    .A1(net8856));
 sg13g2_a21oi_1 _27606_ (.A1(_05765_),
    .A2(_05766_),
    .Y(_01379_),
    .B1(net9055));
 sg13g2_nand2b_1 _27607_ (.Y(_05767_),
    .B(net8725),
    .A_N(_12338_));
 sg13g2_a22oi_1 _27608_ (.Y(_05768_),
    .B1(net8587),
    .B2(net4262),
    .A2(\soc_I.kianv_I.datapath_unit_I.Data[5] ),
    .A1(net8856));
 sg13g2_a21oi_1 _27609_ (.A1(_05767_),
    .A2(_05768_),
    .Y(_01380_),
    .B1(net9047));
 sg13g2_nand2b_1 _27610_ (.Y(_05769_),
    .B(net8725),
    .A_N(_11893_));
 sg13g2_a22oi_1 _27611_ (.Y(_05770_),
    .B1(net8587),
    .B2(net4244),
    .A2(\soc_I.kianv_I.datapath_unit_I.Data[6] ),
    .A1(net8856));
 sg13g2_a21oi_1 _27612_ (.A1(_05769_),
    .A2(_05770_),
    .Y(_01381_),
    .B1(net9047));
 sg13g2_a22oi_1 _27613_ (.Y(_05771_),
    .B1(net8590),
    .B2(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[7] ),
    .A2(_12052_),
    .A1(net8724));
 sg13g2_o21ai_1 _27614_ (.B1(_05771_),
    .Y(_05772_),
    .A1(_10855_),
    .A2(_13808_));
 sg13g2_and2_1 _27615_ (.A(net9392),
    .B(_05772_),
    .X(_01382_));
 sg13g2_nand2_1 _27616_ (.Y(_05773_),
    .A(net2913),
    .B(net8587));
 sg13g2_a22oi_1 _27617_ (.Y(_05774_),
    .B1(\soc_I.kianv_I.datapath_unit_I.Data[8] ),
    .B2(net8856),
    .A2(_11914_),
    .A1(net8725));
 sg13g2_a21oi_1 _27618_ (.A1(_05773_),
    .A2(_05774_),
    .Y(_01383_),
    .B1(net9048));
 sg13g2_nand2_1 _27619_ (.Y(_05775_),
    .A(net8725),
    .B(_12360_));
 sg13g2_a22oi_1 _27620_ (.Y(_05776_),
    .B1(net8588),
    .B2(net4441),
    .A2(\soc_I.kianv_I.datapath_unit_I.Data[9] ),
    .A1(net8857));
 sg13g2_a21oi_1 _27621_ (.A1(_05775_),
    .A2(_05776_),
    .Y(_01384_),
    .B1(net9047));
 sg13g2_nand2_1 _27622_ (.Y(_05777_),
    .A(net3590),
    .B(net8587));
 sg13g2_a22oi_1 _27623_ (.Y(_05778_),
    .B1(\soc_I.kianv_I.datapath_unit_I.Data[10] ),
    .B2(net8856),
    .A2(_12069_),
    .A1(net8726));
 sg13g2_a21oi_1 _27624_ (.A1(_05777_),
    .A2(_05778_),
    .Y(_01385_),
    .B1(net9047));
 sg13g2_nand2_1 _27625_ (.Y(_05779_),
    .A(net3951),
    .B(net8585));
 sg13g2_a22oi_1 _27626_ (.Y(_05780_),
    .B1(\soc_I.kianv_I.datapath_unit_I.Data[11] ),
    .B2(net8854),
    .A2(_12026_),
    .A1(net8724));
 sg13g2_a21oi_1 _27627_ (.A1(_05779_),
    .A2(_05780_),
    .Y(_01386_),
    .B1(net9037));
 sg13g2_nand2b_1 _27628_ (.Y(_05781_),
    .B(net8725),
    .A_N(_12438_));
 sg13g2_a22oi_1 _27629_ (.Y(_05782_),
    .B1(net8587),
    .B2(net4223),
    .A2(\soc_I.kianv_I.datapath_unit_I.Data[12] ),
    .A1(net8856));
 sg13g2_a21oi_1 _27630_ (.A1(_05781_),
    .A2(_05782_),
    .Y(_01387_),
    .B1(net9048));
 sg13g2_nand2_1 _27631_ (.Y(_05783_),
    .A(net8726),
    .B(_12451_));
 sg13g2_a22oi_1 _27632_ (.Y(_05784_),
    .B1(net8587),
    .B2(net4466),
    .A2(\soc_I.kianv_I.datapath_unit_I.Data[13] ),
    .A1(net8856));
 sg13g2_a21oi_1 _27633_ (.A1(_05783_),
    .A2(_05784_),
    .Y(_01388_),
    .B1(net9048));
 sg13g2_nand2b_1 _27634_ (.Y(_05785_),
    .B(net8723),
    .A_N(_12273_));
 sg13g2_a22oi_1 _27635_ (.Y(_05786_),
    .B1(net8586),
    .B2(net4064),
    .A2(\soc_I.kianv_I.datapath_unit_I.Data[14] ),
    .A1(net8855));
 sg13g2_a21oi_1 _27636_ (.A1(_05785_),
    .A2(_05786_),
    .Y(_01389_),
    .B1(net9038));
 sg13g2_nand2b_1 _27637_ (.Y(_05787_),
    .B(net8723),
    .A_N(_12252_));
 sg13g2_a22oi_1 _27638_ (.Y(_05788_),
    .B1(net8585),
    .B2(net4787),
    .A2(\soc_I.kianv_I.datapath_unit_I.Data[15] ),
    .A1(net8854));
 sg13g2_a21oi_1 _27639_ (.A1(_05787_),
    .A2(_05788_),
    .Y(_01390_),
    .B1(net9037));
 sg13g2_nand2b_1 _27640_ (.Y(_05789_),
    .B(net8723),
    .A_N(_12427_));
 sg13g2_a22oi_1 _27641_ (.Y(_05790_),
    .B1(net8585),
    .B2(net5156),
    .A2(\soc_I.kianv_I.datapath_unit_I.Data[16] ),
    .A1(net8854));
 sg13g2_a21oi_1 _27642_ (.A1(_05789_),
    .A2(_05790_),
    .Y(_01391_),
    .B1(net9040));
 sg13g2_nand2b_1 _27643_ (.Y(_05791_),
    .B(net8723),
    .A_N(_12349_));
 sg13g2_a22oi_1 _27644_ (.Y(_05792_),
    .B1(net8585),
    .B2(net5285),
    .A2(\soc_I.kianv_I.datapath_unit_I.Data[17] ),
    .A1(net8855));
 sg13g2_a21oi_1 _27645_ (.A1(_05791_),
    .A2(_05792_),
    .Y(_01392_),
    .B1(net9040));
 sg13g2_nand2b_1 _27646_ (.Y(_05793_),
    .B(net8723),
    .A_N(_12285_));
 sg13g2_a22oi_1 _27647_ (.Y(_05794_),
    .B1(net8585),
    .B2(net5173),
    .A2(\soc_I.kianv_I.datapath_unit_I.Data[18] ),
    .A1(net8854));
 sg13g2_a21oi_1 _27648_ (.A1(_05793_),
    .A2(_05794_),
    .Y(_01393_),
    .B1(net9043));
 sg13g2_nand2b_1 _27649_ (.Y(_05795_),
    .B(net8723),
    .A_N(_12389_));
 sg13g2_a22oi_1 _27650_ (.Y(_05796_),
    .B1(net8585),
    .B2(net5100),
    .A2(\soc_I.kianv_I.datapath_unit_I.Data[19] ),
    .A1(net8854));
 sg13g2_a21oi_1 _27651_ (.A1(_05795_),
    .A2(_05796_),
    .Y(_01394_),
    .B1(net9045));
 sg13g2_nand2_1 _27652_ (.Y(_05797_),
    .A(net4256),
    .B(net8588));
 sg13g2_a22oi_1 _27653_ (.Y(_05798_),
    .B1(\soc_I.kianv_I.datapath_unit_I.Data[20] ),
    .B2(net8857),
    .A2(_12180_),
    .A1(net8726));
 sg13g2_a21oi_1 _27654_ (.A1(_05797_),
    .A2(_05798_),
    .Y(_01395_),
    .B1(net9047));
 sg13g2_nand2b_1 _27655_ (.Y(_05799_),
    .B(net8728),
    .A_N(_12399_));
 sg13g2_a22oi_1 _27656_ (.Y(_05800_),
    .B1(net8588),
    .B2(net5099),
    .A2(\soc_I.kianv_I.datapath_unit_I.Data[21] ),
    .A1(net8856));
 sg13g2_a21oi_1 _27657_ (.A1(_05799_),
    .A2(_05800_),
    .Y(_01396_),
    .B1(net9055));
 sg13g2_nand2b_1 _27658_ (.Y(_05801_),
    .B(net8727),
    .A_N(_12263_));
 sg13g2_a22oi_1 _27659_ (.Y(_05802_),
    .B1(net8589),
    .B2(net4923),
    .A2(\soc_I.kianv_I.datapath_unit_I.Data[22] ),
    .A1(net8858));
 sg13g2_a21oi_1 _27660_ (.A1(_05801_),
    .A2(_05802_),
    .Y(_01397_),
    .B1(net9052));
 sg13g2_nand2b_1 _27661_ (.Y(_05803_),
    .B(net8723),
    .A_N(_12320_));
 sg13g2_a22oi_1 _27662_ (.Y(_05804_),
    .B1(net8585),
    .B2(net5206),
    .A2(\soc_I.kianv_I.datapath_unit_I.Data[23] ),
    .A1(net8854));
 sg13g2_a21oi_1 _27663_ (.A1(_05803_),
    .A2(_05804_),
    .Y(_01398_),
    .B1(net9043));
 sg13g2_nand2_1 _27664_ (.Y(_05805_),
    .A(net3538),
    .B(net8587));
 sg13g2_a22oi_1 _27665_ (.Y(_05806_),
    .B1(\soc_I.kianv_I.datapath_unit_I.Data[24] ),
    .B2(net8858),
    .A2(_12095_),
    .A1(net8727));
 sg13g2_a21oi_1 _27666_ (.A1(_05805_),
    .A2(_05806_),
    .Y(_01399_),
    .B1(net9048));
 sg13g2_nand2_1 _27667_ (.Y(_05807_),
    .A(net8727),
    .B(_12136_));
 sg13g2_a22oi_1 _27668_ (.Y(_05808_),
    .B1(net8589),
    .B2(net4846),
    .A2(\soc_I.kianv_I.datapath_unit_I.Data[25] ),
    .A1(net8858));
 sg13g2_a21oi_1 _27669_ (.A1(_05807_),
    .A2(_05808_),
    .Y(_01400_),
    .B1(net9052));
 sg13g2_nand2b_1 _27670_ (.Y(_05809_),
    .B(net8727),
    .A_N(_12240_));
 sg13g2_a22oi_1 _27671_ (.Y(_05810_),
    .B1(net8589),
    .B2(net4965),
    .A2(\soc_I.kianv_I.datapath_unit_I.Data[26] ),
    .A1(net8858));
 sg13g2_a21oi_1 _27672_ (.A1(_05809_),
    .A2(_05810_),
    .Y(_01401_),
    .B1(net9054));
 sg13g2_nand2_2 _27673_ (.Y(_05811_),
    .A(net8728),
    .B(_12225_));
 sg13g2_a22oi_1 _27674_ (.Y(_05812_),
    .B1(net8586),
    .B2(net4613),
    .A2(\soc_I.kianv_I.datapath_unit_I.Data[27] ),
    .A1(net8855));
 sg13g2_a21oi_1 _27675_ (.A1(_05811_),
    .A2(_05812_),
    .Y(_01402_),
    .B1(net9051));
 sg13g2_nand2_1 _27676_ (.Y(_05813_),
    .A(net3786),
    .B(net8588));
 sg13g2_a22oi_1 _27677_ (.Y(_05814_),
    .B1(\soc_I.kianv_I.datapath_unit_I.Data[28] ),
    .B2(net8858),
    .A2(_12162_),
    .A1(net8728));
 sg13g2_a21oi_1 _27678_ (.A1(_05813_),
    .A2(_05814_),
    .Y(_01403_),
    .B1(net9047));
 sg13g2_nand2_1 _27679_ (.Y(_05815_),
    .A(net4606),
    .B(net8589));
 sg13g2_a22oi_1 _27680_ (.Y(_05816_),
    .B1(\soc_I.kianv_I.datapath_unit_I.Data[29] ),
    .B2(net8858),
    .A2(_12310_),
    .A1(net8727));
 sg13g2_a21oi_1 _27681_ (.A1(_05815_),
    .A2(_05816_),
    .Y(_01404_),
    .B1(net9052));
 sg13g2_nand2_1 _27682_ (.Y(_05817_),
    .A(net4076),
    .B(net8586));
 sg13g2_a22oi_1 _27683_ (.Y(_05818_),
    .B1(\soc_I.kianv_I.datapath_unit_I.Data[30] ),
    .B2(net8855),
    .A2(_11982_),
    .A1(net8724));
 sg13g2_a21oi_1 _27684_ (.A1(_05817_),
    .A2(_05818_),
    .Y(_01405_),
    .B1(net9045));
 sg13g2_nand2_1 _27685_ (.Y(_05819_),
    .A(net4682),
    .B(net8585));
 sg13g2_a22oi_1 _27686_ (.Y(_05820_),
    .B1(\soc_I.kianv_I.datapath_unit_I.Data[31] ),
    .B2(net8854),
    .A2(_12210_),
    .A1(net8723));
 sg13g2_a21oi_1 _27687_ (.A1(_05819_),
    .A2(_05820_),
    .Y(_01406_),
    .B1(net9040));
 sg13g2_o21ai_1 _27688_ (.B1(net9397),
    .Y(_05821_),
    .A1(net4597),
    .A2(net7472));
 sg13g2_a21oi_1 _27689_ (.A1(_11729_),
    .A2(net7472),
    .Y(_01407_),
    .B1(_05821_));
 sg13g2_o21ai_1 _27690_ (.B1(net9406),
    .Y(_05822_),
    .A1(net5056),
    .A2(net7475));
 sg13g2_a21oi_1 _27691_ (.A1(_11837_),
    .A2(net7475),
    .Y(_01408_),
    .B1(_05822_));
 sg13g2_o21ai_1 _27692_ (.B1(net9405),
    .Y(_05823_),
    .A1(net4543),
    .A2(net7475));
 sg13g2_a21oi_1 _27693_ (.A1(_11936_),
    .A2(net7475),
    .Y(_01409_),
    .B1(_05823_));
 sg13g2_o21ai_1 _27694_ (.B1(net9409),
    .Y(_05824_),
    .A1(net4805),
    .A2(net7473));
 sg13g2_a21oi_1 _27695_ (.A1(_12376_),
    .A2(net7473),
    .Y(_01410_),
    .B1(_05824_));
 sg13g2_o21ai_1 _27696_ (.B1(net9408),
    .Y(_05825_),
    .A1(net4336),
    .A2(net7474));
 sg13g2_a21oi_1 _27697_ (.A1(_12416_),
    .A2(net7474),
    .Y(_01411_),
    .B1(_05825_));
 sg13g2_o21ai_1 _27698_ (.B1(net9396),
    .Y(_05826_),
    .A1(net4469),
    .A2(net7474));
 sg13g2_a21oi_1 _27699_ (.A1(_12338_),
    .A2(net7474),
    .Y(_01412_),
    .B1(_05826_));
 sg13g2_o21ai_1 _27700_ (.B1(net9408),
    .Y(_05827_),
    .A1(net4699),
    .A2(net7473));
 sg13g2_a21oi_1 _27701_ (.A1(_11893_),
    .A2(net7473),
    .Y(_01413_),
    .B1(_05827_));
 sg13g2_o21ai_1 _27702_ (.B1(net9396),
    .Y(_05828_),
    .A1(net4197),
    .A2(net7477));
 sg13g2_a21oi_1 _27703_ (.A1(_12051_),
    .A2(net7477),
    .Y(_01414_),
    .B1(_05828_));
 sg13g2_o21ai_1 _27704_ (.B1(net9409),
    .Y(_05829_),
    .A1(_11914_),
    .A2(net7481));
 sg13g2_a21oi_1 _27705_ (.A1(_10506_),
    .A2(net7481),
    .Y(_01415_),
    .B1(_05829_));
 sg13g2_o21ai_1 _27706_ (.B1(net9408),
    .Y(_05830_),
    .A1(_12360_),
    .A2(net7481));
 sg13g2_a21oi_1 _27707_ (.A1(_10505_),
    .A2(net7481),
    .Y(_01416_),
    .B1(_05830_));
 sg13g2_o21ai_1 _27708_ (.B1(net9413),
    .Y(_05831_),
    .A1(net4609),
    .A2(net7474));
 sg13g2_a21oi_1 _27709_ (.A1(_12068_),
    .A2(net7474),
    .Y(_01417_),
    .B1(_05831_));
 sg13g2_o21ai_1 _27710_ (.B1(net9373),
    .Y(_05832_),
    .A1(_12026_),
    .A2(net7484));
 sg13g2_a21oi_1 _27711_ (.A1(_10504_),
    .A2(net7484),
    .Y(_01418_),
    .B1(_05832_));
 sg13g2_o21ai_1 _27712_ (.B1(net9408),
    .Y(_05833_),
    .A1(net4934),
    .A2(net7473));
 sg13g2_a21oi_1 _27713_ (.A1(_12438_),
    .A2(net7473),
    .Y(_01419_),
    .B1(_05833_));
 sg13g2_o21ai_1 _27714_ (.B1(net9413),
    .Y(_05834_),
    .A1(net4792),
    .A2(net7473));
 sg13g2_a21oi_1 _27715_ (.A1(_12450_),
    .A2(net7473),
    .Y(_01420_),
    .B1(_05834_));
 sg13g2_o21ai_1 _27716_ (.B1(net9386),
    .Y(_05835_),
    .A1(net4272),
    .A2(net7478));
 sg13g2_a21oi_1 _27717_ (.A1(_12273_),
    .A2(net7472),
    .Y(_01421_),
    .B1(_05835_));
 sg13g2_o21ai_1 _27718_ (.B1(net9381),
    .Y(_05836_),
    .A1(net4449),
    .A2(net7471));
 sg13g2_a21oi_1 _27719_ (.A1(_12252_),
    .A2(net7471),
    .Y(_01422_),
    .B1(_05836_));
 sg13g2_o21ai_1 _27720_ (.B1(net9381),
    .Y(_05837_),
    .A1(net4750),
    .A2(net7471));
 sg13g2_a21oi_1 _27721_ (.A1(_12427_),
    .A2(net7471),
    .Y(_01423_),
    .B1(_05837_));
 sg13g2_o21ai_1 _27722_ (.B1(net9381),
    .Y(_05838_),
    .A1(net4380),
    .A2(net7471));
 sg13g2_a21oi_1 _27723_ (.A1(_12349_),
    .A2(net7471),
    .Y(_01424_),
    .B1(_05838_));
 sg13g2_o21ai_1 _27724_ (.B1(net9381),
    .Y(_05839_),
    .A1(net4570),
    .A2(net7472));
 sg13g2_a21oi_1 _27725_ (.A1(_12285_),
    .A2(net7472),
    .Y(_01425_),
    .B1(_05839_));
 sg13g2_o21ai_1 _27726_ (.B1(net9386),
    .Y(_05840_),
    .A1(net4235),
    .A2(net7478));
 sg13g2_a21oi_1 _27727_ (.A1(_12389_),
    .A2(net7472),
    .Y(_01426_),
    .B1(_05840_));
 sg13g2_o21ai_1 _27728_ (.B1(net9410),
    .Y(_05841_),
    .A1(net4266),
    .A2(net7475));
 sg13g2_a21oi_1 _27729_ (.A1(_12179_),
    .A2(net7475),
    .Y(_01427_),
    .B1(_05841_));
 sg13g2_o21ai_1 _27730_ (.B1(net9411),
    .Y(_05842_),
    .A1(net4683),
    .A2(net7476));
 sg13g2_a21oi_1 _27731_ (.A1(_12399_),
    .A2(net7476),
    .Y(_01428_),
    .B1(_05842_));
 sg13g2_o21ai_1 _27732_ (.B1(net9410),
    .Y(_05843_),
    .A1(net4811),
    .A2(net7476));
 sg13g2_a21oi_1 _27733_ (.A1(_12263_),
    .A2(net7476),
    .Y(_01429_),
    .B1(_05843_));
 sg13g2_o21ai_1 _27734_ (.B1(net9387),
    .Y(_05844_),
    .A1(net4604),
    .A2(net7471));
 sg13g2_a21oi_1 _27735_ (.A1(_12320_),
    .A2(net7471),
    .Y(_01430_),
    .B1(_05844_));
 sg13g2_o21ai_1 _27736_ (.B1(net9405),
    .Y(_05845_),
    .A1(_12095_),
    .A2(net7481));
 sg13g2_a21oi_1 _27737_ (.A1(_10503_),
    .A2(net7482),
    .Y(_01431_),
    .B1(_05845_));
 sg13g2_o21ai_1 _27738_ (.B1(net9410),
    .Y(_05846_),
    .A1(_12136_),
    .A2(net7482));
 sg13g2_a21oi_1 _27739_ (.A1(_10502_),
    .A2(net7481),
    .Y(_01432_),
    .B1(_05846_));
 sg13g2_o21ai_1 _27740_ (.B1(net9410),
    .Y(_05847_),
    .A1(net4703),
    .A2(net7475));
 sg13g2_a21oi_1 _27741_ (.A1(_12240_),
    .A2(net7475),
    .Y(_01433_),
    .B1(_05847_));
 sg13g2_o21ai_1 _27742_ (.B1(net9401),
    .Y(_05848_),
    .A1(_12225_),
    .A2(net7483));
 sg13g2_a21oi_1 _27743_ (.A1(_10501_),
    .A2(net7483),
    .Y(_01434_),
    .B1(_05848_));
 sg13g2_o21ai_1 _27744_ (.B1(net9404),
    .Y(_05849_),
    .A1(_12162_),
    .A2(net7482));
 sg13g2_a21oi_1 _27745_ (.A1(_10500_),
    .A2(net7481),
    .Y(_01435_),
    .B1(_05849_));
 sg13g2_o21ai_1 _27746_ (.B1(net9405),
    .Y(_05850_),
    .A1(_12310_),
    .A2(net7481));
 sg13g2_a21oi_1 _27747_ (.A1(_10499_),
    .A2(net7482),
    .Y(_01436_),
    .B1(_05850_));
 sg13g2_o21ai_1 _27748_ (.B1(net9386),
    .Y(_05851_),
    .A1(_11982_),
    .A2(net7484));
 sg13g2_a21oi_1 _27749_ (.A1(_10498_),
    .A2(net7484),
    .Y(_01437_),
    .B1(_05851_));
 sg13g2_o21ai_1 _27750_ (.B1(net9386),
    .Y(_05852_),
    .A1(_12210_),
    .A2(net7484));
 sg13g2_a21oi_1 _27751_ (.A1(_10497_),
    .A2(net7484),
    .Y(_01438_),
    .B1(_05852_));
 sg13g2_nor2b_2 _27752_ (.A(_04650_),
    .B_N(_10867_),
    .Y(_05853_));
 sg13g2_o21ai_1 _27753_ (.B1(_10867_),
    .Y(_05854_),
    .A1(_10596_),
    .A2(_13283_));
 sg13g2_o21ai_1 _27754_ (.B1(net9386),
    .Y(_05855_),
    .A1(net4800),
    .A2(net7369));
 sg13g2_a21oi_1 _27755_ (.A1(_10496_),
    .A2(net7369),
    .Y(_01439_),
    .B1(_05855_));
 sg13g2_o21ai_1 _27756_ (.B1(net9377),
    .Y(_05856_),
    .A1(\soc_I.PC[1] ),
    .A2(net7367));
 sg13g2_a21oi_1 _27757_ (.A1(_10495_),
    .A2(net7367),
    .Y(_01440_),
    .B1(_05856_));
 sg13g2_o21ai_1 _27758_ (.B1(net9392),
    .Y(_05857_),
    .A1(\soc_I.PC[2] ),
    .A2(net7368));
 sg13g2_a21oi_1 _27759_ (.A1(_10494_),
    .A2(net7368),
    .Y(_01441_),
    .B1(_05857_));
 sg13g2_o21ai_1 _27760_ (.B1(net9378),
    .Y(_05858_),
    .A1(net4241),
    .A2(net7367));
 sg13g2_a21oi_1 _27761_ (.A1(_10493_),
    .A2(net7367),
    .Y(_01442_),
    .B1(_05858_));
 sg13g2_o21ai_1 _27762_ (.B1(net9394),
    .Y(_05859_),
    .A1(\soc_I.PC[4] ),
    .A2(net7371));
 sg13g2_a21oi_1 _27763_ (.A1(_10492_),
    .A2(net7374),
    .Y(_01443_),
    .B1(_05859_));
 sg13g2_o21ai_1 _27764_ (.B1(net9393),
    .Y(_05860_),
    .A1(\soc_I.PC[5] ),
    .A2(net7371));
 sg13g2_a21oi_1 _27765_ (.A1(_10491_),
    .A2(net7371),
    .Y(_01444_),
    .B1(_05860_));
 sg13g2_o21ai_1 _27766_ (.B1(net9393),
    .Y(_05861_),
    .A1(\soc_I.PC[6] ),
    .A2(net7371));
 sg13g2_a21oi_1 _27767_ (.A1(_10490_),
    .A2(net7371),
    .Y(_01445_),
    .B1(_05861_));
 sg13g2_o21ai_1 _27768_ (.B1(net9346),
    .Y(_05862_),
    .A1(\soc_I.PC[7] ),
    .A2(net7365));
 sg13g2_a21oi_1 _27769_ (.A1(_10489_),
    .A2(net7365),
    .Y(_01446_),
    .B1(_05862_));
 sg13g2_o21ai_1 _27770_ (.B1(net9376),
    .Y(_05863_),
    .A1(\soc_I.PC[8] ),
    .A2(net7368));
 sg13g2_a21oi_1 _27771_ (.A1(_10488_),
    .A2(net7368),
    .Y(_01447_),
    .B1(_05863_));
 sg13g2_o21ai_1 _27772_ (.B1(net9394),
    .Y(_05864_),
    .A1(\soc_I.PC[9] ),
    .A2(net7371));
 sg13g2_a21oi_1 _27773_ (.A1(_10487_),
    .A2(net7371),
    .Y(_01448_),
    .B1(_05864_));
 sg13g2_o21ai_1 _27774_ (.B1(net9349),
    .Y(_05865_),
    .A1(net5441),
    .A2(net7365));
 sg13g2_a21oi_1 _27775_ (.A1(_10486_),
    .A2(net7365),
    .Y(_01449_),
    .B1(_05865_));
 sg13g2_o21ai_1 _27776_ (.B1(net9347),
    .Y(_05866_),
    .A1(\soc_I.PC[11] ),
    .A2(net7365));
 sg13g2_a21oi_1 _27777_ (.A1(_10485_),
    .A2(net7365),
    .Y(_01450_),
    .B1(_05866_));
 sg13g2_o21ai_1 _27778_ (.B1(net9376),
    .Y(_05867_),
    .A1(\soc_I.PC[12] ),
    .A2(net7368));
 sg13g2_a21oi_1 _27779_ (.A1(_10484_),
    .A2(net7368),
    .Y(_01451_),
    .B1(_05867_));
 sg13g2_o21ai_1 _27780_ (.B1(net9406),
    .Y(_05868_),
    .A1(net5385),
    .A2(net7373));
 sg13g2_a21oi_1 _27781_ (.A1(_10483_),
    .A2(net7373),
    .Y(_01452_),
    .B1(_05868_));
 sg13g2_o21ai_1 _27782_ (.B1(net9381),
    .Y(_05869_),
    .A1(net4664),
    .A2(net7366));
 sg13g2_a21oi_1 _27783_ (.A1(_10482_),
    .A2(net7366),
    .Y(_01453_),
    .B1(_05869_));
 sg13g2_o21ai_1 _27784_ (.B1(net9355),
    .Y(_05870_),
    .A1(\soc_I.PC[15] ),
    .A2(net7366));
 sg13g2_a21oi_1 _27785_ (.A1(_10481_),
    .A2(net7366),
    .Y(_01454_),
    .B1(_05870_));
 sg13g2_o21ai_1 _27786_ (.B1(net9343),
    .Y(_05871_),
    .A1(\soc_I.kianv_I.datapath_unit_I.OldPC[16] ),
    .A2(net7349));
 sg13g2_a21oi_1 _27787_ (.A1(_10457_),
    .A2(net7349),
    .Y(_01455_),
    .B1(_05871_));
 sg13g2_o21ai_1 _27788_ (.B1(net9343),
    .Y(_05872_),
    .A1(net5307),
    .A2(net7349));
 sg13g2_a21oi_1 _27789_ (.A1(_10456_),
    .A2(net7348),
    .Y(_01456_),
    .B1(_05872_));
 sg13g2_o21ai_1 _27790_ (.B1(net9343),
    .Y(_05873_),
    .A1(\soc_I.kianv_I.datapath_unit_I.OldPC[18] ),
    .A2(net7348));
 sg13g2_a21oi_1 _27791_ (.A1(_10455_),
    .A2(net7348),
    .Y(_01457_),
    .B1(_05873_));
 sg13g2_o21ai_1 _27792_ (.B1(net9359),
    .Y(_05874_),
    .A1(\soc_I.kianv_I.datapath_unit_I.OldPC[19] ),
    .A2(net7349));
 sg13g2_a21oi_1 _27793_ (.A1(_10454_),
    .A2(net7348),
    .Y(_01458_),
    .B1(_05874_));
 sg13g2_a21oi_1 _27794_ (.A1(net5404),
    .A2(net7370),
    .Y(_05875_),
    .B1(net9045));
 sg13g2_o21ai_1 _27795_ (.B1(_05875_),
    .Y(_01459_),
    .A1(_10453_),
    .A2(net7370));
 sg13g2_o21ai_1 _27796_ (.B1(net9404),
    .Y(_05876_),
    .A1(\soc_I.PC[21] ),
    .A2(net7372));
 sg13g2_a21oi_1 _27797_ (.A1(_10480_),
    .A2(net7373),
    .Y(_01460_),
    .B1(_05876_));
 sg13g2_o21ai_1 _27798_ (.B1(net9404),
    .Y(_05877_),
    .A1(\soc_I.PC[22] ),
    .A2(net7372));
 sg13g2_a21oi_1 _27799_ (.A1(_10479_),
    .A2(net7372),
    .Y(_01461_),
    .B1(_05877_));
 sg13g2_o21ai_1 _27800_ (.B1(net9387),
    .Y(_05878_),
    .A1(\soc_I.PC[23] ),
    .A2(net7370));
 sg13g2_a21oi_1 _27801_ (.A1(_10478_),
    .A2(net7370),
    .Y(_01462_),
    .B1(_05878_));
 sg13g2_o21ai_1 _27802_ (.B1(net9401),
    .Y(_05879_),
    .A1(\soc_I.PC[24] ),
    .A2(net7372));
 sg13g2_a21oi_1 _27803_ (.A1(_10477_),
    .A2(net7372),
    .Y(_01463_),
    .B1(_05879_));
 sg13g2_o21ai_1 _27804_ (.B1(net9404),
    .Y(_05880_),
    .A1(\soc_I.PC[25] ),
    .A2(net7373));
 sg13g2_a21oi_1 _27805_ (.A1(_10476_),
    .A2(net7372),
    .Y(_01464_),
    .B1(_05880_));
 sg13g2_o21ai_1 _27806_ (.B1(net9404),
    .Y(_05881_),
    .A1(\soc_I.PC[26] ),
    .A2(net7372));
 sg13g2_a21oi_1 _27807_ (.A1(_10475_),
    .A2(net7372),
    .Y(_01465_),
    .B1(_05881_));
 sg13g2_o21ai_1 _27808_ (.B1(net9389),
    .Y(_05882_),
    .A1(\soc_I.PC[27] ),
    .A2(net7370));
 sg13g2_a21oi_1 _27809_ (.A1(_10474_),
    .A2(net7375),
    .Y(_01466_),
    .B1(_05882_));
 sg13g2_o21ai_1 _27810_ (.B1(net9387),
    .Y(_05883_),
    .A1(\soc_I.PC[28] ),
    .A2(net7370));
 sg13g2_a21oi_1 _27811_ (.A1(_10473_),
    .A2(net7370),
    .Y(_01467_),
    .B1(_05883_));
 sg13g2_a21oi_1 _27812_ (.A1(\soc_I.kianv_I.datapath_unit_I.OldPC[29] ),
    .A2(net7366),
    .Y(_05884_),
    .B1(net9040));
 sg13g2_o21ai_1 _27813_ (.B1(_05884_),
    .Y(_01468_),
    .A1(_10452_),
    .A2(net7366));
 sg13g2_o21ai_1 _27814_ (.B1(net9382),
    .Y(_05885_),
    .A1(\soc_I.kianv_I.datapath_unit_I.OldPC[30] ),
    .A2(net7360));
 sg13g2_a21oi_1 _27815_ (.A1(_10451_),
    .A2(net7360),
    .Y(_01469_),
    .B1(_05885_));
 sg13g2_o21ai_1 _27816_ (.B1(net9356),
    .Y(_05886_),
    .A1(\soc_I.kianv_I.datapath_unit_I.OldPC[31] ),
    .A2(net7348));
 sg13g2_a21oi_1 _27817_ (.A1(_10450_),
    .A2(net7348),
    .Y(_01470_),
    .B1(_05886_));
 sg13g2_nor3_2 _27818_ (.A(net8977),
    .B(_10847_),
    .C(_10849_),
    .Y(_05887_));
 sg13g2_o21ai_1 _27819_ (.B1(net9398),
    .Y(_05888_),
    .A1(net4795),
    .A2(_05887_));
 sg13g2_nor2_1 _27820_ (.A(_10851_),
    .B(_05888_),
    .Y(_01471_));
 sg13g2_o21ai_1 _27821_ (.B1(net9397),
    .Y(_05889_),
    .A1(net4719),
    .A2(net8846));
 sg13g2_a21oi_1 _27822_ (.A1(net8846),
    .A2(_11729_),
    .Y(_01472_),
    .B1(_05889_));
 sg13g2_o21ai_1 _27823_ (.B1(net9406),
    .Y(_05890_),
    .A1(net4642),
    .A2(net8851));
 sg13g2_a21oi_1 _27824_ (.A1(net8851),
    .A2(_11837_),
    .Y(_01473_),
    .B1(_05890_));
 sg13g2_o21ai_1 _27825_ (.B1(net9405),
    .Y(_05891_),
    .A1(net4411),
    .A2(net8850));
 sg13g2_a21oi_1 _27826_ (.A1(net8850),
    .A2(_11936_),
    .Y(_01474_),
    .B1(_05891_));
 sg13g2_o21ai_1 _27827_ (.B1(net9409),
    .Y(_05892_),
    .A1(net4812),
    .A2(net8847));
 sg13g2_a21oi_1 _27828_ (.A1(net8847),
    .A2(_12376_),
    .Y(_01475_),
    .B1(_05892_));
 sg13g2_o21ai_1 _27829_ (.B1(net9408),
    .Y(_05893_),
    .A1(net4359),
    .A2(net8848));
 sg13g2_a21oi_1 _27830_ (.A1(net8848),
    .A2(_12416_),
    .Y(_01476_),
    .B1(_05893_));
 sg13g2_o21ai_1 _27831_ (.B1(net9408),
    .Y(_05894_),
    .A1(net4384),
    .A2(net8848));
 sg13g2_a21oi_1 _27832_ (.A1(net8848),
    .A2(_12338_),
    .Y(_01477_),
    .B1(_05894_));
 sg13g2_o21ai_1 _27833_ (.B1(net9409),
    .Y(_05895_),
    .A1(net4568),
    .A2(net8847));
 sg13g2_a21oi_1 _27834_ (.A1(net8847),
    .A2(_11893_),
    .Y(_01478_),
    .B1(_05895_));
 sg13g2_o21ai_1 _27835_ (.B1(net9396),
    .Y(_05896_),
    .A1(net4393),
    .A2(net8849));
 sg13g2_a21oi_1 _27836_ (.A1(net8849),
    .A2(_12051_),
    .Y(_01479_),
    .B1(_05896_));
 sg13g2_nor2_1 _27837_ (.A(net8843),
    .B(_11914_),
    .Y(_05897_));
 sg13g2_o21ai_1 _27838_ (.B1(net9408),
    .Y(_05898_),
    .A1(net4898),
    .A2(net8848));
 sg13g2_nor2_1 _27839_ (.A(_05897_),
    .B(_05898_),
    .Y(_01480_));
 sg13g2_nor2_1 _27840_ (.A(net8843),
    .B(_12360_),
    .Y(_05899_));
 sg13g2_o21ai_1 _27841_ (.B1(net9408),
    .Y(_05900_),
    .A1(net4621),
    .A2(net8848));
 sg13g2_nor2_1 _27842_ (.A(_05899_),
    .B(_05900_),
    .Y(_01481_));
 sg13g2_o21ai_1 _27843_ (.B1(net9409),
    .Y(_05901_),
    .A1(net4693),
    .A2(net8847));
 sg13g2_a21oi_1 _27844_ (.A1(net8847),
    .A2(_12068_),
    .Y(_01482_),
    .B1(_05901_));
 sg13g2_nor2_1 _27845_ (.A(net8842),
    .B(_12026_),
    .Y(_05902_));
 sg13g2_o21ai_1 _27846_ (.B1(net9392),
    .Y(_05903_),
    .A1(net4706),
    .A2(net8853));
 sg13g2_nor2_1 _27847_ (.A(_05902_),
    .B(_05903_),
    .Y(_01483_));
 sg13g2_o21ai_1 _27848_ (.B1(net9409),
    .Y(_05904_),
    .A1(net4622),
    .A2(net8847));
 sg13g2_a21oi_1 _27849_ (.A1(net8847),
    .A2(_12438_),
    .Y(_01484_),
    .B1(_05904_));
 sg13g2_o21ai_1 _27850_ (.B1(net9409),
    .Y(_05905_),
    .A1(net4458),
    .A2(net8849));
 sg13g2_a21oi_1 _27851_ (.A1(net8848),
    .A2(_12450_),
    .Y(_01485_),
    .B1(_05905_));
 sg13g2_o21ai_1 _27852_ (.B1(net9399),
    .Y(_05906_),
    .A1(net4625),
    .A2(net8846));
 sg13g2_a21oi_1 _27853_ (.A1(net8846),
    .A2(_12273_),
    .Y(_01486_),
    .B1(_05906_));
 sg13g2_o21ai_1 _27854_ (.B1(net9386),
    .Y(_05907_),
    .A1(net4315),
    .A2(net8844));
 sg13g2_a21oi_1 _27855_ (.A1(net8844),
    .A2(_12252_),
    .Y(_01487_),
    .B1(_05907_));
 sg13g2_o21ai_1 _27856_ (.B1(net9397),
    .Y(_05908_),
    .A1(net4486),
    .A2(net8844));
 sg13g2_a21oi_1 _27857_ (.A1(net8844),
    .A2(_12427_),
    .Y(_01488_),
    .B1(_05908_));
 sg13g2_o21ai_1 _27858_ (.B1(net9397),
    .Y(_05909_),
    .A1(net4410),
    .A2(net8844));
 sg13g2_a21oi_1 _27859_ (.A1(net8844),
    .A2(_12349_),
    .Y(_01489_),
    .B1(_05909_));
 sg13g2_o21ai_1 _27860_ (.B1(net9399),
    .Y(_05910_),
    .A1(net4533),
    .A2(net8845));
 sg13g2_a21oi_1 _27861_ (.A1(net8844),
    .A2(_12285_),
    .Y(_01490_),
    .B1(_05910_));
 sg13g2_o21ai_1 _27862_ (.B1(net9399),
    .Y(_05911_),
    .A1(net4372),
    .A2(net8845));
 sg13g2_a21oi_1 _27863_ (.A1(net8845),
    .A2(_12389_),
    .Y(_01491_),
    .B1(_05911_));
 sg13g2_o21ai_1 _27864_ (.B1(net9410),
    .Y(_05912_),
    .A1(net4626),
    .A2(net8852));
 sg13g2_a21oi_1 _27865_ (.A1(net8852),
    .A2(_12179_),
    .Y(_01492_),
    .B1(_05912_));
 sg13g2_o21ai_1 _27866_ (.B1(net9411),
    .Y(_05913_),
    .A1(net4348),
    .A2(net8853));
 sg13g2_a21oi_1 _27867_ (.A1(net8852),
    .A2(_12399_),
    .Y(_01493_),
    .B1(_05913_));
 sg13g2_o21ai_1 _27868_ (.B1(net9410),
    .Y(_05914_),
    .A1(net4470),
    .A2(net8852));
 sg13g2_a21oi_1 _27869_ (.A1(net8852),
    .A2(_12263_),
    .Y(_01494_),
    .B1(_05914_));
 sg13g2_o21ai_1 _27870_ (.B1(net9405),
    .Y(_05915_),
    .A1(net4379),
    .A2(net8850));
 sg13g2_a21oi_1 _27871_ (.A1(net8850),
    .A2(_12320_),
    .Y(_01495_),
    .B1(_05915_));
 sg13g2_nor2_1 _27872_ (.A(net8842),
    .B(_12095_),
    .Y(_05916_));
 sg13g2_o21ai_1 _27873_ (.B1(net9405),
    .Y(_05917_),
    .A1(net4614),
    .A2(net8850));
 sg13g2_nor2_1 _27874_ (.A(_05916_),
    .B(_05917_),
    .Y(_01496_));
 sg13g2_nor2_1 _27875_ (.A(net8842),
    .B(_12136_),
    .Y(_05918_));
 sg13g2_o21ai_1 _27876_ (.B1(net9411),
    .Y(_05919_),
    .A1(net4431),
    .A2(net8851));
 sg13g2_nor2_1 _27877_ (.A(_05918_),
    .B(_05919_),
    .Y(_01497_));
 sg13g2_o21ai_1 _27878_ (.B1(net9410),
    .Y(_05920_),
    .A1(net4601),
    .A2(net8852));
 sg13g2_a21oi_1 _27879_ (.A1(net8852),
    .A2(_12240_),
    .Y(_01498_),
    .B1(_05920_));
 sg13g2_nor2_1 _27880_ (.A(net8843),
    .B(_12225_),
    .Y(_05921_));
 sg13g2_o21ai_1 _27881_ (.B1(net9405),
    .Y(_05922_),
    .A1(net4618),
    .A2(net8850));
 sg13g2_nor2_1 _27882_ (.A(_05921_),
    .B(_05922_),
    .Y(_01499_));
 sg13g2_nor2_1 _27883_ (.A(net8843),
    .B(_12162_),
    .Y(_05923_));
 sg13g2_o21ai_1 _27884_ (.B1(net9405),
    .Y(_05924_),
    .A1(net4596),
    .A2(net8850));
 sg13g2_nor2_1 _27885_ (.A(_05923_),
    .B(_05924_),
    .Y(_01500_));
 sg13g2_nor2_1 _27886_ (.A(net8842),
    .B(_12310_),
    .Y(_05925_));
 sg13g2_o21ai_1 _27887_ (.B1(net9410),
    .Y(_05926_),
    .A1(net4381),
    .A2(net8850));
 sg13g2_nor2_1 _27888_ (.A(_05925_),
    .B(_05926_),
    .Y(_01501_));
 sg13g2_nor2_1 _27889_ (.A(net8842),
    .B(_11982_),
    .Y(_05927_));
 sg13g2_o21ai_1 _27890_ (.B1(net9389),
    .Y(_05928_),
    .A1(net4437),
    .A2(net8845));
 sg13g2_nor2_1 _27891_ (.A(_05927_),
    .B(_05928_),
    .Y(_01502_));
 sg13g2_nor2_1 _27892_ (.A(net8842),
    .B(_12210_),
    .Y(_05929_));
 sg13g2_o21ai_1 _27893_ (.B1(net9397),
    .Y(_05930_),
    .A1(net4544),
    .A2(net8844));
 sg13g2_nor2_1 _27894_ (.A(_05929_),
    .B(_05930_),
    .Y(_01503_));
 sg13g2_a21oi_1 _27895_ (.A1(_13287_),
    .A2(net7351),
    .Y(_05931_),
    .B1(net9038));
 sg13g2_o21ai_1 _27896_ (.B1(_05931_),
    .Y(_01504_),
    .A1(_10472_),
    .A2(net7351));
 sg13g2_a21oi_1 _27897_ (.A1(_13377_),
    .A2(net7351),
    .Y(_05932_),
    .B1(net9039));
 sg13g2_o21ai_1 _27898_ (.B1(_05932_),
    .Y(_01505_),
    .A1(_10471_),
    .A2(net7352));
 sg13g2_o21ai_1 _27899_ (.B1(net9377),
    .Y(_05933_),
    .A1(net5542),
    .A2(net7352));
 sg13g2_a21oi_1 _27900_ (.A1(_13439_),
    .A2(net7351),
    .Y(_01506_),
    .B1(_05933_));
 sg13g2_o21ai_1 _27901_ (.B1(net9377),
    .Y(_05934_),
    .A1(net4952),
    .A2(net7352));
 sg13g2_a21oi_1 _27902_ (.A1(_13506_),
    .A2(net7352),
    .Y(_01507_),
    .B1(_05934_));
 sg13g2_a21oi_1 _27903_ (.A1(_13571_),
    .A2(net7354),
    .Y(_05935_),
    .B1(net9037));
 sg13g2_o21ai_1 _27904_ (.B1(_05935_),
    .Y(_01508_),
    .A1(_10469_),
    .A2(net7357));
 sg13g2_o21ai_1 _27905_ (.B1(net9392),
    .Y(_05936_),
    .A1(net9714),
    .A2(net7355));
 sg13g2_a21oi_1 _27906_ (.A1(_13634_),
    .A2(net7355),
    .Y(_01509_),
    .B1(_05936_));
 sg13g2_o21ai_1 _27907_ (.B1(net9397),
    .Y(_05937_),
    .A1(net9712),
    .A2(net7356));
 sg13g2_a21oi_1 _27908_ (.A1(_13702_),
    .A2(net7355),
    .Y(_01510_),
    .B1(_05937_));
 sg13g2_o21ai_1 _27909_ (.B1(net9378),
    .Y(_05938_),
    .A1(_13768_),
    .A2(net7367));
 sg13g2_a21oi_1 _27910_ (.A1(_10468_),
    .A2(net7374),
    .Y(_01511_),
    .B1(_05938_));
 sg13g2_o21ai_1 _27911_ (.B1(net9373),
    .Y(_05939_),
    .A1(net5556),
    .A2(net7354));
 sg13g2_a21oi_1 _27912_ (.A1(_13317_),
    .A2(net7354),
    .Y(_01512_),
    .B1(_05939_));
 sg13g2_o21ai_1 _27913_ (.B1(net9394),
    .Y(_05940_),
    .A1(net5539),
    .A2(net7358));
 sg13g2_a21oi_1 _27914_ (.A1(_13397_),
    .A2(net7358),
    .Y(_01513_),
    .B1(_05940_));
 sg13g2_o21ai_1 _27915_ (.B1(net9376),
    .Y(_05941_),
    .A1(net5054),
    .A2(net7351));
 sg13g2_a21oi_1 _27916_ (.A1(_13461_),
    .A2(net7351),
    .Y(_01514_),
    .B1(_05941_));
 sg13g2_o21ai_1 _27917_ (.B1(net9376),
    .Y(_05942_),
    .A1(net9709),
    .A2(net7351));
 sg13g2_a21oi_1 _27918_ (.A1(_13527_),
    .A2(net7351),
    .Y(_01515_),
    .B1(_05942_));
 sg13g2_o21ai_1 _27919_ (.B1(net9382),
    .Y(_05943_),
    .A1(net9707),
    .A2(net7350));
 sg13g2_a21oi_2 _27920_ (.B1(_05943_),
    .Y(_01516_),
    .A2(net7350),
    .A1(_13591_));
 sg13g2_o21ai_1 _27921_ (.B1(net9347),
    .Y(_05944_),
    .A1(net9700),
    .A2(net7348));
 sg13g2_a21oi_1 _27922_ (.A1(_13668_),
    .A2(net7348),
    .Y(_01517_),
    .B1(_05944_));
 sg13g2_o21ai_1 _27923_ (.B1(net9386),
    .Y(_05945_),
    .A1(net9699),
    .A2(net7353));
 sg13g2_a21oi_1 _27924_ (.A1(_13724_),
    .A2(net7353),
    .Y(_01518_),
    .B1(_05945_));
 sg13g2_o21ai_1 _27925_ (.B1(net9346),
    .Y(_05946_),
    .A1(_13787_),
    .A2(net7365));
 sg13g2_a21oi_1 _27926_ (.A1(net9084),
    .A2(net7365),
    .Y(_01519_),
    .B1(_05946_));
 sg13g2_o21ai_1 _27927_ (.B1(net9375),
    .Y(_05947_),
    .A1(net9601),
    .A2(net7354));
 sg13g2_a21oi_1 _27928_ (.A1(_13340_),
    .A2(net7354),
    .Y(_01520_),
    .B1(_05947_));
 sg13g2_o21ai_1 _27929_ (.B1(net9378),
    .Y(_05948_),
    .A1(_13409_),
    .A2(net7367));
 sg13g2_a21oi_2 _27930_ (.B1(_05948_),
    .Y(_01521_),
    .A2(net7367),
    .A1(net9110));
 sg13g2_o21ai_1 _27931_ (.B1(net9350),
    .Y(_05949_),
    .A1(net9554),
    .A2(net7350));
 sg13g2_a21oi_1 _27932_ (.A1(_13473_),
    .A2(net7350),
    .Y(_01522_),
    .B1(_05949_));
 sg13g2_o21ai_1 _27933_ (.B1(net9378),
    .Y(_05950_),
    .A1(_13538_),
    .A2(net7367));
 sg13g2_a21oi_1 _27934_ (.A1(net9112),
    .A2(net7368),
    .Y(_01523_),
    .B1(_05950_));
 sg13g2_o21ai_1 _27935_ (.B1(net9381),
    .Y(_05951_),
    .A1(_13602_),
    .A2(net7366));
 sg13g2_a21oi_1 _27936_ (.A1(net9128),
    .A2(net7369),
    .Y(_01524_),
    .B1(_05951_));
 sg13g2_o21ai_1 _27937_ (.B1(net9392),
    .Y(_05952_),
    .A1(_13653_),
    .A2(net7368));
 sg13g2_a21oi_2 _27938_ (.B1(_05952_),
    .Y(_01525_),
    .A2(net7371),
    .A1(net9160));
 sg13g2_o21ai_1 _27939_ (.B1(net9392),
    .Y(_05953_),
    .A1(net9458),
    .A2(net7356));
 sg13g2_a21oi_1 _27940_ (.A1(_13713_),
    .A2(net7355),
    .Y(_01526_),
    .B1(_05953_));
 sg13g2_o21ai_1 _27941_ (.B1(net9374),
    .Y(_05954_),
    .A1(net9442),
    .A2(net7354));
 sg13g2_a21oi_2 _27942_ (.B1(_05954_),
    .Y(_01527_),
    .A2(net7354),
    .A1(_13777_));
 sg13g2_o21ai_1 _27943_ (.B1(net9392),
    .Y(_05955_),
    .A1(net9434),
    .A2(net7355));
 sg13g2_a21oi_1 _27944_ (.A1(_13330_),
    .A2(net7355),
    .Y(_01528_),
    .B1(_05955_));
 sg13g2_o21ai_1 _27945_ (.B1(net9398),
    .Y(_05956_),
    .A1(net5551),
    .A2(net7358));
 sg13g2_a21oi_1 _27946_ (.A1(_13387_),
    .A2(net7358),
    .Y(_01529_),
    .B1(_05956_));
 sg13g2_o21ai_1 _27947_ (.B1(net9396),
    .Y(_05957_),
    .A1(net5492),
    .A2(net7358));
 sg13g2_a21oi_1 _27948_ (.A1(_13451_),
    .A2(net7358),
    .Y(_01530_),
    .B1(_05957_));
 sg13g2_o21ai_1 _27949_ (.B1(net9393),
    .Y(_05958_),
    .A1(net5237),
    .A2(net7356));
 sg13g2_a21oi_1 _27950_ (.A1(_13516_),
    .A2(net7356),
    .Y(_01531_),
    .B1(_05958_));
 sg13g2_o21ai_1 _27951_ (.B1(net9406),
    .Y(_05959_),
    .A1(net9430),
    .A2(net7359));
 sg13g2_a21oi_1 _27952_ (.A1(_13580_),
    .A2(net7359),
    .Y(_01532_),
    .B1(_05959_));
 sg13g2_o21ai_1 _27953_ (.B1(net9406),
    .Y(_05960_),
    .A1(net9428),
    .A2(net7358));
 sg13g2_a21oi_1 _27954_ (.A1(_13643_),
    .A2(net7358),
    .Y(_01533_),
    .B1(_05960_));
 sg13g2_o21ai_1 _27955_ (.B1(net9403),
    .Y(_05961_),
    .A1(net9426),
    .A2(net7356));
 sg13g2_a21oi_1 _27956_ (.A1(_13734_),
    .A2(net7355),
    .Y(_01534_),
    .B1(_05961_));
 sg13g2_o21ai_1 _27957_ (.B1(net9397),
    .Y(_05962_),
    .A1(net9424),
    .A2(net7357));
 sg13g2_a21oi_1 _27958_ (.A1(_13803_),
    .A2(net7355),
    .Y(_01535_),
    .B1(_05962_));
 sg13g2_and2_1 _27959_ (.A(_10876_),
    .B(_12462_),
    .X(_05963_));
 sg13g2_o21ai_1 _27960_ (.B1(_04656_),
    .Y(_05964_),
    .A1(_10834_),
    .A2(_03811_));
 sg13g2_or4_2 _27961_ (.A(_11017_),
    .B(net7360),
    .C(_05963_),
    .D(_05964_),
    .X(_05965_));
 sg13g2_nor2_1 _27962_ (.A(net9776),
    .B(net7490),
    .Y(_05966_));
 sg13g2_a21oi_2 _27963_ (.B1(_05966_),
    .Y(_05967_),
    .A2(net9776),
    .A1(net3037));
 sg13g2_o21ai_1 _27964_ (.B1(net9397),
    .Y(_05968_),
    .A1(net4800),
    .A2(net7344));
 sg13g2_a21oi_1 _27965_ (.A1(net7344),
    .A2(_05967_),
    .Y(_01536_),
    .B1(_05968_));
 sg13g2_nor2_1 _27966_ (.A(net9776),
    .B(net7668),
    .Y(_05969_));
 sg13g2_a21oi_1 _27967_ (.A1(net2807),
    .A2(net9776),
    .Y(_05970_),
    .B1(_05969_));
 sg13g2_o21ai_1 _27968_ (.B1(net9377),
    .Y(_05971_),
    .A1(net4566),
    .A2(net7342));
 sg13g2_a21oi_1 _27969_ (.A1(net7342),
    .A2(_05970_),
    .Y(_01537_),
    .B1(_05971_));
 sg13g2_nor2_1 _27970_ (.A(net9775),
    .B(net7618),
    .Y(_05972_));
 sg13g2_a21oi_1 _27971_ (.A1(net4321),
    .A2(net9775),
    .Y(_05973_),
    .B1(_05972_));
 sg13g2_o21ai_1 _27972_ (.B1(net9392),
    .Y(_05974_),
    .A1(net4980),
    .A2(net7346));
 sg13g2_a21oi_1 _27973_ (.A1(net7346),
    .A2(_05973_),
    .Y(_01538_),
    .B1(_05974_));
 sg13g2_nor2_1 _27974_ (.A(net9771),
    .B(_12905_),
    .Y(_05975_));
 sg13g2_a21oi_1 _27975_ (.A1(net4144),
    .A2(net9771),
    .Y(_05976_),
    .B1(_05975_));
 sg13g2_o21ai_1 _27976_ (.B1(net9373),
    .Y(_05977_),
    .A1(net4241),
    .A2(net7341));
 sg13g2_a21oi_1 _27977_ (.A1(net7341),
    .A2(_05976_),
    .Y(_01539_),
    .B1(_05977_));
 sg13g2_nand2_1 _27978_ (.Y(_05978_),
    .A(net4847),
    .B(net9775));
 sg13g2_o21ai_1 _27979_ (.B1(_05978_),
    .Y(_05979_),
    .A1(net9775),
    .A2(net7591));
 sg13g2_nor2b_1 _27980_ (.A(_05979_),
    .B_N(net7346),
    .Y(_05980_));
 sg13g2_o21ai_1 _27981_ (.B1(net9394),
    .Y(_05981_),
    .A1(net5426),
    .A2(net7346));
 sg13g2_nor2_1 _27982_ (.A(_05980_),
    .B(_05981_),
    .Y(_01540_));
 sg13g2_nand2_1 _27983_ (.Y(_05982_),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[5] ),
    .B(net9775));
 sg13g2_o21ai_1 _27984_ (.B1(_05982_),
    .Y(_05983_),
    .A1(net9775),
    .A2(_12928_));
 sg13g2_nor2b_1 _27985_ (.A(_05983_),
    .B_N(net7346),
    .Y(_05984_));
 sg13g2_o21ai_1 _27986_ (.B1(net9394),
    .Y(_05985_),
    .A1(net5323),
    .A2(net7346));
 sg13g2_nor2_1 _27987_ (.A(_05984_),
    .B(_05985_),
    .Y(_01541_));
 sg13g2_nand2_1 _27988_ (.Y(_05986_),
    .A(net3923),
    .B(net9775));
 sg13g2_o21ai_1 _27989_ (.B1(_05986_),
    .Y(_05987_),
    .A1(net9775),
    .A2(net7596));
 sg13g2_nor2b_1 _27990_ (.A(_05987_),
    .B_N(net7346),
    .Y(_05988_));
 sg13g2_o21ai_1 _27991_ (.B1(net9394),
    .Y(_05989_),
    .A1(net5272),
    .A2(net7346));
 sg13g2_nor2_1 _27992_ (.A(_05988_),
    .B(_05989_),
    .Y(_01542_));
 sg13g2_nand2_1 _27993_ (.Y(_05990_),
    .A(net4228),
    .B(net9770));
 sg13g2_o21ai_1 _27994_ (.B1(_05990_),
    .Y(_05991_),
    .A1(net9770),
    .A2(net7605));
 sg13g2_nor2b_1 _27995_ (.A(_05991_),
    .B_N(net7337),
    .Y(_05992_));
 sg13g2_o21ai_1 _27996_ (.B1(net9348),
    .Y(_05993_),
    .A1(net5389),
    .A2(net7337));
 sg13g2_nor2_1 _27997_ (.A(_05992_),
    .B(_05993_),
    .Y(_01543_));
 sg13g2_nand2_1 _27998_ (.Y(_05994_),
    .A(net5233),
    .B(net9770));
 sg13g2_o21ai_1 _27999_ (.B1(_05994_),
    .Y(_05995_),
    .A1(net9770),
    .A2(_13007_));
 sg13g2_nor2b_1 _28000_ (.A(_05995_),
    .B_N(net7337),
    .Y(_05996_));
 sg13g2_o21ai_1 _28001_ (.B1(net9348),
    .Y(_05997_),
    .A1(net5501),
    .A2(net7337));
 sg13g2_nor2_1 _28002_ (.A(_05996_),
    .B(_05997_),
    .Y(_01544_));
 sg13g2_nand2_1 _28003_ (.Y(_05998_),
    .A(net5330),
    .B(net9776));
 sg13g2_o21ai_1 _28004_ (.B1(_05998_),
    .Y(_05999_),
    .A1(net9776),
    .A2(net7579));
 sg13g2_nor2b_1 _28005_ (.A(_05999_),
    .B_N(net7342),
    .Y(_06000_));
 sg13g2_o21ai_1 _28006_ (.B1(net9378),
    .Y(_06001_),
    .A1(\soc_I.PC[9] ),
    .A2(net7342));
 sg13g2_nor2_1 _28007_ (.A(_06000_),
    .B(_06001_),
    .Y(_01545_));
 sg13g2_nand2_1 _28008_ (.Y(_06002_),
    .A(net5465),
    .B(net9770));
 sg13g2_o21ai_1 _28009_ (.B1(_06002_),
    .Y(_06003_),
    .A1(net9770),
    .A2(_13029_));
 sg13g2_nor2b_1 _28010_ (.A(_06003_),
    .B_N(net7337),
    .Y(_06004_));
 sg13g2_o21ai_1 _28011_ (.B1(net9346),
    .Y(_06005_),
    .A1(net5441),
    .A2(net7337));
 sg13g2_nor2_1 _28012_ (.A(_06004_),
    .B(_06005_),
    .Y(_01546_));
 sg13g2_nand2_1 _28013_ (.Y(_06006_),
    .A(net4177),
    .B(net9770));
 sg13g2_o21ai_1 _28014_ (.B1(_06006_),
    .Y(_06007_),
    .A1(net9770),
    .A2(net7573));
 sg13g2_nor2b_1 _28015_ (.A(_06007_),
    .B_N(net7337),
    .Y(_06008_));
 sg13g2_o21ai_1 _28016_ (.B1(net9351),
    .Y(_06009_),
    .A1(net5279),
    .A2(net7337));
 sg13g2_nor2_1 _28017_ (.A(_06008_),
    .B(_06009_),
    .Y(_01547_));
 sg13g2_nand2_1 _28018_ (.Y(_06010_),
    .A(net4133),
    .B(net9771));
 sg13g2_o21ai_1 _28019_ (.B1(_06010_),
    .Y(_06011_),
    .A1(net9771),
    .A2(net7545));
 sg13g2_nor2b_1 _28020_ (.A(_06011_),
    .B_N(net7338),
    .Y(_06012_));
 sg13g2_o21ai_1 _28021_ (.B1(net9349),
    .Y(_06013_),
    .A1(net5456),
    .A2(net7338));
 sg13g2_nor2_1 _28022_ (.A(_06012_),
    .B(_06013_),
    .Y(_01548_));
 sg13g2_nand2_1 _28023_ (.Y(_06014_),
    .A(net4123),
    .B(net9772));
 sg13g2_o21ai_1 _28024_ (.B1(_06014_),
    .Y(_06015_),
    .A1(net9771),
    .A2(net7556));
 sg13g2_nor2b_1 _28025_ (.A(_06015_),
    .B_N(net7338),
    .Y(_06016_));
 sg13g2_o21ai_1 _28026_ (.B1(net9362),
    .Y(_06017_),
    .A1(\soc_I.PC[13] ),
    .A2(net7338));
 sg13g2_nor2_1 _28027_ (.A(_06016_),
    .B(net5386),
    .Y(_01549_));
 sg13g2_nor2_1 _28028_ (.A(net9772),
    .B(net7582),
    .Y(_06018_));
 sg13g2_a21oi_1 _28029_ (.A1(net4338),
    .A2(net9772),
    .Y(_06019_),
    .B1(_06018_));
 sg13g2_o21ai_1 _28030_ (.B1(net9363),
    .Y(_06020_),
    .A1(net4664),
    .A2(net7339));
 sg13g2_a21oi_1 _28031_ (.A1(net7339),
    .A2(_06019_),
    .Y(_01550_),
    .B1(_06020_));
 sg13g2_nand2_1 _28032_ (.Y(_06021_),
    .A(net4139),
    .B(net9772));
 sg13g2_o21ai_1 _28033_ (.B1(_06021_),
    .Y(_06022_),
    .A1(net9772),
    .A2(net7566));
 sg13g2_nor2b_1 _28034_ (.A(_06022_),
    .B_N(net7340),
    .Y(_06023_));
 sg13g2_o21ai_1 _28035_ (.B1(net9362),
    .Y(_06024_),
    .A1(net5399),
    .A2(net7340));
 sg13g2_nor2_1 _28036_ (.A(_06023_),
    .B(_06024_),
    .Y(_01551_));
 sg13g2_nand2_1 _28037_ (.Y(_06025_),
    .A(net4203),
    .B(net9773));
 sg13g2_o21ai_1 _28038_ (.B1(_06025_),
    .Y(_06026_),
    .A1(net9773),
    .A2(net7527));
 sg13g2_nor2b_1 _28039_ (.A(_06026_),
    .B_N(net7339),
    .Y(_06027_));
 sg13g2_o21ai_1 _28040_ (.B1(net9366),
    .Y(_06028_),
    .A1(net5226),
    .A2(net7339));
 sg13g2_nor2_1 _28041_ (.A(_06027_),
    .B(_06028_),
    .Y(_01552_));
 sg13g2_nand2_1 _28042_ (.Y(_06029_),
    .A(net4246),
    .B(net9773));
 sg13g2_o21ai_1 _28043_ (.B1(_06029_),
    .Y(_06030_),
    .A1(net9773),
    .A2(net7539));
 sg13g2_nor2b_1 _28044_ (.A(_06030_),
    .B_N(net7340),
    .Y(_06031_));
 sg13g2_o21ai_1 _28045_ (.B1(net9364),
    .Y(_06032_),
    .A1(net5211),
    .A2(net7339));
 sg13g2_nor2_1 _28046_ (.A(_06031_),
    .B(_06032_),
    .Y(_01553_));
 sg13g2_nand2_1 _28047_ (.Y(_06033_),
    .A(net4415),
    .B(net9773));
 sg13g2_o21ai_1 _28048_ (.B1(_06033_),
    .Y(_06034_),
    .A1(net9772),
    .A2(net7533));
 sg13g2_nor2b_1 _28049_ (.A(_06034_),
    .B_N(net7339),
    .Y(_06035_));
 sg13g2_o21ai_1 _28050_ (.B1(net9366),
    .Y(_06036_),
    .A1(net5370),
    .A2(net7339));
 sg13g2_nor2_1 _28051_ (.A(_06035_),
    .B(_06036_),
    .Y(_01554_));
 sg13g2_nand2_1 _28052_ (.Y(_06037_),
    .A(net4550),
    .B(net9773));
 sg13g2_o21ai_1 _28053_ (.B1(_06037_),
    .Y(_06038_),
    .A1(net9773),
    .A2(_13095_));
 sg13g2_nor2b_1 _28054_ (.A(_06038_),
    .B_N(net7340),
    .Y(_06039_));
 sg13g2_o21ai_1 _28055_ (.B1(net9366),
    .Y(_06040_),
    .A1(net5308),
    .A2(net7339));
 sg13g2_nor2_1 _28056_ (.A(_06039_),
    .B(_06040_),
    .Y(_01555_));
 sg13g2_nand2_1 _28057_ (.Y(_06041_),
    .A(net4232),
    .B(net9777));
 sg13g2_o21ai_1 _28058_ (.B1(_06041_),
    .Y(_06042_),
    .A1(net9777),
    .A2(net7510));
 sg13g2_a21oi_1 _28059_ (.A1(net7342),
    .A2(_06042_),
    .Y(_06043_),
    .B1(net9051));
 sg13g2_o21ai_1 _28060_ (.B1(_06043_),
    .Y(_01556_),
    .A1(_10453_),
    .A2(net7342));
 sg13g2_nand2_1 _28061_ (.Y(_06044_),
    .A(net3968),
    .B(net9778));
 sg13g2_o21ai_1 _28062_ (.B1(_06044_),
    .Y(_06045_),
    .A1(net9778),
    .A2(net7515));
 sg13g2_nor2b_1 _28063_ (.A(_06045_),
    .B_N(net7344),
    .Y(_06046_));
 sg13g2_o21ai_1 _28064_ (.B1(net9404),
    .Y(_06047_),
    .A1(net5255),
    .A2(net7344));
 sg13g2_nor2_1 _28065_ (.A(_06046_),
    .B(_06047_),
    .Y(_01557_));
 sg13g2_nand2_1 _28066_ (.Y(_06048_),
    .A(net4403),
    .B(net9778));
 sg13g2_o21ai_1 _28067_ (.B1(_06048_),
    .Y(_06049_),
    .A1(net9778),
    .A2(_13145_));
 sg13g2_nor2b_1 _28068_ (.A(_06049_),
    .B_N(net7345),
    .Y(_06050_));
 sg13g2_o21ai_1 _28069_ (.B1(net9401),
    .Y(_06051_),
    .A1(net5296),
    .A2(net7345));
 sg13g2_nor2_1 _28070_ (.A(_06050_),
    .B(_06051_),
    .Y(_01558_));
 sg13g2_nand2_1 _28071_ (.Y(_06052_),
    .A(net4422),
    .B(net9779));
 sg13g2_o21ai_1 _28072_ (.B1(_06052_),
    .Y(_06053_),
    .A1(net9779),
    .A2(_13132_));
 sg13g2_nor2b_1 _28073_ (.A(_06053_),
    .B_N(net7343),
    .Y(_06054_));
 sg13g2_o21ai_1 _28074_ (.B1(net9387),
    .Y(_06055_),
    .A1(net5258),
    .A2(net7343));
 sg13g2_nor2_1 _28075_ (.A(_06054_),
    .B(_06055_),
    .Y(_01559_));
 sg13g2_nand2_1 _28076_ (.Y(_06056_),
    .A(net4119),
    .B(net9777));
 sg13g2_o21ai_1 _28077_ (.B1(_06056_),
    .Y(_06057_),
    .A1(net9777),
    .A2(net7647));
 sg13g2_nor2b_1 _28078_ (.A(_06057_),
    .B_N(net7344),
    .Y(_06058_));
 sg13g2_o21ai_1 _28079_ (.B1(net9399),
    .Y(_06059_),
    .A1(\soc_I.PC[24] ),
    .A2(net7344));
 sg13g2_nor2_1 _28080_ (.A(_06058_),
    .B(_06059_),
    .Y(_01560_));
 sg13g2_nand2_1 _28081_ (.Y(_06060_),
    .A(net4086),
    .B(net9777));
 sg13g2_o21ai_1 _28082_ (.B1(_06060_),
    .Y(_06061_),
    .A1(net9777),
    .A2(_12497_));
 sg13g2_nor2b_1 _28083_ (.A(_06061_),
    .B_N(net7345),
    .Y(_06062_));
 sg13g2_o21ai_1 _28084_ (.B1(net9404),
    .Y(_06063_),
    .A1(net5383),
    .A2(net7345));
 sg13g2_nor2_1 _28085_ (.A(_06062_),
    .B(_06063_),
    .Y(_01561_));
 sg13g2_nand2_1 _28086_ (.Y(_06064_),
    .A(net4263),
    .B(net9777));
 sg13g2_o21ai_1 _28087_ (.B1(_06064_),
    .Y(_06065_),
    .A1(net9777),
    .A2(_12486_));
 sg13g2_nor2b_1 _28088_ (.A(_06065_),
    .B_N(net7344),
    .Y(_06066_));
 sg13g2_o21ai_1 _28089_ (.B1(net9401),
    .Y(_06067_),
    .A1(net5263),
    .A2(net7344));
 sg13g2_nor2_1 _28090_ (.A(_06066_),
    .B(_06067_),
    .Y(_01562_));
 sg13g2_nor2_1 _28091_ (.A(net9779),
    .B(net7662),
    .Y(_06068_));
 sg13g2_a21oi_1 _28092_ (.A1(net4963),
    .A2(net9779),
    .Y(_06069_),
    .B1(_06068_));
 sg13g2_o21ai_1 _28093_ (.B1(net9389),
    .Y(_06070_),
    .A1(net5097),
    .A2(net7343));
 sg13g2_a21oi_1 _28094_ (.A1(net7343),
    .A2(_06069_),
    .Y(_01563_),
    .B1(_06070_));
 sg13g2_nand2_1 _28095_ (.Y(_06071_),
    .A(net4690),
    .B(net9779));
 sg13g2_o21ai_1 _28096_ (.B1(_06071_),
    .Y(_06072_),
    .A1(net9779),
    .A2(net7641));
 sg13g2_nor2b_1 _28097_ (.A(_06072_),
    .B_N(net7342),
    .Y(_06073_));
 sg13g2_o21ai_1 _28098_ (.B1(net9387),
    .Y(_06074_),
    .A1(net5458),
    .A2(net7342));
 sg13g2_nor2_1 _28099_ (.A(_06073_),
    .B(_06074_),
    .Y(_01564_));
 sg13g2_nand2_1 _28100_ (.Y(_06075_),
    .A(net4672),
    .B(net9774));
 sg13g2_o21ai_1 _28101_ (.B1(_06075_),
    .Y(_06076_),
    .A1(net9774),
    .A2(_12539_));
 sg13g2_a21oi_1 _28102_ (.A1(net7341),
    .A2(_06076_),
    .Y(_06077_),
    .B1(net9040));
 sg13g2_o21ai_1 _28103_ (.B1(_06077_),
    .Y(_01565_),
    .A1(_10452_),
    .A2(net7341));
 sg13g2_nand2_1 _28104_ (.Y(_06078_),
    .A(net3885),
    .B(net9774));
 sg13g2_o21ai_1 _28105_ (.B1(_06078_),
    .Y(_06079_),
    .A1(net9774),
    .A2(net7624));
 sg13g2_nor2b_1 _28106_ (.A(_06079_),
    .B_N(net7341),
    .Y(_06080_));
 sg13g2_o21ai_1 _28107_ (.B1(net9381),
    .Y(_06081_),
    .A1(net4242),
    .A2(net7341));
 sg13g2_nor2_1 _28108_ (.A(_06080_),
    .B(_06081_),
    .Y(_01566_));
 sg13g2_nand2_1 _28109_ (.Y(_06082_),
    .A(net4790),
    .B(net9772));
 sg13g2_o21ai_1 _28110_ (.B1(_06082_),
    .Y(_06083_),
    .A1(net9772),
    .A2(_12530_));
 sg13g2_nor2b_1 _28111_ (.A(_06083_),
    .B_N(net7340),
    .Y(_06084_));
 sg13g2_o21ai_1 _28112_ (.B1(net9354),
    .Y(_06085_),
    .A1(net4981),
    .A2(net7340));
 sg13g2_nor2_1 _28113_ (.A(_06084_),
    .B(_06085_),
    .Y(_01567_));
 sg13g2_nand2_2 _28114_ (.Y(_06086_),
    .A(_14126_),
    .B(_03742_));
 sg13g2_nand2_1 _28115_ (.Y(_06087_),
    .A(net3181),
    .B(net7876));
 sg13g2_o21ai_1 _28116_ (.B1(_06087_),
    .Y(_01568_),
    .A1(net7486),
    .A2(net7876));
 sg13g2_nand2_1 _28117_ (.Y(_06088_),
    .A(net2872),
    .B(net7875));
 sg13g2_o21ai_1 _28118_ (.B1(_06088_),
    .Y(_01569_),
    .A1(net7665),
    .A2(net7875));
 sg13g2_nand2_1 _28119_ (.Y(_06089_),
    .A(net2868),
    .B(net7876));
 sg13g2_o21ai_1 _28120_ (.B1(_06089_),
    .Y(_01570_),
    .A1(net7615),
    .A2(net7876));
 sg13g2_nand2_1 _28121_ (.Y(_06090_),
    .A(net3550),
    .B(net7876));
 sg13g2_o21ai_1 _28122_ (.B1(_06090_),
    .Y(_01571_),
    .A1(net7609),
    .A2(net7877));
 sg13g2_nand2_1 _28123_ (.Y(_06091_),
    .A(net2747),
    .B(net7873));
 sg13g2_o21ai_1 _28124_ (.B1(_06091_),
    .Y(_01572_),
    .A1(net7587),
    .A2(net7873));
 sg13g2_nand2_1 _28125_ (.Y(_06092_),
    .A(net2881),
    .B(net7872));
 sg13g2_o21ai_1 _28126_ (.B1(_06092_),
    .Y(_01573_),
    .A1(net7597),
    .A2(net7872));
 sg13g2_nand2_1 _28127_ (.Y(_06093_),
    .A(net3358),
    .B(net7875));
 sg13g2_o21ai_1 _28128_ (.B1(_06093_),
    .Y(_01574_),
    .A1(net7593),
    .A2(net7875));
 sg13g2_nand2_1 _28129_ (.Y(_06094_),
    .A(net3352),
    .B(net7869));
 sg13g2_o21ai_1 _28130_ (.B1(_06094_),
    .Y(_01575_),
    .A1(net7606),
    .A2(net7868));
 sg13g2_nand2_1 _28131_ (.Y(_06095_),
    .A(net2867),
    .B(net7872));
 sg13g2_o21ai_1 _28132_ (.B1(_06095_),
    .Y(_01576_),
    .A1(net7558),
    .A2(net7872));
 sg13g2_nand2_1 _28133_ (.Y(_06096_),
    .A(net2995),
    .B(net7874));
 sg13g2_o21ai_1 _28134_ (.B1(_06096_),
    .Y(_01577_),
    .A1(net7574),
    .A2(net7874));
 sg13g2_nand2_1 _28135_ (.Y(_06097_),
    .A(net2973),
    .B(net7874));
 sg13g2_o21ai_1 _28136_ (.B1(_06097_),
    .Y(_01578_),
    .A1(net7546),
    .A2(net7874));
 sg13g2_nand2_1 _28137_ (.Y(_06098_),
    .A(net2825),
    .B(net7868));
 sg13g2_o21ai_1 _28138_ (.B1(_06098_),
    .Y(_01579_),
    .A1(net7571),
    .A2(net7868));
 sg13g2_nand2_1 _28139_ (.Y(_06099_),
    .A(net2754),
    .B(net7874));
 sg13g2_o21ai_1 _28140_ (.B1(_06099_),
    .Y(_01580_),
    .A1(net7541),
    .A2(net7874));
 sg13g2_nand2_1 _28141_ (.Y(_06100_),
    .A(net2733),
    .B(net7874));
 sg13g2_o21ai_1 _28142_ (.B1(_06100_),
    .Y(_01581_),
    .A1(net7551),
    .A2(net7874));
 sg13g2_nand2_1 _28143_ (.Y(_06101_),
    .A(net2853),
    .B(net7870));
 sg13g2_o21ai_1 _28144_ (.B1(_06101_),
    .Y(_01582_),
    .A1(net7580),
    .A2(net7870));
 sg13g2_nand2_1 _28145_ (.Y(_06102_),
    .A(net3258),
    .B(net7869));
 sg13g2_o21ai_1 _28146_ (.B1(_06102_),
    .Y(_01583_),
    .A1(net7566),
    .A2(net7869));
 sg13g2_nand2_1 _28147_ (.Y(_06103_),
    .A(net3440),
    .B(net7868));
 sg13g2_o21ai_1 _28148_ (.B1(_06103_),
    .Y(_01584_),
    .A1(net7526),
    .A2(net7868));
 sg13g2_nand2_1 _28149_ (.Y(_06104_),
    .A(net2775),
    .B(net7868));
 sg13g2_o21ai_1 _28150_ (.B1(_06104_),
    .Y(_01585_),
    .A1(net7537),
    .A2(net7868));
 sg13g2_nand2_1 _28151_ (.Y(_06105_),
    .A(net2922),
    .B(net7870));
 sg13g2_o21ai_1 _28152_ (.B1(_06105_),
    .Y(_01586_),
    .A1(net7532),
    .A2(net7870));
 sg13g2_nand2_1 _28153_ (.Y(_06106_),
    .A(net2929),
    .B(net7870));
 sg13g2_o21ai_1 _28154_ (.B1(_06106_),
    .Y(_01587_),
    .A1(net7519),
    .A2(net7870));
 sg13g2_nand2_1 _28155_ (.Y(_06107_),
    .A(net2721),
    .B(net7873));
 sg13g2_o21ai_1 _28156_ (.B1(_06107_),
    .Y(_01588_),
    .A1(net7504),
    .A2(net7873));
 sg13g2_nand2_1 _28157_ (.Y(_06108_),
    .A(net2742),
    .B(_06086_));
 sg13g2_o21ai_1 _28158_ (.B1(_06108_),
    .Y(_01589_),
    .A1(net7512),
    .A2(net7871));
 sg13g2_nand2_1 _28159_ (.Y(_06109_),
    .A(net3014),
    .B(net7877));
 sg13g2_o21ai_1 _28160_ (.B1(_06109_),
    .Y(_01590_),
    .A1(net7494),
    .A2(net7875));
 sg13g2_nand2_1 _28161_ (.Y(_06110_),
    .A(net3489),
    .B(net7869));
 sg13g2_o21ai_1 _28162_ (.B1(_06110_),
    .Y(_01591_),
    .A1(net7503),
    .A2(net7869));
 sg13g2_nand2_1 _28163_ (.Y(_06111_),
    .A(net2912),
    .B(net7872));
 sg13g2_o21ai_1 _28164_ (.B1(_06111_),
    .Y(_01592_),
    .A1(net7646),
    .A2(net7872));
 sg13g2_nand2_1 _28165_ (.Y(_06112_),
    .A(net3713),
    .B(net7876));
 sg13g2_o21ai_1 _28166_ (.B1(_06112_),
    .Y(_01593_),
    .A1(net7651),
    .A2(net7876));
 sg13g2_nand2_1 _28167_ (.Y(_06113_),
    .A(net3747),
    .B(net7875));
 sg13g2_o21ai_1 _28168_ (.B1(_06113_),
    .Y(_01594_),
    .A1(net7653),
    .A2(net7875));
 sg13g2_nand2_1 _28169_ (.Y(_06114_),
    .A(net3450),
    .B(net7871));
 sg13g2_o21ai_1 _28170_ (.B1(_06114_),
    .Y(_01595_),
    .A1(net7661),
    .A2(net7871));
 sg13g2_nand2_1 _28171_ (.Y(_06115_),
    .A(net2752),
    .B(net7871));
 sg13g2_o21ai_1 _28172_ (.B1(_06115_),
    .Y(_01596_),
    .A1(net7640),
    .A2(net7871));
 sg13g2_nand2_1 _28173_ (.Y(_06116_),
    .A(net3137),
    .B(net7872));
 sg13g2_o21ai_1 _28174_ (.B1(_06116_),
    .Y(_01597_),
    .A1(net7625),
    .A2(net7872));
 sg13g2_nand2_1 _28175_ (.Y(_06117_),
    .A(net2924),
    .B(net7871));
 sg13g2_o21ai_1 _28176_ (.B1(_06117_),
    .Y(_01598_),
    .A1(net7619),
    .A2(net7871));
 sg13g2_nand2_1 _28177_ (.Y(_06118_),
    .A(net3337),
    .B(net7868));
 sg13g2_o21ai_1 _28178_ (.B1(_06118_),
    .Y(_01599_),
    .A1(net7633),
    .A2(net7869));
 sg13g2_nor2_1 _28179_ (.A(net4970),
    .B(net9340),
    .Y(_06119_));
 sg13g2_a21oi_1 _28180_ (.A1(net9340),
    .A2(_13182_),
    .Y(_01600_),
    .B1(_06119_));
 sg13g2_nor3_2 _28181_ (.A(\soc_I.clint_I.div[2] ),
    .B(\soc_I.clint_I.div[1] ),
    .C(\soc_I.clint_I.div[0] ),
    .Y(_06120_));
 sg13g2_nor2b_2 _28182_ (.A(\soc_I.clint_I.div[3] ),
    .B_N(_06120_),
    .Y(_06121_));
 sg13g2_nor2_1 _28183_ (.A(\soc_I.clint_I.div[5] ),
    .B(\soc_I.clint_I.div[4] ),
    .Y(_06122_));
 sg13g2_and2_1 _28184_ (.A(_06121_),
    .B(_06122_),
    .X(_06123_));
 sg13g2_nor2b_1 _28185_ (.A(\soc_I.clint_I.div[6] ),
    .B_N(_06123_),
    .Y(_06124_));
 sg13g2_nand2b_1 _28186_ (.Y(_06125_),
    .B(_06124_),
    .A_N(\soc_I.clint_I.div[7] ));
 sg13g2_nor3_1 _28187_ (.A(\soc_I.clint_I.div[9] ),
    .B(\soc_I.clint_I.div[8] ),
    .C(_06125_),
    .Y(_06126_));
 sg13g2_nor2b_1 _28188_ (.A(\soc_I.clint_I.div[10] ),
    .B_N(_06126_),
    .Y(_06127_));
 sg13g2_nor2b_1 _28189_ (.A(\soc_I.clint_I.div[11] ),
    .B_N(_06127_),
    .Y(_06128_));
 sg13g2_nor2_1 _28190_ (.A(\soc_I.clint_I.div[13] ),
    .B(\soc_I.clint_I.div[12] ),
    .Y(_06129_));
 sg13g2_and2_1 _28191_ (.A(_06128_),
    .B(_06129_),
    .X(_06130_));
 sg13g2_nand2b_1 _28192_ (.Y(_06131_),
    .B(_06130_),
    .A_N(\soc_I.clint_I.div[14] ));
 sg13g2_a21oi_2 _28193_ (.B1(_10601_),
    .Y(_06132_),
    .A2(_06131_),
    .A1(\soc_I.clint_I.div[15] ));
 sg13g2_and3_1 _28194_ (.X(_06133_),
    .A(\soc_I.clint_I.div[15] ),
    .B(_10601_),
    .C(_06131_));
 sg13g2_xnor2_1 _28195_ (.Y(_06134_),
    .A(\soc_I.clint_I.div[14] ),
    .B(_06130_));
 sg13g2_nor2_1 _28196_ (.A(\soc_I.clint_I.tick_cnt[14] ),
    .B(_06134_),
    .Y(_06135_));
 sg13g2_nand2_1 _28197_ (.Y(_06136_),
    .A(\soc_I.clint_I.tick_cnt[14] ),
    .B(_06134_));
 sg13g2_inv_1 _28198_ (.Y(_06137_),
    .A(_06136_));
 sg13g2_nor4_1 _28199_ (.A(_06132_),
    .B(_06133_),
    .C(_06135_),
    .D(_06137_),
    .Y(_06138_));
 sg13g2_nand2_1 _28200_ (.Y(_06139_),
    .A(_00248_),
    .B(_06128_));
 sg13g2_xor2_1 _28201_ (.B(\soc_I.clint_I.tick_cnt[13] ),
    .A(\soc_I.clint_I.div[13] ),
    .X(_06140_));
 sg13g2_xnor2_1 _28202_ (.Y(_06141_),
    .A(_06139_),
    .B(_06140_));
 sg13g2_xnor2_1 _28203_ (.Y(_06142_),
    .A(_00248_),
    .B(_06128_));
 sg13g2_and2_1 _28204_ (.A(_10600_),
    .B(_06142_),
    .X(_06143_));
 sg13g2_nor2_1 _28205_ (.A(_10600_),
    .B(_06142_),
    .Y(_06144_));
 sg13g2_nor3_1 _28206_ (.A(_06141_),
    .B(_06143_),
    .C(_06144_),
    .Y(_06145_));
 sg13g2_xnor2_1 _28207_ (.Y(_06146_),
    .A(\soc_I.clint_I.div[11] ),
    .B(_06127_));
 sg13g2_xnor2_1 _28208_ (.Y(_06147_),
    .A(\soc_I.clint_I.tick_cnt[11] ),
    .B(_06146_));
 sg13g2_xnor2_1 _28209_ (.Y(_06148_),
    .A(\soc_I.clint_I.div[10] ),
    .B(_06126_));
 sg13g2_xnor2_1 _28210_ (.Y(_06149_),
    .A(\soc_I.clint_I.tick_cnt[10] ),
    .B(_06148_));
 sg13g2_nor2_1 _28211_ (.A(_06147_),
    .B(_06149_),
    .Y(_06150_));
 sg13g2_nor2_1 _28212_ (.A(\soc_I.clint_I.div[15] ),
    .B(_06131_),
    .Y(_06151_));
 sg13g2_or2_2 _28213_ (.X(_06152_),
    .B(_06125_),
    .A(_10598_));
 sg13g2_xor2_1 _28214_ (.B(\soc_I.clint_I.tick_cnt[9] ),
    .A(\soc_I.clint_I.div[9] ),
    .X(_06153_));
 sg13g2_xor2_1 _28215_ (.B(\soc_I.clint_I.div[0] ),
    .A(\soc_I.clint_I.div[1] ),
    .X(_06154_));
 sg13g2_or2_1 _28216_ (.X(_06155_),
    .B(_06154_),
    .A(\soc_I.clint_I.tick_cnt[1] ));
 sg13g2_nor2_1 _28217_ (.A(\soc_I.clint_I.div[0] ),
    .B(\soc_I.clint_I.tick_cnt[0] ),
    .Y(_06156_));
 sg13g2_nor3_1 _28218_ (.A(\soc_I.clint_I.tick_cnt[16] ),
    .B(\soc_I.clint_I.tick_cnt[17] ),
    .C(_06156_),
    .Y(_06157_));
 sg13g2_a22oi_1 _28219_ (.Y(_06158_),
    .B1(\soc_I.clint_I.tick_cnt[1] ),
    .B2(_06154_),
    .A2(\soc_I.clint_I.tick_cnt[0] ),
    .A1(\soc_I.clint_I.div[0] ));
 sg13g2_o21ai_1 _28220_ (.B1(\soc_I.clint_I.div[2] ),
    .Y(_06159_),
    .A1(\soc_I.clint_I.div[1] ),
    .A2(\soc_I.clint_I.div[0] ));
 sg13g2_nand2b_1 _28221_ (.Y(_06160_),
    .B(_06159_),
    .A_N(_06120_));
 sg13g2_xnor2_1 _28222_ (.Y(_06161_),
    .A(\soc_I.clint_I.tick_cnt[2] ),
    .B(_06160_));
 sg13g2_nand4_1 _28223_ (.B(_06157_),
    .C(_06158_),
    .A(_06155_),
    .Y(_06162_),
    .D(_06161_));
 sg13g2_xnor2_1 _28224_ (.Y(_06163_),
    .A(\soc_I.clint_I.div[3] ),
    .B(_06120_));
 sg13g2_xnor2_1 _28225_ (.Y(_06164_),
    .A(\soc_I.clint_I.tick_cnt[3] ),
    .B(_06163_));
 sg13g2_nor2_1 _28226_ (.A(_06162_),
    .B(_06164_),
    .Y(_06165_));
 sg13g2_xnor2_1 _28227_ (.Y(_06166_),
    .A(\soc_I.clint_I.div[5] ),
    .B(\soc_I.clint_I.tick_cnt[5] ));
 sg13g2_o21ai_1 _28228_ (.B1(_06166_),
    .Y(_06167_),
    .A1(\soc_I.clint_I.tick_cnt[4] ),
    .A2(_06121_));
 sg13g2_a22oi_1 _28229_ (.Y(_06168_),
    .B1(_06166_),
    .B2(_00246_),
    .A2(_06121_),
    .A1(\soc_I.clint_I.tick_cnt[4] ));
 sg13g2_o21ai_1 _28230_ (.B1(_06165_),
    .Y(_06169_),
    .A1(_06167_),
    .A2(_06168_));
 sg13g2_a21oi_1 _28231_ (.A1(_06152_),
    .A2(_06153_),
    .Y(_06170_),
    .B1(_06169_));
 sg13g2_o21ai_1 _28232_ (.B1(_06170_),
    .Y(_06171_),
    .A1(_06152_),
    .A2(_06153_));
 sg13g2_nand2_1 _28233_ (.Y(_06172_),
    .A(_10598_),
    .B(_06125_));
 sg13g2_nand3_1 _28234_ (.B(_06152_),
    .C(_06172_),
    .A(\soc_I.clint_I.tick_cnt[8] ),
    .Y(_06173_));
 sg13g2_xnor2_1 _28235_ (.Y(_06174_),
    .A(\soc_I.clint_I.div[6] ),
    .B(_06123_));
 sg13g2_nor2_1 _28236_ (.A(\soc_I.clint_I.tick_cnt[6] ),
    .B(_06174_),
    .Y(_06175_));
 sg13g2_nand2_1 _28237_ (.Y(_06176_),
    .A(\soc_I.clint_I.tick_cnt[6] ),
    .B(_06174_));
 sg13g2_nand2b_1 _28238_ (.Y(_06177_),
    .B(_06176_),
    .A_N(_06175_));
 sg13g2_o21ai_1 _28239_ (.B1(_06167_),
    .Y(_06178_),
    .A1(_10597_),
    .A2(_06168_));
 sg13g2_nor2b_1 _28240_ (.A(_06177_),
    .B_N(_06178_),
    .Y(_06179_));
 sg13g2_a21o_1 _28241_ (.A2(_06172_),
    .A1(_06152_),
    .B1(\soc_I.clint_I.tick_cnt[8] ),
    .X(_06180_));
 sg13g2_xnor2_1 _28242_ (.Y(_06181_),
    .A(\soc_I.clint_I.div[7] ),
    .B(_06124_));
 sg13g2_xor2_1 _28243_ (.B(_06181_),
    .A(\soc_I.clint_I.tick_cnt[7] ),
    .X(_06182_));
 sg13g2_nand4_1 _28244_ (.B(_06179_),
    .C(_06180_),
    .A(_06173_),
    .Y(_06183_),
    .D(_06182_));
 sg13g2_nor3_1 _28245_ (.A(_06151_),
    .B(_06171_),
    .C(_06183_),
    .Y(_06184_));
 sg13g2_nand4_1 _28246_ (.B(_06145_),
    .C(_06150_),
    .A(_06138_),
    .Y(_06185_),
    .D(_06184_));
 sg13g2_nand2_1 _28247_ (.Y(_06186_),
    .A(\soc_I.clint_I.tick_cnt[7] ),
    .B(_06181_));
 sg13g2_nor2_1 _28248_ (.A(\soc_I.clint_I.tick_cnt[7] ),
    .B(_06181_),
    .Y(_06187_));
 sg13g2_nor4_1 _28249_ (.A(_06162_),
    .B(_06164_),
    .C(_06175_),
    .D(_06187_),
    .Y(_06188_));
 sg13g2_and2_1 _28250_ (.A(\soc_I.clint_I.tick_cnt[10] ),
    .B(_06148_),
    .X(_06189_));
 sg13g2_xnor2_1 _28251_ (.Y(_06190_),
    .A(_06152_),
    .B(_06153_));
 sg13g2_nor2_1 _28252_ (.A(\soc_I.clint_I.tick_cnt[10] ),
    .B(_06148_),
    .Y(_06191_));
 sg13g2_nand2_1 _28253_ (.Y(_06192_),
    .A(_00246_),
    .B(_06121_));
 sg13g2_xnor2_1 _28254_ (.Y(_06193_),
    .A(_00246_),
    .B(_06121_));
 sg13g2_xnor2_1 _28255_ (.Y(_06194_),
    .A(\soc_I.clint_I.tick_cnt[4] ),
    .B(_06193_));
 sg13g2_xnor2_1 _28256_ (.Y(_06195_),
    .A(_06166_),
    .B(_06192_));
 sg13g2_and2_1 _28257_ (.A(_06194_),
    .B(_06195_),
    .X(_06196_));
 sg13g2_nand4_1 _28258_ (.B(_06176_),
    .C(_06180_),
    .A(_06173_),
    .Y(_06197_),
    .D(_06196_));
 sg13g2_nor4_1 _28259_ (.A(_06189_),
    .B(_06190_),
    .C(_06191_),
    .D(_06197_),
    .Y(_06198_));
 sg13g2_nand3_1 _28260_ (.B(_06188_),
    .C(_06198_),
    .A(_06186_),
    .Y(_06199_));
 sg13g2_nor3_1 _28261_ (.A(_06132_),
    .B(_06135_),
    .C(_06199_),
    .Y(_06200_));
 sg13g2_xor2_1 _28262_ (.B(_06139_),
    .A(\soc_I.clint_I.div[13] ),
    .X(_06201_));
 sg13g2_or2_1 _28263_ (.X(_06202_),
    .B(_06201_),
    .A(\soc_I.clint_I.tick_cnt[13] ));
 sg13g2_nor2b_1 _28264_ (.A(_06133_),
    .B_N(_06202_),
    .Y(_06203_));
 sg13g2_and2_1 _28265_ (.A(\soc_I.clint_I.tick_cnt[13] ),
    .B(_06201_),
    .X(_06204_));
 sg13g2_nor4_1 _28266_ (.A(_06143_),
    .B(_06144_),
    .C(_06147_),
    .D(_06151_),
    .Y(_06205_));
 sg13g2_nor2b_1 _28267_ (.A(_06204_),
    .B_N(_06205_),
    .Y(_06206_));
 sg13g2_nand4_1 _28268_ (.B(_06200_),
    .C(_06203_),
    .A(_06136_),
    .Y(_06207_),
    .D(_06206_));
 sg13g2_xor2_1 _28269_ (.B(_06152_),
    .A(\soc_I.clint_I.div[9] ),
    .X(_06208_));
 sg13g2_nor2_1 _28270_ (.A(\soc_I.clint_I.tick_cnt[9] ),
    .B(_06208_),
    .Y(_06209_));
 sg13g2_xor2_1 _28271_ (.B(_06192_),
    .A(\soc_I.clint_I.div[5] ),
    .X(_06210_));
 sg13g2_o21ai_1 _28272_ (.B1(_06194_),
    .Y(_06211_),
    .A1(\soc_I.clint_I.tick_cnt[5] ),
    .A2(_06210_));
 sg13g2_nor2_1 _28273_ (.A(_06177_),
    .B(_06211_),
    .Y(_06212_));
 sg13g2_nand2_1 _28274_ (.Y(_06213_),
    .A(\soc_I.clint_I.tick_cnt[5] ),
    .B(_06210_));
 sg13g2_nand3_1 _28275_ (.B(_06186_),
    .C(_06213_),
    .A(_06165_),
    .Y(_06214_));
 sg13g2_and2_1 _28276_ (.A(\soc_I.clint_I.tick_cnt[9] ),
    .B(_06208_),
    .X(_06215_));
 sg13g2_nor3_1 _28277_ (.A(_06187_),
    .B(_06214_),
    .C(_06215_),
    .Y(_06216_));
 sg13g2_nand4_1 _28278_ (.B(_06180_),
    .C(_06212_),
    .A(_06173_),
    .Y(_06217_),
    .D(_06216_));
 sg13g2_nor4_1 _28279_ (.A(_06189_),
    .B(_06191_),
    .C(_06209_),
    .D(_06217_),
    .Y(_06218_));
 sg13g2_nor2b_1 _28280_ (.A(_06133_),
    .B_N(_06218_),
    .Y(_06219_));
 sg13g2_nand4_1 _28281_ (.B(_06202_),
    .C(_06205_),
    .A(_06136_),
    .Y(_06220_),
    .D(_06219_));
 sg13g2_nor4_2 _28282_ (.A(_06132_),
    .B(_06135_),
    .C(_06204_),
    .Y(_06221_),
    .D(_06220_));
 sg13g2_nand2_1 _28283_ (.Y(_06222_),
    .A(net9001),
    .B(_06207_));
 sg13g2_and3_1 _28284_ (.X(_01601_),
    .A(net9001),
    .B(net2603),
    .C(_06207_));
 sg13g2_xnor2_1 _28285_ (.Y(_06223_),
    .A(\soc_I.clint_I.tick_cnt[0] ),
    .B(net4885));
 sg13g2_nor2_1 _28286_ (.A(net7684),
    .B(net4886),
    .Y(_01602_));
 sg13g2_and3_1 _28287_ (.X(_06224_),
    .A(\soc_I.clint_I.tick_cnt[0] ),
    .B(\soc_I.clint_I.tick_cnt[1] ),
    .C(net3625));
 sg13g2_a21oi_1 _28288_ (.A1(\soc_I.clint_I.tick_cnt[0] ),
    .A2(\soc_I.clint_I.tick_cnt[1] ),
    .Y(_06225_),
    .B1(net3625));
 sg13g2_nor3_1 _28289_ (.A(net7683),
    .B(_06224_),
    .C(net3626),
    .Y(_01603_));
 sg13g2_and2_1 _28290_ (.A(net4432),
    .B(_06224_),
    .X(_06226_));
 sg13g2_nor2_1 _28291_ (.A(net4432),
    .B(_06224_),
    .Y(_06227_));
 sg13g2_nor3_1 _28292_ (.A(net7683),
    .B(_06226_),
    .C(net4433),
    .Y(_01604_));
 sg13g2_and2_1 _28293_ (.A(net4990),
    .B(_06226_),
    .X(_06228_));
 sg13g2_nor2_1 _28294_ (.A(net4990),
    .B(_06226_),
    .Y(_06229_));
 sg13g2_nor3_1 _28295_ (.A(net7684),
    .B(_06228_),
    .C(_06229_),
    .Y(_01605_));
 sg13g2_and2_1 _28296_ (.A(net5031),
    .B(_06228_),
    .X(_06230_));
 sg13g2_nor2_1 _28297_ (.A(net5031),
    .B(_06228_),
    .Y(_06231_));
 sg13g2_nor3_1 _28298_ (.A(_06222_),
    .B(_06230_),
    .C(_06231_),
    .Y(_01606_));
 sg13g2_and2_1 _28299_ (.A(net4607),
    .B(_06230_),
    .X(_06232_));
 sg13g2_nor2_1 _28300_ (.A(net4607),
    .B(_06230_),
    .Y(_06233_));
 sg13g2_nor3_1 _28301_ (.A(_06222_),
    .B(_06232_),
    .C(net4608),
    .Y(_01607_));
 sg13g2_and2_1 _28302_ (.A(net4954),
    .B(_06232_),
    .X(_06234_));
 sg13g2_nor2_1 _28303_ (.A(net4954),
    .B(_06232_),
    .Y(_06235_));
 sg13g2_nor3_1 _28304_ (.A(net7684),
    .B(_06234_),
    .C(_06235_),
    .Y(_01608_));
 sg13g2_and2_1 _28305_ (.A(net4326),
    .B(_06234_),
    .X(_06236_));
 sg13g2_nor2_1 _28306_ (.A(net4326),
    .B(_06234_),
    .Y(_06237_));
 sg13g2_nor3_1 _28307_ (.A(net7684),
    .B(_06236_),
    .C(net4327),
    .Y(_01609_));
 sg13g2_xnor2_1 _28308_ (.Y(_06238_),
    .A(net5270),
    .B(_06236_));
 sg13g2_nor2_1 _28309_ (.A(net7684),
    .B(_06238_),
    .Y(_01610_));
 sg13g2_and3_1 _28310_ (.X(_06239_),
    .A(net5571),
    .B(net4844),
    .C(_06236_));
 sg13g2_a21oi_1 _28311_ (.A1(\soc_I.clint_I.tick_cnt[9] ),
    .A2(_06236_),
    .Y(_06240_),
    .B1(net4844));
 sg13g2_nor3_1 _28312_ (.A(net7684),
    .B(_06239_),
    .C(net4845),
    .Y(_01611_));
 sg13g2_and2_1 _28313_ (.A(net4685),
    .B(_06239_),
    .X(_06241_));
 sg13g2_nor2_1 _28314_ (.A(net4685),
    .B(_06239_),
    .Y(_06242_));
 sg13g2_nor3_1 _28315_ (.A(net7684),
    .B(_06241_),
    .C(net4686),
    .Y(_01612_));
 sg13g2_and2_1 _28316_ (.A(net4155),
    .B(_06241_),
    .X(_06243_));
 sg13g2_nor2_1 _28317_ (.A(net4155),
    .B(_06241_),
    .Y(_06244_));
 sg13g2_nor3_1 _28318_ (.A(net7683),
    .B(_06243_),
    .C(net4156),
    .Y(_01613_));
 sg13g2_and2_1 _28319_ (.A(net5098),
    .B(_06243_),
    .X(_06245_));
 sg13g2_nor2_1 _28320_ (.A(net5098),
    .B(_06243_),
    .Y(_06246_));
 sg13g2_nor3_1 _28321_ (.A(net7683),
    .B(_06245_),
    .C(_06246_),
    .Y(_01614_));
 sg13g2_and2_1 _28322_ (.A(net4947),
    .B(_06245_),
    .X(_06247_));
 sg13g2_nor2_1 _28323_ (.A(net4947),
    .B(_06245_),
    .Y(_06248_));
 sg13g2_nor3_1 _28324_ (.A(net7683),
    .B(_06247_),
    .C(_06248_),
    .Y(_01615_));
 sg13g2_xnor2_1 _28325_ (.Y(_06249_),
    .A(net4838),
    .B(_06247_));
 sg13g2_nor2_1 _28326_ (.A(net7683),
    .B(net4839),
    .Y(_01616_));
 sg13g2_nand3_1 _28327_ (.B(net5118),
    .C(_06247_),
    .A(net4838),
    .Y(_06250_));
 sg13g2_a21oi_1 _28328_ (.A1(net4838),
    .A2(_06247_),
    .Y(_06251_),
    .B1(net5118));
 sg13g2_nor2_1 _28329_ (.A(net7683),
    .B(_06251_),
    .Y(_06252_));
 sg13g2_and2_1 _28330_ (.A(_06250_),
    .B(_06252_),
    .X(_01617_));
 sg13g2_xor2_1 _28331_ (.B(_06250_),
    .A(net4334),
    .X(_06253_));
 sg13g2_nor2_1 _28332_ (.A(net7683),
    .B(net4335),
    .Y(_01618_));
 sg13g2_a21oi_1 _28333_ (.A1(_13225_),
    .A2(_14437_),
    .Y(_06254_),
    .B1(net5145));
 sg13g2_nor4_1 _28334_ (.A(net7468),
    .B(_13212_),
    .C(_13977_),
    .D(_14438_),
    .Y(_06255_));
 sg13g2_nor3_1 _28335_ (.A(net9013),
    .B(_06254_),
    .C(_06255_),
    .Y(_01619_));
 sg13g2_nor2_2 _28336_ (.A(_13187_),
    .B(_14438_),
    .Y(_06256_));
 sg13g2_nor3_1 _28337_ (.A(net7467),
    .B(net7465),
    .C(_14438_),
    .Y(_06257_));
 sg13g2_o21ai_1 _28338_ (.B1(net9322),
    .Y(_06258_),
    .A1(net4799),
    .A2(net7434));
 sg13g2_a21oi_1 _28339_ (.A1(_13978_),
    .A2(_06256_),
    .Y(_01620_),
    .B1(_06258_));
 sg13g2_o21ai_1 _28340_ (.B1(net9322),
    .Y(_06259_),
    .A1(net4510),
    .A2(net7434));
 sg13g2_a21oi_1 _28341_ (.A1(net8612),
    .A2(_06256_),
    .Y(_01621_),
    .B1(_06259_));
 sg13g2_o21ai_1 _28342_ (.B1(net9320),
    .Y(_06260_),
    .A1(net4899),
    .A2(_06257_));
 sg13g2_a21oi_1 _28343_ (.A1(net8610),
    .A2(_06256_),
    .Y(_01622_),
    .B1(_06260_));
 sg13g2_o21ai_1 _28344_ (.B1(net9320),
    .Y(_06261_),
    .A1(net5040),
    .A2(net7434));
 sg13g2_a21oi_1 _28345_ (.A1(net8549),
    .A2(_06257_),
    .Y(_01623_),
    .B1(_06261_));
 sg13g2_o21ai_1 _28346_ (.B1(net9320),
    .Y(_06262_),
    .A1(net4816),
    .A2(net7434));
 sg13g2_a21oi_1 _28347_ (.A1(net8608),
    .A2(_06256_),
    .Y(_01624_),
    .B1(_06262_));
 sg13g2_o21ai_1 _28348_ (.B1(net9320),
    .Y(_06263_),
    .A1(net4708),
    .A2(net7434));
 sg13g2_a21oi_1 _28349_ (.A1(net8606),
    .A2(_06256_),
    .Y(_01625_),
    .B1(_06263_));
 sg13g2_o21ai_1 _28350_ (.B1(net9320),
    .Y(_06264_),
    .A1(net5038),
    .A2(net7434));
 sg13g2_a21oi_1 _28351_ (.A1(net8604),
    .A2(_06256_),
    .Y(_01626_),
    .B1(_06264_));
 sg13g2_o21ai_1 _28352_ (.B1(net9311),
    .Y(_06265_),
    .A1(net4720),
    .A2(net7434));
 sg13g2_a21oi_1 _28353_ (.A1(_14024_),
    .A2(net7434),
    .Y(_01627_),
    .B1(_06265_));
 sg13g2_nand4_1 _28354_ (.B(_14013_),
    .C(_14019_),
    .A(_14006_),
    .Y(_06266_),
    .D(_14029_));
 sg13g2_nand2b_1 _28355_ (.Y(_06267_),
    .B(net8550),
    .A_N(net8611));
 sg13g2_nand3_1 _28356_ (.B(_13977_),
    .C(_13985_),
    .A(net8666),
    .Y(_06268_));
 sg13g2_nor4_1 _28357_ (.A(net8613),
    .B(net8609),
    .C(_06267_),
    .D(_06268_),
    .Y(_06269_));
 sg13g2_nor4_1 _28358_ (.A(_13979_),
    .B(net8607),
    .C(net8605),
    .D(_14025_),
    .Y(_06270_));
 sg13g2_nand4_1 _28359_ (.B(_14001_),
    .C(_06269_),
    .A(_13994_),
    .Y(_06271_),
    .D(_06270_));
 sg13g2_nor4_2 _28360_ (.A(_13134_),
    .B(_13146_),
    .C(_06266_),
    .Y(_06272_),
    .D(_06271_));
 sg13g2_nand4_1 _28361_ (.B(_13123_),
    .C(_13150_),
    .A(_12510_),
    .Y(_06273_),
    .D(_06272_));
 sg13g2_o21ai_1 _28362_ (.B1(net1),
    .Y(_06274_),
    .A1(net7468),
    .A2(_06273_));
 sg13g2_nor2b_2 _28363_ (.A(net9306),
    .B_N(net2794),
    .Y(_06275_));
 sg13g2_nor2_1 _28364_ (.A(net9005),
    .B(net2794),
    .Y(_06276_));
 sg13g2_nor3_1 _28365_ (.A(_06274_),
    .B(_06275_),
    .C(_06276_),
    .Y(_01628_));
 sg13g2_xnor2_1 _28366_ (.Y(_06277_),
    .A(net4480),
    .B(_06275_));
 sg13g2_nor2_1 _28367_ (.A(_06274_),
    .B(_06277_),
    .Y(_01629_));
 sg13g2_nand3_1 _28368_ (.B(net5065),
    .C(_06275_),
    .A(net4480),
    .Y(_06278_));
 sg13g2_a21oi_1 _28369_ (.A1(net4480),
    .A2(_06275_),
    .Y(_06279_),
    .B1(net5065));
 sg13g2_nor2_1 _28370_ (.A(_06274_),
    .B(_06279_),
    .Y(_06280_));
 sg13g2_and2_1 _28371_ (.A(_06278_),
    .B(_06280_),
    .X(_01630_));
 sg13g2_a21oi_1 _28372_ (.A1(net9005),
    .A2(_06278_),
    .Y(_01631_),
    .B1(_06274_));
 sg13g2_o21ai_1 _28373_ (.B1(net9321),
    .Y(_06281_),
    .A1(\soc_I.clint_I.mtime[0] ),
    .A2(_06221_));
 sg13g2_nor2_1 _28374_ (.A(net3910),
    .B(_06207_),
    .Y(_06282_));
 sg13g2_nor2_1 _28375_ (.A(_06281_),
    .B(_06282_),
    .Y(_01632_));
 sg13g2_a21oi_1 _28376_ (.A1(\soc_I.clint_I.mtime[0] ),
    .A2(_06221_),
    .Y(_06283_),
    .B1(net3783));
 sg13g2_nor3_2 _28377_ (.A(_10444_),
    .B(_10445_),
    .C(_06185_),
    .Y(_06284_));
 sg13g2_nor3_1 _28378_ (.A(_10444_),
    .B(_10445_),
    .C(_06207_),
    .Y(_06285_));
 sg13g2_nor3_1 _28379_ (.A(net9014),
    .B(net3784),
    .C(_06285_),
    .Y(_01633_));
 sg13g2_or2_1 _28380_ (.X(_06286_),
    .B(_06284_),
    .A(net5515));
 sg13g2_nand4_1 _28381_ (.B(net3783),
    .C(\soc_I.clint_I.mtime[0] ),
    .A(net5515),
    .Y(_06287_),
    .D(_06221_));
 sg13g2_and3_1 _28382_ (.X(_01634_),
    .A(net9311),
    .B(_06286_),
    .C(_06287_));
 sg13g2_nor2b_1 _28383_ (.A(_00122_),
    .B_N(_06284_),
    .Y(_06288_));
 sg13g2_o21ai_1 _28384_ (.B1(net9311),
    .Y(_06289_),
    .A1(net3694),
    .A2(_06288_));
 sg13g2_a21oi_1 _28385_ (.A1(net3694),
    .A2(_06288_),
    .Y(_01635_),
    .B1(_06289_));
 sg13g2_nand3_1 _28386_ (.B(\soc_I.clint_I.mtime[2] ),
    .C(_06284_),
    .A(net3694),
    .Y(_06290_));
 sg13g2_nor2_1 _28387_ (.A(_10443_),
    .B(_06287_),
    .Y(_06291_));
 sg13g2_o21ai_1 _28388_ (.B1(net9310),
    .Y(_06292_),
    .A1(_10442_),
    .A2(_06290_));
 sg13g2_nand4_1 _28389_ (.B(\soc_I.clint_I.mtime[3] ),
    .C(\soc_I.clint_I.mtime[2] ),
    .A(\soc_I.clint_I.mtime[4] ),
    .Y(_06293_),
    .D(_06285_));
 sg13g2_a21oi_1 _28390_ (.A1(_10442_),
    .A2(_06290_),
    .Y(_01636_),
    .B1(_06292_));
 sg13g2_nor2_1 _28391_ (.A(_00132_),
    .B(_06290_),
    .Y(_06294_));
 sg13g2_o21ai_1 _28392_ (.B1(net9311),
    .Y(_06295_),
    .A1(net3593),
    .A2(_06294_));
 sg13g2_a21oi_1 _28393_ (.A1(net3593),
    .A2(_06294_),
    .Y(_01637_),
    .B1(_06295_));
 sg13g2_or3_1 _28394_ (.A(_10441_),
    .B(_10442_),
    .C(_06290_),
    .X(_06296_));
 sg13g2_nor2_1 _28395_ (.A(_10441_),
    .B(_10442_),
    .Y(_06297_));
 sg13g2_a21oi_1 _28396_ (.A1(_06291_),
    .A2(_06297_),
    .Y(_06298_),
    .B1(net3799));
 sg13g2_nor2_1 _28397_ (.A(_10440_),
    .B(_06296_),
    .Y(_06299_));
 sg13g2_nor3_1 _28398_ (.A(net9006),
    .B(net3800),
    .C(_06299_),
    .Y(_01638_));
 sg13g2_nor2_1 _28399_ (.A(_00142_),
    .B(_06296_),
    .Y(_06300_));
 sg13g2_o21ai_1 _28400_ (.B1(net9308),
    .Y(_06301_),
    .A1(net3413),
    .A2(_06300_));
 sg13g2_a21oi_1 _28401_ (.A1(net3413),
    .A2(_06300_),
    .Y(_01639_),
    .B1(_06301_));
 sg13g2_nor3_2 _28402_ (.A(_10439_),
    .B(_10440_),
    .C(_06296_),
    .Y(_06302_));
 sg13g2_nor4_1 _28403_ (.A(_10439_),
    .B(_10440_),
    .C(_10441_),
    .D(_06293_),
    .Y(_06303_));
 sg13g2_nand4_1 _28404_ (.B(net3799),
    .C(_06291_),
    .A(net3413),
    .Y(_06304_),
    .D(_06297_));
 sg13g2_nand2_2 _28405_ (.Y(_06305_),
    .A(net5087),
    .B(_06302_));
 sg13g2_nand2_1 _28406_ (.Y(_06306_),
    .A(net9308),
    .B(_06305_));
 sg13g2_a21oi_1 _28407_ (.A1(_10438_),
    .A2(_06304_),
    .Y(_01640_),
    .B1(_06306_));
 sg13g2_nor2b_1 _28408_ (.A(_00077_),
    .B_N(_06302_),
    .Y(_06307_));
 sg13g2_o21ai_1 _28409_ (.B1(net9308),
    .Y(_06308_),
    .A1(net4332),
    .A2(_06307_));
 sg13g2_a21oi_1 _28410_ (.A1(net4332),
    .A2(_06307_),
    .Y(_01641_),
    .B1(_06308_));
 sg13g2_nor2_1 _28411_ (.A(_10437_),
    .B(_06305_),
    .Y(_06309_));
 sg13g2_nand3_1 _28412_ (.B(\soc_I.clint_I.mtime[8] ),
    .C(_06303_),
    .A(\soc_I.clint_I.mtime[9] ),
    .Y(_06310_));
 sg13g2_nor2_1 _28413_ (.A(net5125),
    .B(_06309_),
    .Y(_06311_));
 sg13g2_nand2_1 _28414_ (.Y(_06312_),
    .A(\soc_I.clint_I.mtime[10] ),
    .B(_06309_));
 sg13g2_nor4_2 _28415_ (.A(_10436_),
    .B(_10437_),
    .C(_10438_),
    .Y(_06313_),
    .D(_06304_));
 sg13g2_nor3_1 _28416_ (.A(net9004),
    .B(_06311_),
    .C(_06313_),
    .Y(_01642_));
 sg13g2_nor3_1 _28417_ (.A(_10437_),
    .B(_00085_),
    .C(_06305_),
    .Y(_06314_));
 sg13g2_o21ai_1 _28418_ (.B1(net9300),
    .Y(_06315_),
    .A1(net4518),
    .A2(_06314_));
 sg13g2_a21oi_1 _28419_ (.A1(net4518),
    .A2(_06314_),
    .Y(_01643_),
    .B1(_06315_));
 sg13g2_nor3_2 _28420_ (.A(_10435_),
    .B(_10436_),
    .C(_06310_),
    .Y(_06316_));
 sg13g2_nand4_1 _28421_ (.B(\soc_I.clint_I.mtime[11] ),
    .C(\soc_I.clint_I.mtime[10] ),
    .A(\soc_I.clint_I.mtime[12] ),
    .Y(_06317_),
    .D(_06309_));
 sg13g2_o21ai_1 _28422_ (.B1(net9301),
    .Y(_06318_),
    .A1(net5188),
    .A2(_06316_));
 sg13g2_a21oi_1 _28423_ (.A1(net5188),
    .A2(_06316_),
    .Y(_01644_),
    .B1(_06318_));
 sg13g2_nor3_1 _28424_ (.A(_10435_),
    .B(net4501),
    .C(_06312_),
    .Y(_06319_));
 sg13g2_o21ai_1 _28425_ (.B1(net9301),
    .Y(_06320_),
    .A1(\soc_I.clint_I.mtime[13] ),
    .A2(net4502));
 sg13g2_a21oi_1 _28426_ (.A1(\soc_I.clint_I.mtime[13] ),
    .A2(net4502),
    .Y(_01645_),
    .B1(_06320_));
 sg13g2_nor2_1 _28427_ (.A(_10434_),
    .B(_06317_),
    .Y(_06321_));
 sg13g2_nand3_1 _28428_ (.B(net5188),
    .C(_06316_),
    .A(\soc_I.clint_I.mtime[13] ),
    .Y(_06322_));
 sg13g2_and4_1 _28429_ (.A(\soc_I.clint_I.mtime[13] ),
    .B(\soc_I.clint_I.mtime[12] ),
    .C(\soc_I.clint_I.mtime[11] ),
    .D(_06313_),
    .X(_06323_));
 sg13g2_nand2_1 _28430_ (.Y(_06324_),
    .A(net5243),
    .B(_06321_));
 sg13g2_nand2_1 _28431_ (.Y(_06325_),
    .A(net9316),
    .B(_06324_));
 sg13g2_a21oi_1 _28432_ (.A1(_10433_),
    .A2(_06322_),
    .Y(_01646_),
    .B1(_06325_));
 sg13g2_nor3_1 _28433_ (.A(_10434_),
    .B(_00101_),
    .C(_06317_),
    .Y(_06326_));
 sg13g2_o21ai_1 _28434_ (.B1(net9301),
    .Y(_06327_),
    .A1(net4602),
    .A2(_06326_));
 sg13g2_a21oi_1 _28435_ (.A1(net4602),
    .A2(_06326_),
    .Y(_01647_),
    .B1(_06327_));
 sg13g2_nor3_1 _28436_ (.A(_10432_),
    .B(_10433_),
    .C(_06322_),
    .Y(_06328_));
 sg13g2_nand3_1 _28437_ (.B(net5243),
    .C(_06323_),
    .A(net4602),
    .Y(_06329_));
 sg13g2_nand2b_1 _28438_ (.Y(_06330_),
    .B(_06329_),
    .A_N(net5428));
 sg13g2_nand4_1 _28439_ (.B(\soc_I.clint_I.mtime[15] ),
    .C(\soc_I.clint_I.mtime[14] ),
    .A(\soc_I.clint_I.mtime[16] ),
    .Y(_06331_),
    .D(_06321_));
 sg13g2_and3_1 _28440_ (.X(_01648_),
    .A(net9316),
    .B(_06330_),
    .C(_06331_));
 sg13g2_nor3_1 _28441_ (.A(_10432_),
    .B(_00015_),
    .C(_06324_),
    .Y(_06332_));
 sg13g2_o21ai_1 _28442_ (.B1(net9316),
    .Y(_06333_),
    .A1(net4497),
    .A2(_06332_));
 sg13g2_a21oi_1 _28443_ (.A1(net4497),
    .A2(_06332_),
    .Y(_01649_),
    .B1(_06333_));
 sg13g2_nand3_1 _28444_ (.B(\soc_I.clint_I.mtime[16] ),
    .C(_06328_),
    .A(net4497),
    .Y(_06334_));
 sg13g2_nand2_1 _28445_ (.Y(_06335_),
    .A(\soc_I.clint_I.mtime[17] ),
    .B(\soc_I.clint_I.mtime[16] ));
 sg13g2_nor3_1 _28446_ (.A(_10430_),
    .B(_06329_),
    .C(_06335_),
    .Y(_06336_));
 sg13g2_a21o_1 _28447_ (.A2(_06334_),
    .A1(_10430_),
    .B1(_06336_),
    .X(_06337_));
 sg13g2_nor2_1 _28448_ (.A(net9009),
    .B(net5391),
    .Y(_01650_));
 sg13g2_nor3_1 _28449_ (.A(_10431_),
    .B(_00030_),
    .C(_06331_),
    .Y(_06338_));
 sg13g2_o21ai_1 _28450_ (.B1(net9317),
    .Y(_06339_),
    .A1(net3943),
    .A2(_06338_));
 sg13g2_a21oi_1 _28451_ (.A1(net3943),
    .A2(_06338_),
    .Y(_01651_),
    .B1(_06339_));
 sg13g2_nor4_2 _28452_ (.A(_10429_),
    .B(_10430_),
    .C(_10431_),
    .Y(_06340_),
    .D(_06331_));
 sg13g2_and2_1 _28453_ (.A(net3943),
    .B(_06336_),
    .X(_06341_));
 sg13g2_nor4_1 _28454_ (.A(_10428_),
    .B(_10429_),
    .C(_10430_),
    .D(_06334_),
    .Y(_06342_));
 sg13g2_o21ai_1 _28455_ (.B1(net9317),
    .Y(_06343_),
    .A1(net5119),
    .A2(_06341_));
 sg13g2_nor2_1 _28456_ (.A(_06342_),
    .B(_06343_),
    .Y(_01652_));
 sg13g2_and2_1 _28457_ (.A(_10662_),
    .B(_06340_),
    .X(_06344_));
 sg13g2_o21ai_1 _28458_ (.B1(net9318),
    .Y(_06345_),
    .A1(net5003),
    .A2(_06344_));
 sg13g2_a21oi_1 _28459_ (.A1(net5003),
    .A2(_06344_),
    .Y(_01653_),
    .B1(_06345_));
 sg13g2_and3_1 _28460_ (.X(_06346_),
    .A(\soc_I.clint_I.mtime[21] ),
    .B(\soc_I.clint_I.mtime[20] ),
    .C(_06340_));
 sg13g2_and2_1 _28461_ (.A(\soc_I.clint_I.mtime[21] ),
    .B(\soc_I.clint_I.mtime[20] ),
    .X(_06347_));
 sg13g2_or2_1 _28462_ (.X(_06348_),
    .B(_06346_),
    .A(net5511));
 sg13g2_nand2_1 _28463_ (.Y(_06349_),
    .A(net5511),
    .B(_06346_));
 sg13g2_and3_1 _28464_ (.X(_01654_),
    .A(net9318),
    .B(_06348_),
    .C(_06349_));
 sg13g2_and2_1 _28465_ (.A(_10666_),
    .B(_06346_),
    .X(_06350_));
 sg13g2_o21ai_1 _28466_ (.B1(net9318),
    .Y(_06351_),
    .A1(\soc_I.clint_I.mtime[23] ),
    .A2(_06350_));
 sg13g2_a21oi_1 _28467_ (.A1(\soc_I.clint_I.mtime[23] ),
    .A2(_06350_),
    .Y(_01655_),
    .B1(_06351_));
 sg13g2_nand4_1 _28468_ (.B(\soc_I.clint_I.mtime[22] ),
    .C(net5003),
    .A(\soc_I.clint_I.mtime[23] ),
    .Y(_06352_),
    .D(_06342_));
 sg13g2_nand4_1 _28469_ (.B(\soc_I.clint_I.mtime[22] ),
    .C(_06341_),
    .A(\soc_I.clint_I.mtime[23] ),
    .Y(_06353_),
    .D(_06347_));
 sg13g2_nor3_1 _28470_ (.A(_10426_),
    .B(_10427_),
    .C(_06349_),
    .Y(_06354_));
 sg13g2_xnor2_1 _28471_ (.Y(_06355_),
    .A(_10426_),
    .B(_06353_));
 sg13g2_nor2_1 _28472_ (.A(net9008),
    .B(net5298),
    .Y(_01656_));
 sg13g2_nor3_1 _28473_ (.A(_10427_),
    .B(net4171),
    .C(_06349_),
    .Y(_06356_));
 sg13g2_o21ai_1 _28474_ (.B1(net9318),
    .Y(_06357_),
    .A1(\soc_I.clint_I.mtime[25] ),
    .A2(net4172));
 sg13g2_a21oi_1 _28475_ (.A1(\soc_I.clint_I.mtime[25] ),
    .A2(net4172),
    .Y(_01657_),
    .B1(_06357_));
 sg13g2_and2_1 _28476_ (.A(\soc_I.clint_I.mtime[25] ),
    .B(_06354_),
    .X(_06358_));
 sg13g2_nand2_1 _28477_ (.Y(_06359_),
    .A(\soc_I.clint_I.mtime[25] ),
    .B(_06354_));
 sg13g2_nor4_2 _28478_ (.A(_10424_),
    .B(_10425_),
    .C(_10426_),
    .Y(_06360_),
    .D(_06352_));
 sg13g2_o21ai_1 _28479_ (.B1(net9317),
    .Y(_06361_),
    .A1(net5194),
    .A2(_06358_));
 sg13g2_nor4_1 _28480_ (.A(_10424_),
    .B(_10425_),
    .C(_10426_),
    .D(_06353_),
    .Y(_06362_));
 sg13g2_nor2_1 _28481_ (.A(_06360_),
    .B(net5195),
    .Y(_01658_));
 sg13g2_nor2_1 _28482_ (.A(_00034_),
    .B(_06359_),
    .Y(_06363_));
 sg13g2_o21ai_1 _28483_ (.B1(net9319),
    .Y(_06364_),
    .A1(net4901),
    .A2(_06363_));
 sg13g2_a21oi_1 _28484_ (.A1(net4901),
    .A2(_06363_),
    .Y(_01659_),
    .B1(_06364_));
 sg13g2_and3_1 _28485_ (.X(_06365_),
    .A(\soc_I.clint_I.mtime[27] ),
    .B(\soc_I.clint_I.mtime[26] ),
    .C(_06358_));
 sg13g2_or2_1 _28486_ (.X(_06366_),
    .B(_06365_),
    .A(net5474));
 sg13g2_nand2_1 _28487_ (.Y(_06367_),
    .A(net5474),
    .B(_06365_));
 sg13g2_and3_1 _28488_ (.X(_01660_),
    .A(net9326),
    .B(net5475),
    .C(_06367_));
 sg13g2_nor2b_1 _28489_ (.A(_00048_),
    .B_N(_06365_),
    .Y(_06368_));
 sg13g2_o21ai_1 _28490_ (.B1(net9322),
    .Y(_06369_),
    .A1(net4555),
    .A2(_06368_));
 sg13g2_a21oi_1 _28491_ (.A1(net4555),
    .A2(_06368_),
    .Y(_01661_),
    .B1(_06369_));
 sg13g2_nand4_1 _28492_ (.B(net5474),
    .C(net4901),
    .A(net4555),
    .Y(_06370_),
    .D(_06360_));
 sg13g2_and4_1 _28493_ (.A(net4555),
    .B(\soc_I.clint_I.mtime[28] ),
    .C(\soc_I.clint_I.mtime[27] ),
    .D(_06362_),
    .X(_06371_));
 sg13g2_nor3_1 _28494_ (.A(_10422_),
    .B(_10423_),
    .C(_06367_),
    .Y(_06372_));
 sg13g2_xnor2_1 _28495_ (.Y(_06373_),
    .A(net4765),
    .B(_06371_));
 sg13g2_nor2_1 _28496_ (.A(net9008),
    .B(net4766),
    .Y(_01662_));
 sg13g2_nor3_1 _28497_ (.A(_10423_),
    .B(_00064_),
    .C(_06367_),
    .Y(_06374_));
 sg13g2_o21ai_1 _28498_ (.B1(net9322),
    .Y(_06375_),
    .A1(net4582),
    .A2(_06374_));
 sg13g2_a21oi_1 _28499_ (.A1(net4582),
    .A2(_06374_),
    .Y(_01663_),
    .B1(_06375_));
 sg13g2_nand3_1 _28500_ (.B(net4765),
    .C(_06371_),
    .A(net4582),
    .Y(_06376_));
 sg13g2_and2_1 _28501_ (.A(_10420_),
    .B(_06376_),
    .X(_06377_));
 sg13g2_nor4_2 _28502_ (.A(_10420_),
    .B(_10421_),
    .C(_10422_),
    .Y(_06378_),
    .D(_06370_));
 sg13g2_nor3_1 _28503_ (.A(net9008),
    .B(_06377_),
    .C(net5510),
    .Y(_01664_));
 sg13g2_nor2_1 _28504_ (.A(net4494),
    .B(_06376_),
    .Y(_06379_));
 sg13g2_o21ai_1 _28505_ (.B1(net9322),
    .Y(_06380_),
    .A1(\soc_I.clint_I.mtime[33] ),
    .A2(net4495));
 sg13g2_a21oi_1 _28506_ (.A1(\soc_I.clint_I.mtime[33] ),
    .A2(net4495),
    .Y(_01665_),
    .B1(_06380_));
 sg13g2_nand4_1 _28507_ (.B(net4996),
    .C(net4582),
    .A(\soc_I.clint_I.mtime[33] ),
    .Y(_06381_),
    .D(_06372_));
 sg13g2_nand3_1 _28508_ (.B(\soc_I.clint_I.mtime[33] ),
    .C(_06378_),
    .A(net5536),
    .Y(_06382_));
 sg13g2_nand2_1 _28509_ (.Y(_06383_),
    .A(net9320),
    .B(_06382_));
 sg13g2_a21oi_1 _28510_ (.A1(_10419_),
    .A2(net4997),
    .Y(_01666_),
    .B1(_06383_));
 sg13g2_nor3_1 _28511_ (.A(_10418_),
    .B(_10419_),
    .C(_06381_),
    .Y(_06384_));
 sg13g2_nor2_1 _28512_ (.A(_10418_),
    .B(_06382_),
    .Y(_06385_));
 sg13g2_a21oi_1 _28513_ (.A1(_10418_),
    .A2(_06382_),
    .Y(_06386_),
    .B1(net9008));
 sg13g2_nor2b_1 _28514_ (.A(_06385_),
    .B_N(net5537),
    .Y(_01667_));
 sg13g2_o21ai_1 _28515_ (.B1(_10417_),
    .Y(_06387_),
    .A1(_10418_),
    .A2(_06382_));
 sg13g2_nand2_2 _28516_ (.Y(_06388_),
    .A(net5546),
    .B(_06385_));
 sg13g2_and3_1 _28517_ (.X(_01668_),
    .A(net9320),
    .B(_06387_),
    .C(_06388_));
 sg13g2_nand3_1 _28518_ (.B(\soc_I.clint_I.mtime[36] ),
    .C(_06384_),
    .A(net5166),
    .Y(_06389_));
 sg13g2_nand2_1 _28519_ (.Y(_06390_),
    .A(net9320),
    .B(_06389_));
 sg13g2_a21oi_1 _28520_ (.A1(_10416_),
    .A2(_06388_),
    .Y(_01669_),
    .B1(_06390_));
 sg13g2_and2_1 _28521_ (.A(_10415_),
    .B(_06389_),
    .X(_06391_));
 sg13g2_nor3_2 _28522_ (.A(_10415_),
    .B(_10416_),
    .C(_06388_),
    .Y(_06392_));
 sg13g2_nor3_1 _28523_ (.A(net9004),
    .B(_06391_),
    .C(_06392_),
    .Y(_01670_));
 sg13g2_nor2_1 _28524_ (.A(net5061),
    .B(_06392_),
    .Y(_06393_));
 sg13g2_nor3_2 _28525_ (.A(_10414_),
    .B(_10415_),
    .C(_06389_),
    .Y(_06394_));
 sg13g2_nor3_1 _28526_ (.A(net9007),
    .B(net5062),
    .C(_06394_),
    .Y(_01671_));
 sg13g2_nor2_1 _28527_ (.A(net5149),
    .B(_06394_),
    .Y(_06395_));
 sg13g2_nand2_1 _28528_ (.Y(_06396_),
    .A(net5149),
    .B(_06394_));
 sg13g2_inv_1 _28529_ (.Y(_06397_),
    .A(_06396_));
 sg13g2_nor3_1 _28530_ (.A(net9003),
    .B(net5150),
    .C(_06397_),
    .Y(_01672_));
 sg13g2_and4_2 _28531_ (.A(net5317),
    .B(net5149),
    .C(\soc_I.clint_I.mtime[39] ),
    .D(_06392_),
    .X(_06398_));
 sg13g2_o21ai_1 _28532_ (.B1(net9305),
    .Y(_06399_),
    .A1(net5317),
    .A2(_06397_));
 sg13g2_nor2_1 _28533_ (.A(_06398_),
    .B(_06399_),
    .Y(_01673_));
 sg13g2_nor2_1 _28534_ (.A(net5117),
    .B(_06398_),
    .Y(_06400_));
 sg13g2_and3_1 _28535_ (.X(_06401_),
    .A(net5117),
    .B(\soc_I.clint_I.mtime[41] ),
    .C(_06397_));
 sg13g2_nor3_1 _28536_ (.A(net9003),
    .B(_06400_),
    .C(_06401_),
    .Y(_01674_));
 sg13g2_or2_1 _28537_ (.X(_06402_),
    .B(_06401_),
    .A(net5169));
 sg13g2_nand2_2 _28538_ (.Y(_06403_),
    .A(net5169),
    .B(_06401_));
 sg13g2_and3_1 _28539_ (.X(_01675_),
    .A(net9300),
    .B(_06402_),
    .C(_06403_));
 sg13g2_nand4_1 _28540_ (.B(\soc_I.clint_I.mtime[43] ),
    .C(\soc_I.clint_I.mtime[42] ),
    .A(\soc_I.clint_I.mtime[44] ),
    .Y(_06404_),
    .D(_06398_));
 sg13g2_nand2_1 _28541_ (.Y(_06405_),
    .A(net9300),
    .B(_06404_));
 sg13g2_a21oi_1 _28542_ (.A1(_10413_),
    .A2(_06403_),
    .Y(_01676_),
    .B1(_06405_));
 sg13g2_and2_1 _28543_ (.A(_10412_),
    .B(_06404_),
    .X(_06406_));
 sg13g2_nor3_2 _28544_ (.A(_10412_),
    .B(_10413_),
    .C(_06403_),
    .Y(_06407_));
 sg13g2_nor3_1 _28545_ (.A(net9004),
    .B(net5499),
    .C(_06407_),
    .Y(_01677_));
 sg13g2_o21ai_1 _28546_ (.B1(_10411_),
    .Y(_06408_),
    .A1(_10412_),
    .A2(_06404_));
 sg13g2_nand2_1 _28547_ (.Y(_06409_),
    .A(net5552),
    .B(_06407_));
 sg13g2_and3_1 _28548_ (.X(_01678_),
    .A(net9301),
    .B(_06408_),
    .C(_06409_));
 sg13g2_a21oi_1 _28549_ (.A1(\soc_I.clint_I.mtime[46] ),
    .A2(_06407_),
    .Y(_06410_),
    .B1(net4001));
 sg13g2_nor4_2 _28550_ (.A(_10410_),
    .B(_10411_),
    .C(_10412_),
    .Y(_06411_),
    .D(_06404_));
 sg13g2_nor3_1 _28551_ (.A(net9004),
    .B(net4002),
    .C(_06411_),
    .Y(_01679_));
 sg13g2_nor2_1 _28552_ (.A(net5079),
    .B(_06411_),
    .Y(_06412_));
 sg13g2_nor3_2 _28553_ (.A(_10409_),
    .B(_10410_),
    .C(_06409_),
    .Y(_06413_));
 sg13g2_nor3_1 _28554_ (.A(net9004),
    .B(_06412_),
    .C(_06413_),
    .Y(_01680_));
 sg13g2_or2_1 _28555_ (.X(_06414_),
    .B(_06413_),
    .A(net5444));
 sg13g2_nand2_1 _28556_ (.Y(_06415_),
    .A(net5444),
    .B(_06413_));
 sg13g2_and3_1 _28557_ (.X(_01681_),
    .A(net9315),
    .B(_06414_),
    .C(_06415_));
 sg13g2_nand2b_1 _28558_ (.Y(_06416_),
    .B(_06415_),
    .A_N(net5174));
 sg13g2_nand4_1 _28559_ (.B(\soc_I.clint_I.mtime[49] ),
    .C(net5079),
    .A(net5174),
    .Y(_06417_),
    .D(_06411_));
 sg13g2_and3_1 _28560_ (.X(_01682_),
    .A(net9315),
    .B(_06416_),
    .C(_06417_));
 sg13g2_nor2b_1 _28561_ (.A(net4819),
    .B_N(_06417_),
    .Y(_06418_));
 sg13g2_and4_2 _28562_ (.A(net4819),
    .B(\soc_I.clint_I.mtime[50] ),
    .C(\soc_I.clint_I.mtime[49] ),
    .D(_06413_),
    .X(_06419_));
 sg13g2_nor3_1 _28563_ (.A(net9009),
    .B(net4820),
    .C(net5175),
    .Y(_01683_));
 sg13g2_nor2_1 _28564_ (.A(net4721),
    .B(_06419_),
    .Y(_06420_));
 sg13g2_nand2_2 _28565_ (.Y(_06421_),
    .A(net4721),
    .B(net5175));
 sg13g2_inv_1 _28566_ (.Y(_06422_),
    .A(_06421_));
 sg13g2_nor3_1 _28567_ (.A(net9012),
    .B(net4722),
    .C(_06422_),
    .Y(_01684_));
 sg13g2_o21ai_1 _28568_ (.B1(net9318),
    .Y(_06423_),
    .A1(_10407_),
    .A2(_06421_));
 sg13g2_a21oi_1 _28569_ (.A1(_10407_),
    .A2(_06421_),
    .Y(_01685_),
    .B1(_06423_));
 sg13g2_a21oi_1 _28570_ (.A1(\soc_I.clint_I.mtime[53] ),
    .A2(_06422_),
    .Y(_06424_),
    .B1(net4274));
 sg13g2_nor3_2 _28571_ (.A(_10406_),
    .B(_10407_),
    .C(_06421_),
    .Y(_06425_));
 sg13g2_nor3_1 _28572_ (.A(net9012),
    .B(net4275),
    .C(_06425_),
    .Y(_01686_));
 sg13g2_nor2_1 _28573_ (.A(net4971),
    .B(_06425_),
    .Y(_06426_));
 sg13g2_nand2_2 _28574_ (.Y(_06427_),
    .A(net4971),
    .B(_06425_));
 sg13g2_inv_1 _28575_ (.Y(_06428_),
    .A(_06427_));
 sg13g2_nor3_1 _28576_ (.A(net9010),
    .B(_06426_),
    .C(_06428_),
    .Y(_01687_));
 sg13g2_o21ai_1 _28577_ (.B1(net9319),
    .Y(_06429_),
    .A1(_10405_),
    .A2(_06427_));
 sg13g2_a21oi_1 _28578_ (.A1(_10405_),
    .A2(_06427_),
    .Y(_01688_),
    .B1(_06429_));
 sg13g2_a21oi_1 _28579_ (.A1(\soc_I.clint_I.mtime[56] ),
    .A2(_06428_),
    .Y(_06430_),
    .B1(net4268));
 sg13g2_nor3_2 _28580_ (.A(_10404_),
    .B(_10405_),
    .C(_06427_),
    .Y(_06431_));
 sg13g2_nor3_1 _28581_ (.A(net9010),
    .B(net4269),
    .C(_06431_),
    .Y(_01689_));
 sg13g2_nor2_1 _28582_ (.A(net4825),
    .B(_06431_),
    .Y(_06432_));
 sg13g2_nand2_2 _28583_ (.Y(_06433_),
    .A(net4825),
    .B(_06431_));
 sg13g2_inv_1 _28584_ (.Y(_06434_),
    .A(_06433_));
 sg13g2_nor3_1 _28585_ (.A(net9011),
    .B(_06432_),
    .C(_06434_),
    .Y(_01690_));
 sg13g2_o21ai_1 _28586_ (.B1(net9319),
    .Y(_06435_),
    .A1(_10403_),
    .A2(_06433_));
 sg13g2_a21oi_1 _28587_ (.A1(_10403_),
    .A2(net4826),
    .Y(_01691_),
    .B1(_06435_));
 sg13g2_a21oi_1 _28588_ (.A1(\soc_I.clint_I.mtime[59] ),
    .A2(_06434_),
    .Y(_06436_),
    .B1(net4304));
 sg13g2_nor3_2 _28589_ (.A(_10402_),
    .B(_10403_),
    .C(_06433_),
    .Y(_06437_));
 sg13g2_nor3_1 _28590_ (.A(net9010),
    .B(net4305),
    .C(_06437_),
    .Y(_01692_));
 sg13g2_or2_1 _28591_ (.X(_06438_),
    .B(_06437_),
    .A(net5532));
 sg13g2_nand2_1 _28592_ (.Y(_06439_),
    .A(net5532),
    .B(_06437_));
 sg13g2_and3_1 _28593_ (.X(_01693_),
    .A(net9318),
    .B(_06438_),
    .C(_06439_));
 sg13g2_nand3_1 _28594_ (.B(\soc_I.clint_I.mtime[61] ),
    .C(_06437_),
    .A(net4564),
    .Y(_06440_));
 sg13g2_nand2_1 _28595_ (.Y(_06441_),
    .A(net9327),
    .B(_06440_));
 sg13g2_a21oi_1 _28596_ (.A1(_10400_),
    .A2(_06439_),
    .Y(_01694_),
    .B1(_06441_));
 sg13g2_o21ai_1 _28597_ (.B1(net9318),
    .Y(_06442_),
    .A1(_10399_),
    .A2(_06440_));
 sg13g2_a21oi_1 _28598_ (.A1(_10399_),
    .A2(_06440_),
    .Y(_01695_),
    .B1(_06442_));
 sg13g2_and3_2 _28599_ (.X(_06443_),
    .A(_13173_),
    .B(_13176_),
    .C(_14437_));
 sg13g2_and3_1 _28600_ (.X(_06444_),
    .A(_13173_),
    .B(_13260_),
    .C(_14437_));
 sg13g2_o21ai_1 _28601_ (.B1(net9331),
    .Y(_06445_),
    .A1(net4796),
    .A2(net7420));
 sg13g2_a21oi_1 _28602_ (.A1(_13978_),
    .A2(_06443_),
    .Y(_01696_),
    .B1(_06445_));
 sg13g2_o21ai_1 _28603_ (.B1(net9332),
    .Y(_06446_),
    .A1(net3405),
    .A2(_06444_));
 sg13g2_a21oi_1 _28604_ (.A1(net8612),
    .A2(_06443_),
    .Y(_01697_),
    .B1(_06446_));
 sg13g2_o21ai_1 _28605_ (.B1(net9331),
    .Y(_06447_),
    .A1(net4747),
    .A2(net7420));
 sg13g2_a21oi_1 _28606_ (.A1(net8610),
    .A2(_06443_),
    .Y(_01698_),
    .B1(_06447_));
 sg13g2_o21ai_1 _28607_ (.B1(net9331),
    .Y(_06448_),
    .A1(net4966),
    .A2(net7420));
 sg13g2_a21oi_1 _28608_ (.A1(net8549),
    .A2(net7420),
    .Y(_01699_),
    .B1(_06448_));
 sg13g2_o21ai_1 _28609_ (.B1(net9331),
    .Y(_06449_),
    .A1(net3918),
    .A2(_06444_));
 sg13g2_a21oi_1 _28610_ (.A1(net8608),
    .A2(_06443_),
    .Y(_01700_),
    .B1(_06449_));
 sg13g2_o21ai_1 _28611_ (.B1(net9332),
    .Y(_06450_),
    .A1(net3802),
    .A2(net7420));
 sg13g2_a21oi_1 _28612_ (.A1(net8606),
    .A2(_06443_),
    .Y(_01701_),
    .B1(_06450_));
 sg13g2_o21ai_1 _28613_ (.B1(net9331),
    .Y(_06451_),
    .A1(net4709),
    .A2(net7420));
 sg13g2_a21oi_1 _28614_ (.A1(net8604),
    .A2(_06443_),
    .Y(_01702_),
    .B1(_06451_));
 sg13g2_o21ai_1 _28615_ (.B1(net9332),
    .Y(_06452_),
    .A1(net4061),
    .A2(net7420));
 sg13g2_a21oi_1 _28616_ (.A1(_14024_),
    .A2(net7420),
    .Y(_01703_),
    .B1(_06452_));
 sg13g2_nor2_1 _28617_ (.A(net9016),
    .B(_13196_),
    .Y(_01704_));
 sg13g2_and3_2 _28618_ (.X(_06453_),
    .A(_13173_),
    .B(_13177_),
    .C(_14437_));
 sg13g2_and3_1 _28619_ (.X(_06454_),
    .A(_13173_),
    .B(_13261_),
    .C(_14437_));
 sg13g2_o21ai_1 _28620_ (.B1(net9331),
    .Y(_06455_),
    .A1(net4863),
    .A2(_06454_));
 sg13g2_a21oi_1 _28621_ (.A1(_13978_),
    .A2(_06453_),
    .Y(_01705_),
    .B1(_06455_));
 sg13g2_o21ai_1 _28622_ (.B1(net9334),
    .Y(_06456_),
    .A1(net4967),
    .A2(net7419));
 sg13g2_a21oi_1 _28623_ (.A1(net8612),
    .A2(_06453_),
    .Y(_01706_),
    .B1(_06456_));
 sg13g2_o21ai_1 _28624_ (.B1(net9331),
    .Y(_06457_),
    .A1(net5039),
    .A2(_06454_));
 sg13g2_a21oi_1 _28625_ (.A1(net8610),
    .A2(_06453_),
    .Y(_01707_),
    .B1(_06457_));
 sg13g2_o21ai_1 _28626_ (.B1(net9340),
    .Y(_06458_),
    .A1(net4892),
    .A2(net7419));
 sg13g2_a21oi_1 _28627_ (.A1(net8549),
    .A2(net7419),
    .Y(_01708_),
    .B1(_06458_));
 sg13g2_o21ai_1 _28628_ (.B1(net9334),
    .Y(_06459_),
    .A1(net5010),
    .A2(net7419));
 sg13g2_a21oi_1 _28629_ (.A1(net8608),
    .A2(_06453_),
    .Y(_01709_),
    .B1(_06459_));
 sg13g2_o21ai_1 _28630_ (.B1(net9332),
    .Y(_06460_),
    .A1(net4991),
    .A2(net7419));
 sg13g2_a21oi_1 _28631_ (.A1(net8606),
    .A2(_06453_),
    .Y(_01710_),
    .B1(_06460_));
 sg13g2_o21ai_1 _28632_ (.B1(net9340),
    .Y(_06461_),
    .A1(net4951),
    .A2(net7419));
 sg13g2_a21oi_1 _28633_ (.A1(net8604),
    .A2(_06453_),
    .Y(_01711_),
    .B1(_06461_));
 sg13g2_o21ai_1 _28634_ (.B1(net9331),
    .Y(_06462_),
    .A1(net5151),
    .A2(net7419));
 sg13g2_a21oi_1 _28635_ (.A1(_14024_),
    .A2(net7419),
    .Y(_01712_),
    .B1(_06462_));
 sg13g2_nor4_2 _28636_ (.A(_10466_),
    .B(net9710),
    .C(_00185_),
    .Y(_06463_),
    .D(_14128_));
 sg13g2_nand2_1 _28637_ (.Y(_06464_),
    .A(net8961),
    .B(_06463_));
 sg13g2_nand2_1 _28638_ (.Y(_06465_),
    .A(net2749),
    .B(net8106));
 sg13g2_o21ai_1 _28639_ (.B1(_06465_),
    .Y(_01713_),
    .A1(net7487),
    .A2(net8106));
 sg13g2_nand2_1 _28640_ (.Y(_06466_),
    .A(net3340),
    .B(net8103));
 sg13g2_o21ai_1 _28641_ (.B1(_06466_),
    .Y(_01714_),
    .A1(net7665),
    .A2(net8103));
 sg13g2_nand2_1 _28642_ (.Y(_06467_),
    .A(net2969),
    .B(net8105));
 sg13g2_o21ai_1 _28643_ (.B1(_06467_),
    .Y(_01715_),
    .A1(net7613),
    .A2(net8103));
 sg13g2_nand2_1 _28644_ (.Y(_06468_),
    .A(net3531),
    .B(net8105));
 sg13g2_o21ai_1 _28645_ (.B1(_06468_),
    .Y(_01716_),
    .A1(net7608),
    .A2(net8105));
 sg13g2_nand2_1 _28646_ (.Y(_06469_),
    .A(net3454),
    .B(net8101));
 sg13g2_o21ai_1 _28647_ (.B1(_06469_),
    .Y(_01717_),
    .A1(net7586),
    .A2(net8101));
 sg13g2_nand2_1 _28648_ (.Y(_06470_),
    .A(net2963),
    .B(net8101));
 sg13g2_o21ai_1 _28649_ (.B1(_06470_),
    .Y(_01718_),
    .A1(net7597),
    .A2(net8101));
 sg13g2_nand2_1 _28650_ (.Y(_06471_),
    .A(net3404),
    .B(net8104));
 sg13g2_o21ai_1 _28651_ (.B1(_06471_),
    .Y(_01719_),
    .A1(net7593),
    .A2(net8104));
 sg13g2_nand2_1 _28652_ (.Y(_06472_),
    .A(net3141),
    .B(net8099));
 sg13g2_o21ai_1 _28653_ (.B1(_06472_),
    .Y(_01720_),
    .A1(net7604),
    .A2(net8099));
 sg13g2_nand2_1 _28654_ (.Y(_06473_),
    .A(net3064),
    .B(net8102));
 sg13g2_o21ai_1 _28655_ (.B1(_06473_),
    .Y(_01721_),
    .A1(net7560),
    .A2(net8102));
 sg13g2_nand2_1 _28656_ (.Y(_06474_),
    .A(net2944),
    .B(net8105));
 sg13g2_o21ai_1 _28657_ (.B1(_06474_),
    .Y(_01722_),
    .A1(net7578),
    .A2(net8103));
 sg13g2_nand2_1 _28658_ (.Y(_06475_),
    .A(net2971),
    .B(net8104));
 sg13g2_o21ai_1 _28659_ (.B1(_06475_),
    .Y(_01723_),
    .A1(net7547),
    .A2(net8104));
 sg13g2_nand2_1 _28660_ (.Y(_06476_),
    .A(net4023),
    .B(net8097));
 sg13g2_o21ai_1 _28661_ (.B1(_06476_),
    .Y(_01724_),
    .A1(net7570),
    .A2(net8097));
 sg13g2_nand2_1 _28662_ (.Y(_06477_),
    .A(net3848),
    .B(net8103));
 sg13g2_o21ai_1 _28663_ (.B1(_06477_),
    .Y(_01725_),
    .A1(net7540),
    .A2(net8103));
 sg13g2_nand2_1 _28664_ (.Y(_06478_),
    .A(net3946),
    .B(net8103));
 sg13g2_o21ai_1 _28665_ (.B1(_06478_),
    .Y(_01726_),
    .A1(net7551),
    .A2(net8103));
 sg13g2_nand2_1 _28666_ (.Y(_06479_),
    .A(net3810),
    .B(net8107));
 sg13g2_o21ai_1 _28667_ (.B1(_06479_),
    .Y(_01727_),
    .A1(net7580),
    .A2(net8100));
 sg13g2_nand2_1 _28668_ (.Y(_06480_),
    .A(net3825),
    .B(net8097));
 sg13g2_o21ai_1 _28669_ (.B1(_06480_),
    .Y(_01728_),
    .A1(net7567),
    .A2(net8097));
 sg13g2_nand2_1 _28670_ (.Y(_06481_),
    .A(net3589),
    .B(net8097));
 sg13g2_o21ai_1 _28671_ (.B1(_06481_),
    .Y(_01729_),
    .A1(net7524),
    .A2(net8097));
 sg13g2_nand2_1 _28672_ (.Y(_06482_),
    .A(net2776),
    .B(net8097));
 sg13g2_o21ai_1 _28673_ (.B1(_06482_),
    .Y(_01730_),
    .A1(net7537),
    .A2(net8097));
 sg13g2_nand2_1 _28674_ (.Y(_06483_),
    .A(net3892),
    .B(net8099));
 sg13g2_o21ai_1 _28675_ (.B1(_06483_),
    .Y(_01731_),
    .A1(net7531),
    .A2(net8099));
 sg13g2_nand2_1 _28676_ (.Y(_06484_),
    .A(net3233),
    .B(net8099));
 sg13g2_o21ai_1 _28677_ (.B1(_06484_),
    .Y(_01732_),
    .A1(net7517),
    .A2(net8099));
 sg13g2_nand2_1 _28678_ (.Y(_06485_),
    .A(net3390),
    .B(net8106));
 sg13g2_o21ai_1 _28679_ (.B1(_06485_),
    .Y(_01733_),
    .A1(net7504),
    .A2(net8106));
 sg13g2_nand2_1 _28680_ (.Y(_06486_),
    .A(net3448),
    .B(net8101));
 sg13g2_o21ai_1 _28681_ (.B1(_06486_),
    .Y(_01734_),
    .A1(net7512),
    .A2(net8101));
 sg13g2_nand2_1 _28682_ (.Y(_06487_),
    .A(net3201),
    .B(net8104));
 sg13g2_o21ai_1 _28683_ (.B1(_06487_),
    .Y(_01735_),
    .A1(net7494),
    .A2(net8104));
 sg13g2_nand2_1 _28684_ (.Y(_06488_),
    .A(net3679),
    .B(net8098));
 sg13g2_o21ai_1 _28685_ (.B1(_06488_),
    .Y(_01736_),
    .A1(net7502),
    .A2(net8098));
 sg13g2_nand2_1 _28686_ (.Y(_06489_),
    .A(net2958),
    .B(net8101));
 sg13g2_o21ai_1 _28687_ (.B1(_06489_),
    .Y(_01737_),
    .A1(net7646),
    .A2(net8101));
 sg13g2_nand2_1 _28688_ (.Y(_06490_),
    .A(net3325),
    .B(net8106));
 sg13g2_o21ai_1 _28689_ (.B1(_06490_),
    .Y(_01738_),
    .A1(net7649),
    .A2(net8106));
 sg13g2_nand2_1 _28690_ (.Y(_06491_),
    .A(net3186),
    .B(net8104));
 sg13g2_o21ai_1 _28691_ (.B1(_06491_),
    .Y(_01739_),
    .A1(net7657),
    .A2(net8104));
 sg13g2_nand2_1 _28692_ (.Y(_06492_),
    .A(net3586),
    .B(net8100));
 sg13g2_o21ai_1 _28693_ (.B1(_06492_),
    .Y(_01740_),
    .A1(net7662),
    .A2(net8100));
 sg13g2_nand2_1 _28694_ (.Y(_06493_),
    .A(net3246),
    .B(net8100));
 sg13g2_o21ai_1 _28695_ (.B1(_06493_),
    .Y(_01741_),
    .A1(net7637),
    .A2(net8100));
 sg13g2_nand2_1 _28696_ (.Y(_06494_),
    .A(net3831),
    .B(net8102));
 sg13g2_o21ai_1 _28697_ (.B1(_06494_),
    .Y(_01742_),
    .A1(net7626),
    .A2(net8102));
 sg13g2_nand2_1 _28698_ (.Y(_06495_),
    .A(net3386),
    .B(net8100));
 sg13g2_o21ai_1 _28699_ (.B1(_06495_),
    .Y(_01743_),
    .A1(net7623),
    .A2(net8100));
 sg13g2_nand2_1 _28700_ (.Y(_06496_),
    .A(net3175),
    .B(net8098));
 sg13g2_o21ai_1 _28701_ (.B1(_06496_),
    .Y(_01744_),
    .A1(net7631),
    .A2(net8098));
 sg13g2_nand2_2 _28702_ (.Y(_06497_),
    .A(net4771),
    .B(_13795_));
 sg13g2_inv_2 _28703_ (.Y(_06498_),
    .A(_06497_));
 sg13g2_nor3_2 _28704_ (.A(\soc_I.spi0_I.div[2] ),
    .B(\soc_I.spi0_I.div[1] ),
    .C(\soc_I.spi0_I.div[0] ),
    .Y(_06499_));
 sg13g2_nor2b_1 _28705_ (.A(\soc_I.spi0_I.div[3] ),
    .B_N(_06499_),
    .Y(_06500_));
 sg13g2_nor2b_1 _28706_ (.A(\soc_I.spi0_I.div[4] ),
    .B_N(_06500_),
    .Y(_06501_));
 sg13g2_nor2b_1 _28707_ (.A(\soc_I.spi0_I.div[5] ),
    .B_N(_06501_),
    .Y(_06502_));
 sg13g2_nor2b_2 _28708_ (.A(\soc_I.spi0_I.div[6] ),
    .B_N(_06502_),
    .Y(_06503_));
 sg13g2_nand2b_1 _28709_ (.Y(_06504_),
    .B(_06503_),
    .A_N(\soc_I.spi0_I.div[7] ));
 sg13g2_nor3_1 _28710_ (.A(\soc_I.spi0_I.div[9] ),
    .B(\soc_I.spi0_I.div[8] ),
    .C(_06504_),
    .Y(_06505_));
 sg13g2_nor2b_1 _28711_ (.A(\soc_I.spi0_I.div[10] ),
    .B_N(_06505_),
    .Y(_06506_));
 sg13g2_nand2b_1 _28712_ (.Y(_06507_),
    .B(_06506_),
    .A_N(\soc_I.spi0_I.div[11] ));
 sg13g2_nor3_1 _28713_ (.A(\soc_I.spi0_I.div[13] ),
    .B(\soc_I.spi0_I.div[12] ),
    .C(_06507_),
    .Y(_06508_));
 sg13g2_nor2b_1 _28714_ (.A(\soc_I.spi0_I.div[14] ),
    .B_N(_06508_),
    .Y(_06509_));
 sg13g2_nor2b_2 _28715_ (.A(\soc_I.spi0_I.div[15] ),
    .B_N(_06509_),
    .Y(_06510_));
 sg13g2_xnor2_1 _28716_ (.Y(_06511_),
    .A(\soc_I.spi0_I.div[14] ),
    .B(_06508_));
 sg13g2_nand3b_1 _28717_ (.B(_00288_),
    .C(_06506_),
    .Y(_06512_),
    .A_N(\soc_I.spi0_I.div[11] ));
 sg13g2_xor2_1 _28718_ (.B(_06512_),
    .A(\soc_I.spi0_I.div[13] ),
    .X(_06513_));
 sg13g2_xnor2_1 _28719_ (.Y(_06514_),
    .A(_00288_),
    .B(_06507_));
 sg13g2_xnor2_1 _28720_ (.Y(_06515_),
    .A(\soc_I.spi0_I.div[11] ),
    .B(_06506_));
 sg13g2_nor2_1 _28721_ (.A(\soc_I.spi0_I.tick_cnt[11] ),
    .B(_06515_),
    .Y(_06516_));
 sg13g2_nand2_1 _28722_ (.Y(_06517_),
    .A(\soc_I.spi0_I.tick_cnt[11] ),
    .B(_06515_));
 sg13g2_nand2b_1 _28723_ (.Y(_06518_),
    .B(\soc_I.spi0_I.div[15] ),
    .A_N(_06509_));
 sg13g2_nor2_1 _28724_ (.A(\soc_I.spi0_I.tick_cnt[13] ),
    .B(_06513_),
    .Y(_06519_));
 sg13g2_a21oi_1 _28725_ (.A1(\soc_I.spi0_I.tick_cnt[15] ),
    .A2(_06518_),
    .Y(_06520_),
    .B1(_06519_));
 sg13g2_xor2_1 _28726_ (.B(\soc_I.spi0_I.tick_cnt[9] ),
    .A(\soc_I.spi0_I.div[9] ),
    .X(_06521_));
 sg13g2_nand3b_1 _28727_ (.B(_00287_),
    .C(_06503_),
    .Y(_06522_),
    .A_N(\soc_I.spi0_I.div[7] ));
 sg13g2_xnor2_1 _28728_ (.Y(_06523_),
    .A(\soc_I.spi0_I.div[10] ),
    .B(_06505_));
 sg13g2_xnor2_1 _28729_ (.Y(_06524_),
    .A(\soc_I.spi0_I.div[7] ),
    .B(_06503_));
 sg13g2_xnor2_1 _28730_ (.Y(_06525_),
    .A(\soc_I.spi0_I.tick_cnt[7] ),
    .B(_06524_));
 sg13g2_xnor2_1 _28731_ (.Y(_06526_),
    .A(\soc_I.spi0_I.div[5] ),
    .B(_06501_));
 sg13g2_xnor2_1 _28732_ (.Y(_06527_),
    .A(\soc_I.spi0_I.tick_cnt[5] ),
    .B(_06526_));
 sg13g2_xor2_1 _28733_ (.B(\soc_I.spi0_I.div[0] ),
    .A(\soc_I.spi0_I.div[1] ),
    .X(_06528_));
 sg13g2_nor2_1 _28734_ (.A(\soc_I.spi0_I.div[0] ),
    .B(\soc_I.spi0_I.tick_cnt[0] ),
    .Y(_06529_));
 sg13g2_nor3_1 _28735_ (.A(\soc_I.spi0_I.tick_cnt[17] ),
    .B(\soc_I.spi0_I.tick_cnt[16] ),
    .C(_06529_),
    .Y(_06530_));
 sg13g2_o21ai_1 _28736_ (.B1(_06530_),
    .Y(_06531_),
    .A1(\soc_I.spi0_I.tick_cnt[1] ),
    .A2(_06528_));
 sg13g2_a221oi_1 _28737_ (.B2(\soc_I.spi0_I.tick_cnt[1] ),
    .C1(_06531_),
    .B1(_06528_),
    .A1(\soc_I.spi0_I.div[0] ),
    .Y(_06532_),
    .A2(\soc_I.spi0_I.tick_cnt[0] ));
 sg13g2_o21ai_1 _28738_ (.B1(\soc_I.spi0_I.div[2] ),
    .Y(_06533_),
    .A1(\soc_I.spi0_I.div[1] ),
    .A2(\soc_I.spi0_I.div[0] ));
 sg13g2_nand2b_1 _28739_ (.Y(_06534_),
    .B(_06533_),
    .A_N(_06499_));
 sg13g2_xnor2_1 _28740_ (.Y(_06535_),
    .A(\soc_I.spi0_I.tick_cnt[2] ),
    .B(_06534_));
 sg13g2_xor2_1 _28741_ (.B(_06499_),
    .A(\soc_I.spi0_I.div[3] ),
    .X(_06536_));
 sg13g2_xnor2_1 _28742_ (.Y(_06537_),
    .A(\soc_I.spi0_I.tick_cnt[3] ),
    .B(_06536_));
 sg13g2_xor2_1 _28743_ (.B(_06500_),
    .A(\soc_I.spi0_I.div[4] ),
    .X(_06538_));
 sg13g2_xnor2_1 _28744_ (.Y(_06539_),
    .A(\soc_I.spi0_I.tick_cnt[4] ),
    .B(_06538_));
 sg13g2_nand4_1 _28745_ (.B(_06535_),
    .C(_06537_),
    .A(_06532_),
    .Y(_06540_),
    .D(_06539_));
 sg13g2_xnor2_1 _28746_ (.Y(_06541_),
    .A(\soc_I.spi0_I.div[6] ),
    .B(_06502_));
 sg13g2_xnor2_1 _28747_ (.Y(_06542_),
    .A(\soc_I.spi0_I.tick_cnt[6] ),
    .B(_06541_));
 sg13g2_nor4_1 _28748_ (.A(_06525_),
    .B(_06527_),
    .C(_06540_),
    .D(_06542_),
    .Y(_06543_));
 sg13g2_o21ai_1 _28749_ (.B1(_06543_),
    .Y(_06544_),
    .A1(\soc_I.spi0_I.tick_cnt[10] ),
    .A2(_06523_));
 sg13g2_a21oi_1 _28750_ (.A1(\soc_I.spi0_I.tick_cnt[10] ),
    .A2(_06523_),
    .Y(_06545_),
    .B1(_06544_));
 sg13g2_xnor2_1 _28751_ (.Y(_06546_),
    .A(\soc_I.spi0_I.tick_cnt[14] ),
    .B(_06511_));
 sg13g2_xnor2_1 _28752_ (.Y(_06547_),
    .A(\soc_I.spi0_I.tick_cnt[12] ),
    .B(_06514_));
 sg13g2_a21oi_1 _28753_ (.A1(\soc_I.spi0_I.tick_cnt[13] ),
    .A2(_06513_),
    .Y(_06548_),
    .B1(_06547_));
 sg13g2_o21ai_1 _28754_ (.B1(_06548_),
    .Y(_06549_),
    .A1(\soc_I.spi0_I.tick_cnt[15] ),
    .A2(_06518_));
 sg13g2_xnor2_1 _28755_ (.Y(_06550_),
    .A(_06521_),
    .B(_06522_));
 sg13g2_xnor2_1 _28756_ (.Y(_06551_),
    .A(_00287_),
    .B(_06504_));
 sg13g2_and2_1 _28757_ (.A(\soc_I.spi0_I.tick_cnt[8] ),
    .B(_06551_),
    .X(_06552_));
 sg13g2_o21ai_1 _28758_ (.B1(_06517_),
    .Y(_06553_),
    .A1(\soc_I.spi0_I.tick_cnt[8] ),
    .A2(_06551_));
 sg13g2_nor4_1 _28759_ (.A(_06516_),
    .B(_06550_),
    .C(_06552_),
    .D(_06553_),
    .Y(_06554_));
 sg13g2_nand3_1 _28760_ (.B(_06545_),
    .C(_06554_),
    .A(_06520_),
    .Y(_06555_));
 sg13g2_nor4_2 _28761_ (.A(_06510_),
    .B(_06546_),
    .C(_06549_),
    .Y(_06556_),
    .D(_06555_));
 sg13g2_o21ai_1 _28762_ (.B1(net8828),
    .Y(_06557_),
    .A1(_06510_),
    .A2(_06556_));
 sg13g2_nand2_1 _28763_ (.Y(_06558_),
    .A(_06497_),
    .B(_06557_));
 sg13g2_nand2_2 _28764_ (.Y(_06559_),
    .A(net7493),
    .B(_13266_));
 sg13g2_or3_1 _28765_ (.A(net3856),
    .B(net8830),
    .C(_06559_),
    .X(_06560_));
 sg13g2_nand2_1 _28766_ (.Y(_06561_),
    .A(_06558_),
    .B(_06560_));
 sg13g2_nor2_1 _28767_ (.A(\soc_I.spi0_I.sclk ),
    .B(_06557_),
    .Y(_06562_));
 sg13g2_nor2_2 _28768_ (.A(_06498_),
    .B(_06562_),
    .Y(_06563_));
 sg13g2_inv_1 _28769_ (.Y(_06564_),
    .A(_06563_));
 sg13g2_a22oi_1 _28770_ (.Y(_06565_),
    .B1(_06564_),
    .B2(_06560_),
    .A2(_06561_),
    .A1(net4307));
 sg13g2_nand2_1 _28771_ (.Y(_01745_),
    .A(net9325),
    .B(net4308));
 sg13g2_nand2_2 _28772_ (.Y(_06566_),
    .A(net9323),
    .B(_06497_));
 sg13g2_xor2_1 _28773_ (.B(_06563_),
    .A(net5044),
    .X(_06567_));
 sg13g2_nor2_1 _28774_ (.A(_06566_),
    .B(_06567_),
    .Y(_01746_));
 sg13g2_nor3_1 _28775_ (.A(net5041),
    .B(\soc_I.spi0_I.xfer_cycles[0] ),
    .C(_06563_),
    .Y(_06568_));
 sg13g2_o21ai_1 _28776_ (.B1(net5041),
    .Y(_06569_),
    .A1(\soc_I.spi0_I.xfer_cycles[0] ),
    .A2(_06563_));
 sg13g2_nor2b_1 _28777_ (.A(net5042),
    .B_N(_06569_),
    .Y(_06570_));
 sg13g2_nor2_1 _28778_ (.A(_06566_),
    .B(net5043),
    .Y(_01747_));
 sg13g2_xnor2_1 _28779_ (.Y(_06571_),
    .A(net4675),
    .B(_06568_));
 sg13g2_nor2_1 _28780_ (.A(_06566_),
    .B(net4676),
    .Y(_01748_));
 sg13g2_nor4_1 _28781_ (.A(\soc_I.spi0_I.xfer_cycles[2] ),
    .B(\soc_I.spi0_I.xfer_cycles[1] ),
    .C(\soc_I.spi0_I.xfer_cycles[0] ),
    .D(_06563_),
    .Y(_06572_));
 sg13g2_o21ai_1 _28782_ (.B1(net9324),
    .Y(_06573_),
    .A1(net3190),
    .A2(_06572_));
 sg13g2_nand3_1 _28783_ (.B(_13154_),
    .C(_14437_),
    .A(net7491),
    .Y(_06574_));
 sg13g2_o21ai_1 _28784_ (.B1(_06498_),
    .Y(_06575_),
    .A1(_14438_),
    .A2(_06559_));
 sg13g2_a221oi_1 _28785_ (.B2(_06498_),
    .C1(_06573_),
    .B1(_06574_),
    .A1(net3190),
    .Y(_01749_),
    .A2(_06572_));
 sg13g2_nand2_1 _28786_ (.Y(_06576_),
    .A(net4292),
    .B(_06563_));
 sg13g2_xnor2_1 _28787_ (.Y(_06577_),
    .A(_10693_),
    .B(_13794_));
 sg13g2_nand2_1 _28788_ (.Y(_06578_),
    .A(_06562_),
    .B(_06577_));
 sg13g2_a21oi_1 _28789_ (.A1(_06576_),
    .A2(_06578_),
    .Y(_01750_),
    .B1(net9014));
 sg13g2_nor3_1 _28790_ (.A(_10693_),
    .B(_13794_),
    .C(_06563_),
    .Y(_06579_));
 sg13g2_xnor2_1 _28791_ (.Y(_06580_),
    .A(net4738),
    .B(_06579_));
 sg13g2_nor2_1 _28792_ (.A(_06566_),
    .B(net4739),
    .Y(_01751_));
 sg13g2_o21ai_1 _28793_ (.B1(net4537),
    .Y(_06581_),
    .A1(net3856),
    .A2(net8830));
 sg13g2_a21oi_1 _28794_ (.A1(_06560_),
    .A2(_06581_),
    .Y(_01752_),
    .B1(net9014));
 sg13g2_o21ai_1 _28795_ (.B1(net9334),
    .Y(_06582_),
    .A1(\soc_I.spi0_I.spi_buf[7] ),
    .A2(_06557_));
 sg13g2_a21oi_1 _28796_ (.A1(_10398_),
    .A2(_06557_),
    .Y(_01753_),
    .B1(_06582_));
 sg13g2_nand2_1 _28797_ (.Y(_06583_),
    .A(net3856),
    .B(net8830));
 sg13g2_a21oi_1 _28798_ (.A1(_06560_),
    .A2(_06583_),
    .Y(_01754_),
    .B1(net9014));
 sg13g2_a21oi_2 _28799_ (.B1(_06563_),
    .Y(_06584_),
    .A2(_06574_),
    .A1(_06498_));
 sg13g2_and2_2 _28800_ (.A(_06564_),
    .B(_06575_),
    .X(_06585_));
 sg13g2_o21ai_1 _28801_ (.B1(net9325),
    .Y(_06586_),
    .A1(net4828),
    .A2(_06585_));
 sg13g2_nor2_1 _28802_ (.A(net8831),
    .B(_13978_),
    .Y(_06587_));
 sg13g2_a21oi_1 _28803_ (.A1(net4),
    .A2(net8830),
    .Y(_06588_),
    .B1(_06587_));
 sg13g2_a21oi_1 _28804_ (.A1(_06584_),
    .A2(_06588_),
    .Y(_01755_),
    .B1(_06586_));
 sg13g2_o21ai_1 _28805_ (.B1(net9326),
    .Y(_06589_),
    .A1(net3719),
    .A2(_06585_));
 sg13g2_nor2_1 _28806_ (.A(net8831),
    .B(net8612),
    .Y(_06590_));
 sg13g2_a21oi_1 _28807_ (.A1(net4828),
    .A2(net8830),
    .Y(_06591_),
    .B1(_06590_));
 sg13g2_a21oi_1 _28808_ (.A1(_06584_),
    .A2(_06591_),
    .Y(_01756_),
    .B1(_06589_));
 sg13g2_o21ai_1 _28809_ (.B1(net9325),
    .Y(_06592_),
    .A1(net3947),
    .A2(_06585_));
 sg13g2_nor2_1 _28810_ (.A(net8830),
    .B(net8610),
    .Y(_06593_));
 sg13g2_a21oi_1 _28811_ (.A1(net3719),
    .A2(net8830),
    .Y(_06594_),
    .B1(_06593_));
 sg13g2_a21oi_1 _28812_ (.A1(_06584_),
    .A2(_06594_),
    .Y(_01757_),
    .B1(_06592_));
 sg13g2_o21ai_1 _28813_ (.B1(net9324),
    .Y(_06595_),
    .A1(net4316),
    .A2(_06585_));
 sg13g2_nor2_1 _28814_ (.A(net8829),
    .B(net8549),
    .Y(_06596_));
 sg13g2_a21oi_1 _28815_ (.A1(net3947),
    .A2(net8828),
    .Y(_06597_),
    .B1(_06596_));
 sg13g2_a21oi_1 _28816_ (.A1(_06584_),
    .A2(_06597_),
    .Y(_01758_),
    .B1(_06595_));
 sg13g2_o21ai_1 _28817_ (.B1(net9324),
    .Y(_06598_),
    .A1(net4008),
    .A2(_06585_));
 sg13g2_nor2_1 _28818_ (.A(net8829),
    .B(net8608),
    .Y(_06599_));
 sg13g2_a21oi_1 _28819_ (.A1(net4316),
    .A2(net8828),
    .Y(_06600_),
    .B1(_06599_));
 sg13g2_a21oi_1 _28820_ (.A1(_06584_),
    .A2(_06600_),
    .Y(_01759_),
    .B1(_06598_));
 sg13g2_o21ai_1 _28821_ (.B1(net9324),
    .Y(_06601_),
    .A1(net4102),
    .A2(_06585_));
 sg13g2_nor2_1 _28822_ (.A(net8829),
    .B(net8606),
    .Y(_06602_));
 sg13g2_a21oi_1 _28823_ (.A1(net4008),
    .A2(net8828),
    .Y(_06603_),
    .B1(_06602_));
 sg13g2_a21oi_1 _28824_ (.A1(_06584_),
    .A2(_06603_),
    .Y(_01760_),
    .B1(_06601_));
 sg13g2_o21ai_1 _28825_ (.B1(net9326),
    .Y(_06604_),
    .A1(net4645),
    .A2(_06585_));
 sg13g2_nor2_1 _28826_ (.A(net8829),
    .B(net8604),
    .Y(_06605_));
 sg13g2_a21oi_1 _28827_ (.A1(net4102),
    .A2(net8829),
    .Y(_06606_),
    .B1(_06605_));
 sg13g2_a21oi_1 _28828_ (.A1(_06584_),
    .A2(_06606_),
    .Y(_01761_),
    .B1(_06604_));
 sg13g2_o21ai_1 _28829_ (.B1(net9334),
    .Y(_06607_),
    .A1(net3705),
    .A2(_06585_));
 sg13g2_nor2_1 _28830_ (.A(_10379_),
    .B(_13795_),
    .Y(_06608_));
 sg13g2_a21oi_1 _28831_ (.A1(_13795_),
    .A2(_14025_),
    .Y(_06609_),
    .B1(_06608_));
 sg13g2_a21oi_1 _28832_ (.A1(_06584_),
    .A2(_06609_),
    .Y(_01762_),
    .B1(_06607_));
 sg13g2_nor2_1 _28833_ (.A(net9297),
    .B(_06556_),
    .Y(_06610_));
 sg13g2_nand2_1 _28834_ (.Y(_06611_),
    .A(net8828),
    .B(_06610_));
 sg13g2_and3_1 _28835_ (.X(_01763_),
    .A(net2598),
    .B(net8828),
    .C(_06610_));
 sg13g2_xnor2_1 _28836_ (.Y(_06612_),
    .A(\soc_I.spi0_I.tick_cnt[1] ),
    .B(net4988));
 sg13g2_nor2_1 _28837_ (.A(net7682),
    .B(net4989),
    .Y(_01764_));
 sg13g2_and3_1 _28838_ (.X(_06613_),
    .A(net3819),
    .B(\soc_I.spi0_I.tick_cnt[1] ),
    .C(\soc_I.spi0_I.tick_cnt[0] ));
 sg13g2_a21oi_1 _28839_ (.A1(\soc_I.spi0_I.tick_cnt[1] ),
    .A2(\soc_I.spi0_I.tick_cnt[0] ),
    .Y(_06614_),
    .B1(net3819));
 sg13g2_nor3_1 _28840_ (.A(net7682),
    .B(_06613_),
    .C(net3820),
    .Y(_01765_));
 sg13g2_and3_1 _28841_ (.X(_06615_),
    .A(net3871),
    .B(net8828),
    .C(_06613_));
 sg13g2_a21oi_1 _28842_ (.A1(net8828),
    .A2(_06613_),
    .Y(_06616_),
    .B1(net3871));
 sg13g2_nor3_1 _28843_ (.A(net7682),
    .B(_06615_),
    .C(net3872),
    .Y(_01766_));
 sg13g2_and2_1 _28844_ (.A(net4413),
    .B(_06615_),
    .X(_06617_));
 sg13g2_nor2_1 _28845_ (.A(net4413),
    .B(_06615_),
    .Y(_06618_));
 sg13g2_nor3_1 _28846_ (.A(net7682),
    .B(_06617_),
    .C(_06618_),
    .Y(_01767_));
 sg13g2_xnor2_1 _28847_ (.Y(_06619_),
    .A(net5012),
    .B(_06617_));
 sg13g2_nor2_1 _28848_ (.A(_06611_),
    .B(_06619_),
    .Y(_01768_));
 sg13g2_and3_1 _28849_ (.X(_06620_),
    .A(net3425),
    .B(\soc_I.spi0_I.tick_cnt[5] ),
    .C(_06617_));
 sg13g2_a21oi_1 _28850_ (.A1(\soc_I.spi0_I.tick_cnt[5] ),
    .A2(_06617_),
    .Y(_06621_),
    .B1(net3425));
 sg13g2_nor3_1 _28851_ (.A(_06611_),
    .B(_06620_),
    .C(net3426),
    .Y(_01769_));
 sg13g2_and2_1 _28852_ (.A(net4279),
    .B(_06620_),
    .X(_06622_));
 sg13g2_nor2_1 _28853_ (.A(net4279),
    .B(_06620_),
    .Y(_06623_));
 sg13g2_nor3_1 _28854_ (.A(net7681),
    .B(_06622_),
    .C(net4280),
    .Y(_01770_));
 sg13g2_and2_1 _28855_ (.A(net4571),
    .B(_06622_),
    .X(_06624_));
 sg13g2_nor2_1 _28856_ (.A(net4571),
    .B(_06622_),
    .Y(_06625_));
 sg13g2_nor3_1 _28857_ (.A(net7681),
    .B(_06624_),
    .C(_06625_),
    .Y(_01771_));
 sg13g2_and2_1 _28858_ (.A(net4287),
    .B(_06624_),
    .X(_06626_));
 sg13g2_nor2_1 _28859_ (.A(net4287),
    .B(_06624_),
    .Y(_06627_));
 sg13g2_nor3_1 _28860_ (.A(net7681),
    .B(_06626_),
    .C(net4288),
    .Y(_01772_));
 sg13g2_and2_1 _28861_ (.A(net4189),
    .B(_06626_),
    .X(_06628_));
 sg13g2_nor2_1 _28862_ (.A(net4189),
    .B(_06626_),
    .Y(_06629_));
 sg13g2_nor3_1 _28863_ (.A(net7681),
    .B(_06628_),
    .C(net4190),
    .Y(_01773_));
 sg13g2_and2_1 _28864_ (.A(net4434),
    .B(_06628_),
    .X(_06630_));
 sg13g2_nor2_1 _28865_ (.A(net4434),
    .B(_06628_),
    .Y(_06631_));
 sg13g2_nor3_1 _28866_ (.A(net7681),
    .B(_06630_),
    .C(_06631_),
    .Y(_01774_));
 sg13g2_and2_1 _28867_ (.A(net4467),
    .B(_06630_),
    .X(_06632_));
 sg13g2_nor2_1 _28868_ (.A(net4467),
    .B(_06630_),
    .Y(_06633_));
 sg13g2_nor3_1 _28869_ (.A(net7681),
    .B(_06632_),
    .C(_06633_),
    .Y(_01775_));
 sg13g2_and2_1 _28870_ (.A(net4346),
    .B(_06632_),
    .X(_06634_));
 sg13g2_nor2_1 _28871_ (.A(net4346),
    .B(_06632_),
    .Y(_06635_));
 sg13g2_nor3_1 _28872_ (.A(net7681),
    .B(_06634_),
    .C(net4347),
    .Y(_01776_));
 sg13g2_and2_1 _28873_ (.A(net4251),
    .B(_06634_),
    .X(_06636_));
 sg13g2_nor2_1 _28874_ (.A(net4251),
    .B(_06634_),
    .Y(_06637_));
 sg13g2_nor3_1 _28875_ (.A(net7681),
    .B(_06636_),
    .C(net4252),
    .Y(_01777_));
 sg13g2_and2_1 _28876_ (.A(net4656),
    .B(_06636_),
    .X(_06638_));
 sg13g2_nor2_1 _28877_ (.A(net4656),
    .B(_06636_),
    .Y(_06639_));
 sg13g2_nor3_1 _28878_ (.A(net7682),
    .B(_06638_),
    .C(_06639_),
    .Y(_01778_));
 sg13g2_nand2_1 _28879_ (.Y(_06640_),
    .A(\soc_I.spi0_I.tick_cnt[16] ),
    .B(_06638_));
 sg13g2_xnor2_1 _28880_ (.Y(_06641_),
    .A(net4508),
    .B(_06638_));
 sg13g2_nor2_1 _28881_ (.A(net7682),
    .B(net4509),
    .Y(_01779_));
 sg13g2_xor2_1 _28882_ (.B(_06640_),
    .A(net4487),
    .X(_06642_));
 sg13g2_nor2_1 _28883_ (.A(net7682),
    .B(net4488),
    .Y(_01780_));
 sg13g2_nand3_1 _28884_ (.B(_13154_),
    .C(_14437_),
    .A(_12895_),
    .Y(_06643_));
 sg13g2_a21oi_1 _28885_ (.A1(net4561),
    .A2(_06643_),
    .Y(_06644_),
    .B1(net9020));
 sg13g2_o21ai_1 _28886_ (.B1(_06644_),
    .Y(_01781_),
    .A1(_13977_),
    .A2(_06643_));
 sg13g2_nor2_2 _28887_ (.A(_00292_),
    .B(_13237_),
    .Y(_06645_));
 sg13g2_or2_2 _28888_ (.X(_06646_),
    .B(_13237_),
    .A(_00292_));
 sg13g2_nand2b_1 _28889_ (.Y(_06647_),
    .B(net8819),
    .A_N(net4164));
 sg13g2_a21oi_1 _28890_ (.A1(net4164),
    .A2(_14121_),
    .Y(_06648_),
    .B1(_06646_));
 sg13g2_o21ai_1 _28891_ (.B1(_06647_),
    .Y(_06649_),
    .A1(\soc_I.rx_uart_i.fifo_i.cnt[0] ),
    .A2(net8819));
 sg13g2_a221oi_1 _28892_ (.B2(_06646_),
    .C1(net9002),
    .B1(_06649_),
    .A1(_06647_),
    .Y(_01782_),
    .A2(_06648_));
 sg13g2_a21oi_1 _28893_ (.A1(\soc_I.rx_uart_i.ready ),
    .A2(\soc_I.rx_uart_i.fifo_i.cnt[0] ),
    .Y(_06650_),
    .B1(net5203));
 sg13g2_nand3_1 _28894_ (.B(\soc_I.rx_uart_i.fifo_i.cnt[1] ),
    .C(\soc_I.rx_uart_i.fifo_i.cnt[0] ),
    .A(\soc_I.rx_uart_i.ready ),
    .Y(_06651_));
 sg13g2_nand2b_1 _28895_ (.Y(_06652_),
    .B(_06651_),
    .A_N(_06650_));
 sg13g2_o21ai_1 _28896_ (.B1(net5203),
    .Y(_06653_),
    .A1(\soc_I.rx_uart_i.ready ),
    .A2(\soc_I.rx_uart_i.fifo_i.cnt[0] ));
 sg13g2_nor3_1 _28897_ (.A(net5203),
    .B(\soc_I.rx_uart_i.fifo_i.cnt[0] ),
    .C(net8819),
    .Y(_06654_));
 sg13g2_nor2_1 _28898_ (.A(_06646_),
    .B(_06654_),
    .Y(_06655_));
 sg13g2_a221oi_1 _28899_ (.B2(_06655_),
    .C1(net9002),
    .B1(net5204),
    .A1(_06646_),
    .Y(_01783_),
    .A2(_06652_));
 sg13g2_a21oi_1 _28900_ (.A1(_06646_),
    .A2(_06651_),
    .Y(_06656_),
    .B1(_06655_));
 sg13g2_o21ai_1 _28901_ (.B1(net9298),
    .Y(_06657_),
    .A1(net4249),
    .A2(_06656_));
 sg13g2_a21oi_1 _28902_ (.A1(net4249),
    .A2(_06656_),
    .Y(_01784_),
    .B1(_06657_));
 sg13g2_nor3_1 _28903_ (.A(_10650_),
    .B(_06645_),
    .C(_06651_),
    .Y(_06658_));
 sg13g2_nor3_1 _28904_ (.A(\soc_I.rx_uart_i.fifo_i.cnt[0] ),
    .B(net8819),
    .C(_06646_),
    .Y(_06659_));
 sg13g2_a21o_1 _28905_ (.A2(_06659_),
    .A1(_13235_),
    .B1(_06658_),
    .X(_06660_));
 sg13g2_o21ai_1 _28906_ (.B1(net9298),
    .Y(_06661_),
    .A1(net3837),
    .A2(_06660_));
 sg13g2_a21oi_1 _28907_ (.A1(net3837),
    .A2(_06660_),
    .Y(_01785_),
    .B1(_06661_));
 sg13g2_nand2_1 _28908_ (.Y(_06662_),
    .A(net3837),
    .B(_06658_));
 sg13g2_o21ai_1 _28909_ (.B1(net9298),
    .Y(_06663_),
    .A1(net4012),
    .A2(_14119_));
 sg13g2_xor2_1 _28910_ (.B(_06662_),
    .A(net5106),
    .X(_06664_));
 sg13g2_nor2_1 _28911_ (.A(_06663_),
    .B(_06664_),
    .Y(_01786_));
 sg13g2_nor2_1 _28912_ (.A(_13182_),
    .B(_14437_),
    .Y(_06665_));
 sg13g2_nand3_1 _28913_ (.B(_13263_),
    .C(_14438_),
    .A(_13173_),
    .Y(_06666_));
 sg13g2_nor2_1 _28914_ (.A(net4216),
    .B(net7364),
    .Y(_06667_));
 sg13g2_nand2_1 _28915_ (.Y(_06668_),
    .A(\gpio_uo_en[0] ),
    .B(_13177_));
 sg13g2_a22oi_1 _28916_ (.Y(_06669_),
    .B1(_13180_),
    .B2(net2),
    .A2(_13176_),
    .A1(\gpio_uo_out[0] ));
 sg13g2_and3_1 _28917_ (.X(_06670_),
    .A(net7364),
    .B(_06668_),
    .C(_06669_));
 sg13g2_nor3_1 _28918_ (.A(net9013),
    .B(_06667_),
    .C(_06670_),
    .Y(_01787_));
 sg13g2_o21ai_1 _28919_ (.B1(net9334),
    .Y(_06671_),
    .A1(\soc_I.gpio0_I.rdata[1] ),
    .A2(net7363));
 sg13g2_nand2_1 _28920_ (.Y(_06672_),
    .A(net3405),
    .B(_13260_));
 sg13g2_a221oi_1 _28921_ (.B2(net3),
    .C1(_06666_),
    .B1(_13262_),
    .A1(\gpio_uo_en[1] ),
    .Y(_06673_),
    .A2(_13261_));
 sg13g2_a21oi_1 _28922_ (.A1(_06672_),
    .A2(_06673_),
    .Y(_01788_),
    .B1(_06671_));
 sg13g2_nor2_1 _28923_ (.A(net4640),
    .B(net7363),
    .Y(_06674_));
 sg13g2_nand2_1 _28924_ (.Y(_06675_),
    .A(\gpio_uo_out[2] ),
    .B(_13176_));
 sg13g2_a22oi_1 _28925_ (.Y(_06676_),
    .B1(_13180_),
    .B2(net4),
    .A2(_13177_),
    .A1(\gpio_uo_en[2] ));
 sg13g2_and3_1 _28926_ (.X(_06677_),
    .A(net7363),
    .B(_06675_),
    .C(_06676_));
 sg13g2_nor3_1 _28927_ (.A(net9014),
    .B(_06674_),
    .C(_06677_),
    .Y(_01789_));
 sg13g2_nor2_1 _28928_ (.A(net4634),
    .B(net7364),
    .Y(_06678_));
 sg13g2_nand2_1 _28929_ (.Y(_06679_),
    .A(\gpio_uo_out[3] ),
    .B(_13176_));
 sg13g2_a22oi_1 _28930_ (.Y(_06680_),
    .B1(_13180_),
    .B2(net5),
    .A2(_13177_),
    .A1(\gpio_uo_en[3] ));
 sg13g2_and3_1 _28931_ (.X(_06681_),
    .A(net7364),
    .B(_06679_),
    .C(_06680_));
 sg13g2_nor3_1 _28932_ (.A(net9013),
    .B(_06678_),
    .C(_06681_),
    .Y(_01790_));
 sg13g2_o21ai_1 _28933_ (.B1(net9334),
    .Y(_06682_),
    .A1(\soc_I.gpio0_I.rdata[4] ),
    .A2(net7363));
 sg13g2_nand2_1 _28934_ (.Y(_06683_),
    .A(net3918),
    .B(_13260_));
 sg13g2_a221oi_1 _28935_ (.B2(net6),
    .C1(_06666_),
    .B1(_13262_),
    .A1(\gpio_uo_en[4] ),
    .Y(_06684_),
    .A2(_13261_));
 sg13g2_a21oi_1 _28936_ (.A1(_06683_),
    .A2(_06684_),
    .Y(_01791_),
    .B1(_06682_));
 sg13g2_o21ai_1 _28937_ (.B1(net9334),
    .Y(_06685_),
    .A1(\soc_I.gpio0_I.rdata[5] ),
    .A2(net7363));
 sg13g2_nand2_1 _28938_ (.Y(_06686_),
    .A(net3802),
    .B(_13260_));
 sg13g2_a221oi_1 _28939_ (.B2(net7),
    .C1(_06666_),
    .B1(_13262_),
    .A1(\gpio_uo_en[5] ),
    .Y(_06687_),
    .A2(_13261_));
 sg13g2_a21oi_1 _28940_ (.A1(_06686_),
    .A2(_06687_),
    .Y(_01792_),
    .B1(_06685_));
 sg13g2_nor2_1 _28941_ (.A(net4277),
    .B(net7363),
    .Y(_06688_));
 sg13g2_nand2_1 _28942_ (.Y(_06689_),
    .A(\gpio_uo_out[6] ),
    .B(_13176_));
 sg13g2_a22oi_1 _28943_ (.Y(_06690_),
    .B1(_13180_),
    .B2(net8),
    .A2(_13177_),
    .A1(\gpio_uo_en[6] ));
 sg13g2_and3_1 _28944_ (.X(_06691_),
    .A(net7363),
    .B(_06689_),
    .C(_06690_));
 sg13g2_nor3_1 _28945_ (.A(net9013),
    .B(_06688_),
    .C(_06691_),
    .Y(_01793_));
 sg13g2_o21ai_1 _28946_ (.B1(net9334),
    .Y(_06692_),
    .A1(\soc_I.gpio0_I.rdata[7] ),
    .A2(net7363));
 sg13g2_nand2_1 _28947_ (.Y(_06693_),
    .A(net4061),
    .B(_13260_));
 sg13g2_a221oi_1 _28948_ (.B2(net9),
    .C1(_06666_),
    .B1(_13262_),
    .A1(\gpio_uo_en[7] ),
    .Y(_06694_),
    .A2(_13261_));
 sg13g2_a21oi_1 _28949_ (.A1(_06693_),
    .A2(_06694_),
    .Y(_01794_),
    .B1(_06692_));
 sg13g2_nor2_2 _28950_ (.A(\soc_I.rx_uart_i.state[1] ),
    .B(\soc_I.rx_uart_i.state[0] ),
    .Y(_06695_));
 sg13g2_and2_1 _28951_ (.A(\soc_I.rx_uart_i.state[2] ),
    .B(_06695_),
    .X(_06696_));
 sg13g2_nand2_2 _28952_ (.Y(_06697_),
    .A(net3400),
    .B(_06695_));
 sg13g2_nor2_1 _28953_ (.A(\soc_I.rx_uart_i.wait_states[7] ),
    .B(\soc_I.rx_uart_i.wait_states[6] ),
    .Y(_06698_));
 sg13g2_nor2_1 _28954_ (.A(\soc_I.rx_uart_i.wait_states[3] ),
    .B(\soc_I.rx_uart_i.wait_states[2] ),
    .Y(_06699_));
 sg13g2_nor4_2 _28955_ (.A(\soc_I.rx_uart_i.wait_states[15] ),
    .B(\soc_I.rx_uart_i.wait_states[14] ),
    .C(\soc_I.rx_uart_i.wait_states[13] ),
    .Y(_06700_),
    .D(\soc_I.rx_uart_i.wait_states[12] ));
 sg13g2_nor2_1 _28956_ (.A(\soc_I.rx_uart_i.wait_states[11] ),
    .B(\soc_I.rx_uart_i.wait_states[10] ),
    .Y(_06701_));
 sg13g2_nor3_1 _28957_ (.A(\soc_I.rx_uart_i.wait_states[8] ),
    .B(\soc_I.rx_uart_i.wait_states[7] ),
    .C(\soc_I.rx_uart_i.wait_states[6] ),
    .Y(_06702_));
 sg13g2_nor3_1 _28958_ (.A(\soc_I.rx_uart_i.wait_states[11] ),
    .B(\soc_I.rx_uart_i.wait_states[10] ),
    .C(\soc_I.rx_uart_i.wait_states[9] ),
    .Y(_06703_));
 sg13g2_nand3_1 _28959_ (.B(_00290_),
    .C(_06699_),
    .A(\soc_I.rx_uart_i.wait_states[0] ),
    .Y(_06704_));
 sg13g2_nor4_1 _28960_ (.A(\soc_I.rx_uart_i.wait_states[5] ),
    .B(\soc_I.rx_uart_i.wait_states[4] ),
    .C(\soc_I.rx_uart_i.wait_states[1] ),
    .D(_06704_),
    .Y(_06705_));
 sg13g2_nand4_1 _28961_ (.B(_06702_),
    .C(_06703_),
    .A(_06700_),
    .Y(_06706_),
    .D(_06705_));
 sg13g2_nand2_1 _28962_ (.Y(_06707_),
    .A(net8800),
    .B(_06706_));
 sg13g2_nor2_1 _28963_ (.A(net3009),
    .B(net2611),
    .Y(_06708_));
 sg13g2_nand3_1 _28964_ (.B(_06707_),
    .C(_06708_),
    .A(_06695_),
    .Y(_06709_));
 sg13g2_a221oi_1 _28965_ (.B2(_10397_),
    .C1(net9003),
    .B1(_06709_),
    .A1(_10395_),
    .Y(_01795_),
    .A2(_06695_));
 sg13g2_nand2_1 _28966_ (.Y(_06710_),
    .A(net2859),
    .B(net8553));
 sg13g2_nor2_1 _28967_ (.A(\soc_I.qqspi_I.spi_buf[24] ),
    .B(net7464),
    .Y(_06711_));
 sg13g2_o21ai_1 _28968_ (.B1(net8557),
    .Y(_06712_),
    .A1(\soc_I.qqspi_I.spi_buf[0] ),
    .A2(net7454));
 sg13g2_o21ai_1 _28969_ (.B1(_06710_),
    .Y(_01796_),
    .A1(_06711_),
    .A2(_06712_));
 sg13g2_nand2_1 _28970_ (.Y(_06713_),
    .A(net2849),
    .B(net8552));
 sg13g2_nor2_1 _28971_ (.A(\soc_I.qqspi_I.spi_buf[25] ),
    .B(net7460),
    .Y(_06714_));
 sg13g2_o21ai_1 _28972_ (.B1(net8557),
    .Y(_06715_),
    .A1(\soc_I.qqspi_I.spi_buf[1] ),
    .A2(net7455));
 sg13g2_o21ai_1 _28973_ (.B1(_06713_),
    .Y(_01797_),
    .A1(_06714_),
    .A2(_06715_));
 sg13g2_nand2_1 _28974_ (.Y(_06716_),
    .A(net2677),
    .B(net8551));
 sg13g2_nor2_1 _28975_ (.A(\soc_I.qqspi_I.spi_buf[26] ),
    .B(net7461),
    .Y(_06717_));
 sg13g2_o21ai_1 _28976_ (.B1(net8558),
    .Y(_06718_),
    .A1(\soc_I.qqspi_I.spi_buf[2] ),
    .A2(net7454));
 sg13g2_o21ai_1 _28977_ (.B1(_06716_),
    .Y(_01798_),
    .A1(_06717_),
    .A2(_06718_));
 sg13g2_nand2_1 _28978_ (.Y(_06719_),
    .A(net3444),
    .B(net8552));
 sg13g2_nor2_1 _28979_ (.A(\soc_I.qqspi_I.spi_buf[27] ),
    .B(net7460),
    .Y(_06720_));
 sg13g2_o21ai_1 _28980_ (.B1(net8556),
    .Y(_06721_),
    .A1(\soc_I.qqspi_I.spi_buf[3] ),
    .A2(net7454));
 sg13g2_o21ai_1 _28981_ (.B1(_06719_),
    .Y(_01799_),
    .A1(_06720_),
    .A2(_06721_));
 sg13g2_nand2_1 _28982_ (.Y(_06722_),
    .A(net2813),
    .B(net8552));
 sg13g2_nor2_1 _28983_ (.A(\soc_I.qqspi_I.spi_buf[28] ),
    .B(net7459),
    .Y(_06723_));
 sg13g2_o21ai_1 _28984_ (.B1(net8556),
    .Y(_06724_),
    .A1(\soc_I.qqspi_I.spi_buf[4] ),
    .A2(net7455));
 sg13g2_o21ai_1 _28985_ (.B1(_06722_),
    .Y(_01800_),
    .A1(_06723_),
    .A2(_06724_));
 sg13g2_nand2_1 _28986_ (.Y(_06725_),
    .A(net2783),
    .B(net8551));
 sg13g2_nor2_1 _28987_ (.A(\soc_I.qqspi_I.spi_buf[29] ),
    .B(net7459),
    .Y(_06726_));
 sg13g2_o21ai_1 _28988_ (.B1(net8556),
    .Y(_06727_),
    .A1(\soc_I.qqspi_I.spi_buf[5] ),
    .A2(net7454));
 sg13g2_o21ai_1 _28989_ (.B1(_06725_),
    .Y(_01801_),
    .A1(_06726_),
    .A2(_06727_));
 sg13g2_nand2_1 _28990_ (.Y(_06728_),
    .A(net2697),
    .B(net8551));
 sg13g2_nor2_1 _28991_ (.A(\soc_I.qqspi_I.spi_buf[30] ),
    .B(net7459),
    .Y(_06729_));
 sg13g2_o21ai_1 _28992_ (.B1(net8556),
    .Y(_06730_),
    .A1(\soc_I.qqspi_I.spi_buf[6] ),
    .A2(net7454));
 sg13g2_o21ai_1 _28993_ (.B1(_06728_),
    .Y(_01802_),
    .A1(_06729_),
    .A2(_06730_));
 sg13g2_nand2_1 _28994_ (.Y(_06731_),
    .A(net2949),
    .B(net8552));
 sg13g2_nor2_1 _28995_ (.A(\soc_I.qqspi_I.spi_buf[31] ),
    .B(net7459),
    .Y(_06732_));
 sg13g2_o21ai_1 _28996_ (.B1(net8557),
    .Y(_06733_),
    .A1(\soc_I.qqspi_I.spi_buf[7] ),
    .A2(net7455));
 sg13g2_o21ai_1 _28997_ (.B1(_06731_),
    .Y(_01803_),
    .A1(_06732_),
    .A2(_06733_));
 sg13g2_nand2_1 _28998_ (.Y(_06734_),
    .A(net3745),
    .B(net8551));
 sg13g2_nor2_1 _28999_ (.A(\soc_I.qqspi_I.spi_buf[16] ),
    .B(net7461),
    .Y(_06735_));
 sg13g2_o21ai_1 _29000_ (.B1(net8558),
    .Y(_06736_),
    .A1(\soc_I.qqspi_I.spi_buf[8] ),
    .A2(net7456));
 sg13g2_o21ai_1 _29001_ (.B1(_06734_),
    .Y(_01804_),
    .A1(_06735_),
    .A2(_06736_));
 sg13g2_nand2_1 _29002_ (.Y(_06737_),
    .A(net3883),
    .B(net8554));
 sg13g2_nor2_1 _29003_ (.A(\soc_I.qqspi_I.spi_buf[17] ),
    .B(net7463),
    .Y(_06738_));
 sg13g2_o21ai_1 _29004_ (.B1(net8560),
    .Y(_06739_),
    .A1(\soc_I.qqspi_I.spi_buf[9] ),
    .A2(net7457));
 sg13g2_o21ai_1 _29005_ (.B1(_06737_),
    .Y(_01805_),
    .A1(_06738_),
    .A2(_06739_));
 sg13g2_nand2_1 _29006_ (.Y(_06740_),
    .A(net3976),
    .B(net8554));
 sg13g2_nor2_1 _29007_ (.A(\soc_I.qqspi_I.spi_buf[18] ),
    .B(net7463),
    .Y(_06741_));
 sg13g2_o21ai_1 _29008_ (.B1(net8560),
    .Y(_06742_),
    .A1(\soc_I.qqspi_I.spi_buf[10] ),
    .A2(net7457));
 sg13g2_o21ai_1 _29009_ (.B1(_06740_),
    .Y(_01806_),
    .A1(_06741_),
    .A2(_06742_));
 sg13g2_nand2_1 _29010_ (.Y(_06743_),
    .A(net2654),
    .B(net8553));
 sg13g2_nor2_1 _29011_ (.A(\soc_I.qqspi_I.spi_buf[19] ),
    .B(net7462),
    .Y(_06744_));
 sg13g2_o21ai_1 _29012_ (.B1(net8559),
    .Y(_06745_),
    .A1(\soc_I.qqspi_I.spi_buf[11] ),
    .A2(net7456));
 sg13g2_o21ai_1 _29013_ (.B1(_06743_),
    .Y(_01807_),
    .A1(_06744_),
    .A2(_06745_));
 sg13g2_nand2_1 _29014_ (.Y(_06746_),
    .A(net3651),
    .B(net8553));
 sg13g2_nor2_1 _29015_ (.A(\soc_I.qqspi_I.spi_buf[20] ),
    .B(net7462),
    .Y(_06747_));
 sg13g2_o21ai_1 _29016_ (.B1(net8559),
    .Y(_06748_),
    .A1(\soc_I.qqspi_I.spi_buf[12] ),
    .A2(net7456));
 sg13g2_o21ai_1 _29017_ (.B1(_06746_),
    .Y(_01808_),
    .A1(_06747_),
    .A2(_06748_));
 sg13g2_nand2_1 _29018_ (.Y(_06749_),
    .A(net3145),
    .B(net8553));
 sg13g2_nor2_1 _29019_ (.A(\soc_I.qqspi_I.spi_buf[21] ),
    .B(net7462),
    .Y(_06750_));
 sg13g2_o21ai_1 _29020_ (.B1(net8559),
    .Y(_06751_),
    .A1(\soc_I.qqspi_I.spi_buf[13] ),
    .A2(net7457));
 sg13g2_o21ai_1 _29021_ (.B1(_06749_),
    .Y(_01809_),
    .A1(_06750_),
    .A2(_06751_));
 sg13g2_nand2_1 _29022_ (.Y(_06752_),
    .A(net4166),
    .B(net8554));
 sg13g2_nor2_1 _29023_ (.A(\soc_I.qqspi_I.spi_buf[22] ),
    .B(net7463),
    .Y(_06753_));
 sg13g2_o21ai_1 _29024_ (.B1(net8559),
    .Y(_06754_),
    .A1(\soc_I.qqspi_I.spi_buf[14] ),
    .A2(net7457));
 sg13g2_o21ai_1 _29025_ (.B1(_06752_),
    .Y(_01810_),
    .A1(_06753_),
    .A2(_06754_));
 sg13g2_nand2_1 _29026_ (.Y(_06755_),
    .A(net2640),
    .B(net8554));
 sg13g2_nor2_1 _29027_ (.A(\soc_I.qqspi_I.spi_buf[23] ),
    .B(net7462),
    .Y(_06756_));
 sg13g2_o21ai_1 _29028_ (.B1(net8559),
    .Y(_06757_),
    .A1(\soc_I.qqspi_I.spi_buf[15] ),
    .A2(net7456));
 sg13g2_o21ai_1 _29029_ (.B1(_06755_),
    .Y(_01811_),
    .A1(_06756_),
    .A2(_06757_));
 sg13g2_nand2_1 _29030_ (.Y(_06758_),
    .A(net2705),
    .B(net8553));
 sg13g2_nor2_1 _29031_ (.A(\soc_I.qqspi_I.spi_buf[8] ),
    .B(net7462),
    .Y(_06759_));
 sg13g2_o21ai_1 _29032_ (.B1(net8558),
    .Y(_06760_),
    .A1(\soc_I.qqspi_I.spi_buf[16] ),
    .A2(net7456));
 sg13g2_o21ai_1 _29033_ (.B1(_06758_),
    .Y(_01812_),
    .A1(_06759_),
    .A2(_06760_));
 sg13g2_nand2_1 _29034_ (.Y(_06761_),
    .A(net3494),
    .B(net8553));
 sg13g2_nor2_1 _29035_ (.A(\soc_I.qqspi_I.spi_buf[9] ),
    .B(net7462),
    .Y(_06762_));
 sg13g2_o21ai_1 _29036_ (.B1(net8559),
    .Y(_06763_),
    .A1(\soc_I.qqspi_I.spi_buf[17] ),
    .A2(net7456));
 sg13g2_o21ai_1 _29037_ (.B1(_06761_),
    .Y(_01813_),
    .A1(_06762_),
    .A2(_06763_));
 sg13g2_nand2_1 _29038_ (.Y(_06764_),
    .A(net2781),
    .B(net8554));
 sg13g2_nor2_1 _29039_ (.A(\soc_I.qqspi_I.spi_buf[10] ),
    .B(net7464),
    .Y(_06765_));
 sg13g2_o21ai_1 _29040_ (.B1(net8560),
    .Y(_06766_),
    .A1(\soc_I.qqspi_I.spi_buf[18] ),
    .A2(net7457));
 sg13g2_o21ai_1 _29041_ (.B1(_06764_),
    .Y(_01814_),
    .A1(_06765_),
    .A2(_06766_));
 sg13g2_nand2_1 _29042_ (.Y(_06767_),
    .A(net2719),
    .B(net8555));
 sg13g2_nor2_1 _29043_ (.A(\soc_I.qqspi_I.spi_buf[11] ),
    .B(net7463),
    .Y(_06768_));
 sg13g2_o21ai_1 _29044_ (.B1(net8560),
    .Y(_06769_),
    .A1(\soc_I.qqspi_I.spi_buf[19] ),
    .A2(net7457));
 sg13g2_o21ai_1 _29045_ (.B1(_06767_),
    .Y(_01815_),
    .A1(_06768_),
    .A2(_06769_));
 sg13g2_nand2_1 _29046_ (.Y(_06770_),
    .A(net3629),
    .B(net8553));
 sg13g2_nor2_1 _29047_ (.A(\soc_I.qqspi_I.spi_buf[12] ),
    .B(net7462),
    .Y(_06771_));
 sg13g2_o21ai_1 _29048_ (.B1(net8559),
    .Y(_06772_),
    .A1(\soc_I.qqspi_I.spi_buf[20] ),
    .A2(net7456));
 sg13g2_o21ai_1 _29049_ (.B1(_06770_),
    .Y(_01816_),
    .A1(_06771_),
    .A2(_06772_));
 sg13g2_nand2_1 _29050_ (.Y(_06773_),
    .A(net2767),
    .B(net8553));
 sg13g2_nor2_1 _29051_ (.A(\soc_I.qqspi_I.spi_buf[13] ),
    .B(net7462),
    .Y(_06774_));
 sg13g2_o21ai_1 _29052_ (.B1(net8559),
    .Y(_06775_),
    .A1(\soc_I.qqspi_I.spi_buf[21] ),
    .A2(net7456));
 sg13g2_o21ai_1 _29053_ (.B1(_06773_),
    .Y(_01817_),
    .A1(_06774_),
    .A2(_06775_));
 sg13g2_nand2_1 _29054_ (.Y(_06776_),
    .A(net3085),
    .B(net8554));
 sg13g2_nor2_1 _29055_ (.A(\soc_I.qqspi_I.spi_buf[14] ),
    .B(net7463),
    .Y(_06777_));
 sg13g2_o21ai_1 _29056_ (.B1(net8560),
    .Y(_06778_),
    .A1(\soc_I.qqspi_I.spi_buf[22] ),
    .A2(net7457));
 sg13g2_o21ai_1 _29057_ (.B1(_06776_),
    .Y(_01818_),
    .A1(_06777_),
    .A2(_06778_));
 sg13g2_a21oi_1 _29058_ (.A1(_10375_),
    .A2(net7463),
    .Y(_06779_),
    .B1(net8554));
 sg13g2_o21ai_1 _29059_ (.B1(_06779_),
    .Y(_06780_),
    .A1(\soc_I.qqspi_I.spi_buf[15] ),
    .A2(net7463));
 sg13g2_o21ai_1 _29060_ (.B1(_06780_),
    .Y(_01819_),
    .A1(_10670_),
    .A2(net8560));
 sg13g2_a21oi_1 _29061_ (.A1(_10376_),
    .A2(net7464),
    .Y(_06781_),
    .B1(net8555));
 sg13g2_o21ai_1 _29062_ (.B1(_06781_),
    .Y(_06782_),
    .A1(\soc_I.qqspi_I.spi_buf[0] ),
    .A2(net7460));
 sg13g2_o21ai_1 _29063_ (.B1(_06782_),
    .Y(_01820_),
    .A1(_10656_),
    .A2(net8558));
 sg13g2_nand2_1 _29064_ (.Y(_06783_),
    .A(net2669),
    .B(net8551));
 sg13g2_nor2_1 _29065_ (.A(\soc_I.qqspi_I.spi_buf[1] ),
    .B(net7459),
    .Y(_06784_));
 sg13g2_o21ai_1 _29066_ (.B1(net8556),
    .Y(_06785_),
    .A1(\soc_I.qqspi_I.spi_buf[25] ),
    .A2(net7455));
 sg13g2_o21ai_1 _29067_ (.B1(_06783_),
    .Y(_01821_),
    .A1(_06784_),
    .A2(_06785_));
 sg13g2_nand2_1 _29068_ (.Y(_06786_),
    .A(net2779),
    .B(net8551));
 sg13g2_nor2_1 _29069_ (.A(\soc_I.qqspi_I.spi_buf[2] ),
    .B(net7461),
    .Y(_06787_));
 sg13g2_o21ai_1 _29070_ (.B1(net8558),
    .Y(_06788_),
    .A1(\soc_I.qqspi_I.spi_buf[26] ),
    .A2(net7454));
 sg13g2_o21ai_1 _29071_ (.B1(_06786_),
    .Y(_01822_),
    .A1(_06787_),
    .A2(_06788_));
 sg13g2_nand2_1 _29072_ (.Y(_06789_),
    .A(net2690),
    .B(net8552));
 sg13g2_nor2_1 _29073_ (.A(\soc_I.qqspi_I.spi_buf[3] ),
    .B(net7459),
    .Y(_06790_));
 sg13g2_o21ai_1 _29074_ (.B1(net8556),
    .Y(_06791_),
    .A1(\soc_I.qqspi_I.spi_buf[27] ),
    .A2(net7455));
 sg13g2_o21ai_1 _29075_ (.B1(_06789_),
    .Y(_01823_),
    .A1(_06790_),
    .A2(_06791_));
 sg13g2_nand2_1 _29076_ (.Y(_06792_),
    .A(net2693),
    .B(net8555));
 sg13g2_nor2_1 _29077_ (.A(\soc_I.qqspi_I.spi_buf[4] ),
    .B(net7464),
    .Y(_06793_));
 sg13g2_o21ai_1 _29078_ (.B1(net8561),
    .Y(_06794_),
    .A1(\soc_I.qqspi_I.spi_buf[28] ),
    .A2(net7458));
 sg13g2_o21ai_1 _29079_ (.B1(_06792_),
    .Y(_01824_),
    .A1(_06793_),
    .A2(_06794_));
 sg13g2_nand2_1 _29080_ (.Y(_06795_),
    .A(net2856),
    .B(net8555));
 sg13g2_nor2_1 _29081_ (.A(\soc_I.qqspi_I.spi_buf[5] ),
    .B(net7464),
    .Y(_06796_));
 sg13g2_o21ai_1 _29082_ (.B1(net8561),
    .Y(_06797_),
    .A1(\soc_I.qqspi_I.spi_buf[29] ),
    .A2(net7458));
 sg13g2_o21ai_1 _29083_ (.B1(_06795_),
    .Y(_01825_),
    .A1(_06796_),
    .A2(_06797_));
 sg13g2_nand2_1 _29084_ (.Y(_06798_),
    .A(net2773),
    .B(net8551));
 sg13g2_nor2_1 _29085_ (.A(\soc_I.qqspi_I.spi_buf[6] ),
    .B(net7459),
    .Y(_06799_));
 sg13g2_o21ai_1 _29086_ (.B1(net8556),
    .Y(_06800_),
    .A1(\soc_I.qqspi_I.spi_buf[30] ),
    .A2(net7454));
 sg13g2_o21ai_1 _29087_ (.B1(_06798_),
    .Y(_01826_),
    .A1(_06799_),
    .A2(_06800_));
 sg13g2_nand2_1 _29088_ (.Y(_06801_),
    .A(net2790),
    .B(net8551));
 sg13g2_nor2_1 _29089_ (.A(\soc_I.qqspi_I.spi_buf[7] ),
    .B(net7459),
    .Y(_06802_));
 sg13g2_o21ai_1 _29090_ (.B1(net8556),
    .Y(_06803_),
    .A1(\soc_I.qqspi_I.spi_buf[31] ),
    .A2(net7454));
 sg13g2_o21ai_1 _29091_ (.B1(_06801_),
    .Y(_01827_),
    .A1(_06802_),
    .A2(_06803_));
 sg13g2_nor2b_1 _29092_ (.A(\soc_I.rx_uart_i.state[0] ),
    .B_N(\soc_I.rx_uart_i.state[1] ),
    .Y(_06804_));
 sg13g2_and2_2 _29093_ (.A(_00249_),
    .B(_06804_),
    .X(_06805_));
 sg13g2_nand2_2 _29094_ (.Y(_06806_),
    .A(net4524),
    .B(_06804_));
 sg13g2_nor2_1 _29095_ (.A(\soc_I.rx_uart_i.bit_idx[1] ),
    .B(net9274),
    .Y(_06807_));
 sg13g2_nor3_1 _29096_ (.A(net4472),
    .B(net4545),
    .C(\soc_I.rx_uart_i.bit_idx[0] ),
    .Y(_06808_));
 sg13g2_nand2_1 _29097_ (.Y(_06809_),
    .A(_06805_),
    .B(_06808_));
 sg13g2_o21ai_1 _29098_ (.B1(net9302),
    .Y(_06810_),
    .A1(net5142),
    .A2(_06809_));
 sg13g2_a21oi_1 _29099_ (.A1(net9170),
    .A2(_06809_),
    .Y(_01828_),
    .B1(net5143));
 sg13g2_and2_1 _29100_ (.A(\soc_I.rx_uart_i.bit_idx[1] ),
    .B(net9274),
    .X(_06811_));
 sg13g2_nor2_1 _29101_ (.A(_06807_),
    .B(_06811_),
    .Y(_06812_));
 sg13g2_nor3_1 _29102_ (.A(net3095),
    .B(_06807_),
    .C(_06811_),
    .Y(_06813_));
 sg13g2_o21ai_1 _29103_ (.B1(\soc_I.rx_uart_i.bit_idx[2] ),
    .Y(_06814_),
    .A1(\soc_I.rx_uart_i.bit_idx[1] ),
    .A2(net9274));
 sg13g2_nor2_1 _29104_ (.A(_06806_),
    .B(_06808_),
    .Y(_06815_));
 sg13g2_and2_2 _29105_ (.A(_06814_),
    .B(_06815_),
    .X(_06816_));
 sg13g2_nand2_1 _29106_ (.Y(_06817_),
    .A(_06813_),
    .B(_06816_));
 sg13g2_nand2_1 _29107_ (.Y(_06818_),
    .A(net9274),
    .B(net5142));
 sg13g2_nor2_1 _29108_ (.A(net4545),
    .B(_06818_),
    .Y(_06819_));
 sg13g2_a22oi_1 _29109_ (.Y(_06820_),
    .B1(_06819_),
    .B2(_06816_),
    .A2(_06817_),
    .A1(net9288));
 sg13g2_nor2_1 _29110_ (.A(net9003),
    .B(_06820_),
    .Y(_01829_));
 sg13g2_nor2_1 _29111_ (.A(_10393_),
    .B(net9274),
    .Y(_06821_));
 sg13g2_nand2_1 _29112_ (.Y(_06822_),
    .A(_06816_),
    .B(_06821_));
 sg13g2_nor3_2 _29113_ (.A(_10393_),
    .B(net9274),
    .C(net4313),
    .Y(_06823_));
 sg13g2_a22oi_1 _29114_ (.Y(_06824_),
    .B1(net4314),
    .B2(_06816_),
    .A2(_06822_),
    .A1(net9287));
 sg13g2_nor2_1 _29115_ (.A(net9002),
    .B(_06824_),
    .Y(_01830_));
 sg13g2_nor2_1 _29116_ (.A(net3095),
    .B(_06812_),
    .Y(_06825_));
 sg13g2_nand2_1 _29117_ (.Y(_06826_),
    .A(_06816_),
    .B(_06825_));
 sg13g2_nor2_1 _29118_ (.A(_10393_),
    .B(_06818_),
    .Y(_06827_));
 sg13g2_a22oi_1 _29119_ (.Y(_06828_),
    .B1(_06827_),
    .B2(_06816_),
    .A2(_06826_),
    .A1(net9284));
 sg13g2_nor2_1 _29120_ (.A(net9002),
    .B(_06828_),
    .Y(_01831_));
 sg13g2_nor3_1 _29121_ (.A(\soc_I.rx_uart_i.bit_idx[1] ),
    .B(net9274),
    .C(net4313),
    .Y(_06829_));
 sg13g2_nand3_1 _29122_ (.B(_06805_),
    .C(_06807_),
    .A(net4472),
    .Y(_06830_));
 sg13g2_a22oi_1 _29123_ (.Y(_06831_),
    .B1(_06830_),
    .B2(net9283),
    .A2(_06829_),
    .A1(_06815_));
 sg13g2_nor2_1 _29124_ (.A(net9002),
    .B(net4473),
    .Y(_01832_));
 sg13g2_o21ai_1 _29125_ (.B1(_06809_),
    .Y(_06832_),
    .A1(_06806_),
    .A2(_06814_));
 sg13g2_nand2_1 _29126_ (.Y(_06833_),
    .A(_06813_),
    .B(_06832_));
 sg13g2_a22oi_1 _29127_ (.Y(_06834_),
    .B1(_06833_),
    .B2(net9281),
    .A2(_06832_),
    .A1(_06819_));
 sg13g2_nor2_1 _29128_ (.A(net9002),
    .B(_06834_),
    .Y(_01833_));
 sg13g2_nand2_1 _29129_ (.Y(_06835_),
    .A(_06821_),
    .B(_06832_));
 sg13g2_a22oi_1 _29130_ (.Y(_06836_),
    .B1(_06835_),
    .B2(net9278),
    .A2(_06832_),
    .A1(_06823_));
 sg13g2_nor2_1 _29131_ (.A(net9002),
    .B(_06836_),
    .Y(_01834_));
 sg13g2_or4_1 _29132_ (.A(net3095),
    .B(_06806_),
    .C(_06812_),
    .D(_06814_),
    .X(_06837_));
 sg13g2_a22oi_1 _29133_ (.Y(_06838_),
    .B1(_06837_),
    .B2(net9276),
    .A2(_06832_),
    .A1(_06827_));
 sg13g2_nor2_1 _29134_ (.A(net9002),
    .B(_06838_),
    .Y(_01835_));
 sg13g2_nand2b_1 _29135_ (.Y(_06839_),
    .B(\soc_I.rx_uart_i.rx_in_sync[2] ),
    .A_N(\soc_I.rx_uart_i.rx_in_sync[1] ));
 sg13g2_nand3_1 _29136_ (.B(_06695_),
    .C(_06839_),
    .A(_00249_),
    .Y(_06840_));
 sg13g2_and2_1 _29137_ (.A(_06707_),
    .B(_06840_),
    .X(_06841_));
 sg13g2_nand2_1 _29138_ (.Y(_06842_),
    .A(net3400),
    .B(net9303));
 sg13g2_and4_1 _29139_ (.A(net9303),
    .B(net2611),
    .C(net8800),
    .D(_06841_),
    .X(_01836_));
 sg13g2_and4_1 _29140_ (.A(net9303),
    .B(net3009),
    .C(net8800),
    .D(_06841_),
    .X(_01837_));
 sg13g2_nand2_1 _29141_ (.Y(_06843_),
    .A(\soc_I.rx_uart_i.state[0] ),
    .B(_00249_));
 sg13g2_a21oi_1 _29142_ (.A1(\soc_I.rx_uart_i.state[1] ),
    .A2(\soc_I.rx_uart_i.rx_in_sync[2] ),
    .Y(_06844_),
    .B1(_06843_));
 sg13g2_o21ai_1 _29143_ (.B1(_06844_),
    .Y(_06845_),
    .A1(\soc_I.rx_uart_i.state[1] ),
    .A2(\soc_I.rx_uart_i.rx_in_sync[2] ));
 sg13g2_and2_1 _29144_ (.A(_06840_),
    .B(_06845_),
    .X(_06846_));
 sg13g2_nand3_1 _29145_ (.B(_00249_),
    .C(_06846_),
    .A(net9303),
    .Y(_06847_));
 sg13g2_nand2b_1 _29146_ (.Y(_06848_),
    .B(_06707_),
    .A_N(_06847_));
 sg13g2_o21ai_1 _29147_ (.B1(_06848_),
    .Y(_01838_),
    .A1(_06841_),
    .A2(_06842_));
 sg13g2_o21ai_1 _29148_ (.B1(net9299),
    .Y(_06849_),
    .A1(net9274),
    .A2(_06805_));
 sg13g2_a21oi_1 _29149_ (.A1(_10394_),
    .A2(_06805_),
    .Y(_01839_),
    .B1(_06849_));
 sg13g2_o21ai_1 _29150_ (.B1(net9299),
    .Y(_06850_),
    .A1(_06806_),
    .A2(_06812_));
 sg13g2_a21oi_1 _29151_ (.A1(_10393_),
    .A2(_06806_),
    .Y(_01840_),
    .B1(_06850_));
 sg13g2_a21oi_1 _29152_ (.A1(_06805_),
    .A2(net4546),
    .Y(_06851_),
    .B1(net4472));
 sg13g2_nand3_1 _29153_ (.B(_06805_),
    .C(_06811_),
    .A(net4472),
    .Y(_06852_));
 sg13g2_nand2_1 _29154_ (.Y(_06853_),
    .A(net9299),
    .B(_06852_));
 sg13g2_nor2_1 _29155_ (.A(_06851_),
    .B(_06853_),
    .Y(_01841_));
 sg13g2_a22oi_1 _29156_ (.Y(_06854_),
    .B1(_06804_),
    .B2(_10395_),
    .A2(_06695_),
    .A1(_00249_));
 sg13g2_nand3_1 _29157_ (.B(_06843_),
    .C(_06854_),
    .A(_06697_),
    .Y(_06855_));
 sg13g2_and2_1 _29158_ (.A(_06846_),
    .B(_06855_),
    .X(_06856_));
 sg13g2_nand2_1 _29159_ (.Y(_06857_),
    .A(_06846_),
    .B(_06855_));
 sg13g2_nor2b_1 _29160_ (.A(_06695_),
    .B_N(_00249_),
    .Y(_06858_));
 sg13g2_nor2_1 _29161_ (.A(net8799),
    .B(net8797),
    .Y(_06859_));
 sg13g2_nor2_1 _29162_ (.A(net5220),
    .B(_06697_),
    .Y(_06860_));
 sg13g2_a221oi_1 _29163_ (.B2(\soc_I.div_reg[1] ),
    .C1(_06860_),
    .B1(net8672),
    .A1(\soc_I.div_reg[0] ),
    .Y(_06861_),
    .A2(net8796));
 sg13g2_a21oi_1 _29164_ (.A1(net5220),
    .A2(net8539),
    .Y(_06862_),
    .B1(net9005));
 sg13g2_o21ai_1 _29165_ (.B1(_06862_),
    .Y(_01842_),
    .A1(net8539),
    .A2(_06861_));
 sg13g2_nor2_2 _29166_ (.A(\soc_I.rx_uart_i.wait_states[1] ),
    .B(\soc_I.rx_uart_i.wait_states[0] ),
    .Y(_06863_));
 sg13g2_and2_1 _29167_ (.A(net5246),
    .B(net5220),
    .X(_06864_));
 sg13g2_o21ai_1 _29168_ (.B1(net8799),
    .Y(_06865_),
    .A1(_06863_),
    .A2(_06864_));
 sg13g2_a221oi_1 _29169_ (.B2(\soc_I.div_reg[2] ),
    .C1(net8539),
    .B1(net8671),
    .A1(\soc_I.div_reg[1] ),
    .Y(_06866_),
    .A2(net8796));
 sg13g2_o21ai_1 _29170_ (.B1(net9305),
    .Y(_06867_),
    .A1(net5246),
    .A2(net8541));
 sg13g2_a21oi_1 _29171_ (.A1(_06865_),
    .A2(_06866_),
    .Y(_01843_),
    .B1(_06867_));
 sg13g2_xor2_1 _29172_ (.B(_06863_),
    .A(_00153_),
    .X(_06868_));
 sg13g2_nor2_1 _29173_ (.A(_06697_),
    .B(_06868_),
    .Y(_06869_));
 sg13g2_a221oi_1 _29174_ (.B2(\soc_I.div_reg[3] ),
    .C1(_06869_),
    .B1(net8671),
    .A1(\soc_I.div_reg[2] ),
    .Y(_06870_),
    .A2(net8797));
 sg13g2_o21ai_1 _29175_ (.B1(net9304),
    .Y(_06871_),
    .A1(net4534),
    .A2(net8541));
 sg13g2_a21oi_1 _29176_ (.A1(net8541),
    .A2(_06870_),
    .Y(_01844_),
    .B1(_06871_));
 sg13g2_a22oi_1 _29177_ (.Y(_06872_),
    .B1(net8671),
    .B2(\soc_I.div_reg[4] ),
    .A2(net8797),
    .A1(\soc_I.div_reg[3] ));
 sg13g2_a21oi_1 _29178_ (.A1(_00153_),
    .A2(_06863_),
    .Y(_06873_),
    .B1(net4983));
 sg13g2_nand3_1 _29179_ (.B(_00153_),
    .C(_06863_),
    .A(\soc_I.rx_uart_i.wait_states[3] ),
    .Y(_06874_));
 sg13g2_a21oi_1 _29180_ (.A1(net8799),
    .A2(_06874_),
    .Y(_06875_),
    .B1(net8538));
 sg13g2_o21ai_1 _29181_ (.B1(_06872_),
    .Y(_06876_),
    .A1(_06873_),
    .A2(_06875_));
 sg13g2_o21ai_1 _29182_ (.B1(_06876_),
    .Y(_06877_),
    .A1(net4983),
    .A2(net8542));
 sg13g2_nor2_1 _29183_ (.A(net9005),
    .B(net4984),
    .Y(_01845_));
 sg13g2_and2_1 _29184_ (.A(_06699_),
    .B(_06863_),
    .X(_06878_));
 sg13g2_inv_1 _29185_ (.Y(_06879_),
    .A(_06878_));
 sg13g2_xor2_1 _29186_ (.B(_06878_),
    .A(_00154_),
    .X(_06880_));
 sg13g2_nor2_1 _29187_ (.A(_06697_),
    .B(_06880_),
    .Y(_06881_));
 sg13g2_a221oi_1 _29188_ (.B2(\soc_I.div_reg[5] ),
    .C1(_06881_),
    .B1(net8671),
    .A1(\soc_I.div_reg[4] ),
    .Y(_06882_),
    .A2(net8797));
 sg13g2_o21ai_1 _29189_ (.B1(net9304),
    .Y(_06883_),
    .A1(net5015),
    .A2(net8542));
 sg13g2_a21oi_1 _29190_ (.A1(net8541),
    .A2(_06882_),
    .Y(_01846_),
    .B1(_06883_));
 sg13g2_nand3_1 _29191_ (.B(_00154_),
    .C(_06878_),
    .A(\soc_I.rx_uart_i.wait_states[5] ),
    .Y(_06884_));
 sg13g2_a21oi_1 _29192_ (.A1(net8799),
    .A2(_06884_),
    .Y(_06885_),
    .B1(net8538));
 sg13g2_a21oi_1 _29193_ (.A1(_00154_),
    .A2(_06878_),
    .Y(_06886_),
    .B1(net5267));
 sg13g2_a22oi_1 _29194_ (.Y(_06887_),
    .B1(net8671),
    .B2(\soc_I.div_reg[6] ),
    .A2(net8798),
    .A1(\soc_I.div_reg[5] ));
 sg13g2_o21ai_1 _29195_ (.B1(_06887_),
    .Y(_06888_),
    .A1(_06885_),
    .A2(_06886_));
 sg13g2_o21ai_1 _29196_ (.B1(_06888_),
    .Y(_06889_),
    .A1(net5267),
    .A2(net8541));
 sg13g2_nor2_1 _29197_ (.A(net9005),
    .B(net5268),
    .Y(_01847_));
 sg13g2_nor3_2 _29198_ (.A(\soc_I.rx_uart_i.wait_states[5] ),
    .B(\soc_I.rx_uart_i.wait_states[4] ),
    .C(_06879_),
    .Y(_06890_));
 sg13g2_xnor2_1 _29199_ (.Y(_06891_),
    .A(_00155_),
    .B(_06890_));
 sg13g2_nand2_1 _29200_ (.Y(_06892_),
    .A(net8800),
    .B(_06891_));
 sg13g2_a221oi_1 _29201_ (.B2(\soc_I.div_reg[7] ),
    .C1(net8538),
    .B1(net8672),
    .A1(\soc_I.div_reg[6] ),
    .Y(_06893_),
    .A2(net8797));
 sg13g2_o21ai_1 _29202_ (.B1(net9304),
    .Y(_06894_),
    .A1(net4888),
    .A2(_06856_));
 sg13g2_a21oi_1 _29203_ (.A1(_06892_),
    .A2(_06893_),
    .Y(_01848_),
    .B1(_06894_));
 sg13g2_nand3_1 _29204_ (.B(_00155_),
    .C(_06890_),
    .A(\soc_I.rx_uart_i.wait_states[7] ),
    .Y(_06895_));
 sg13g2_nand2_1 _29205_ (.Y(_06896_),
    .A(net8799),
    .B(_06895_));
 sg13g2_a21oi_1 _29206_ (.A1(_00155_),
    .A2(_06890_),
    .Y(_06897_),
    .B1(net5162));
 sg13g2_a21oi_1 _29207_ (.A1(_06856_),
    .A2(_06896_),
    .Y(_06898_),
    .B1(_06897_));
 sg13g2_a221oi_1 _29208_ (.B2(\soc_I.div_reg[8] ),
    .C1(_06898_),
    .B1(net8672),
    .A1(\soc_I.div_reg[7] ),
    .Y(_06899_),
    .A2(net8798));
 sg13g2_o21ai_1 _29209_ (.B1(net9305),
    .Y(_06900_),
    .A1(net5162),
    .A2(net8542));
 sg13g2_nor2_1 _29210_ (.A(_06899_),
    .B(_06900_),
    .Y(_01849_));
 sg13g2_nand2_1 _29211_ (.Y(_06901_),
    .A(_06698_),
    .B(_06890_));
 sg13g2_nand2_1 _29212_ (.Y(_06902_),
    .A(_06702_),
    .B(_06890_));
 sg13g2_nand2_1 _29213_ (.Y(_06903_),
    .A(net4850),
    .B(_06901_));
 sg13g2_a21o_1 _29214_ (.A2(_06903_),
    .A1(_06902_),
    .B1(_06697_),
    .X(_06904_));
 sg13g2_a221oi_1 _29215_ (.B2(\soc_I.div_reg[9] ),
    .C1(net8539),
    .B1(net8672),
    .A1(\soc_I.div_reg[8] ),
    .Y(_06905_),
    .A2(net8796));
 sg13g2_o21ai_1 _29216_ (.B1(net9304),
    .Y(_06906_),
    .A1(net4850),
    .A2(net8542));
 sg13g2_a21oi_1 _29217_ (.A1(_06904_),
    .A2(_06905_),
    .Y(_01850_),
    .B1(_06906_));
 sg13g2_nor2_2 _29218_ (.A(net5109),
    .B(_06902_),
    .Y(_06907_));
 sg13g2_and2_1 _29219_ (.A(net5109),
    .B(_06902_),
    .X(_06908_));
 sg13g2_o21ai_1 _29220_ (.B1(net8799),
    .Y(_06909_),
    .A1(_06907_),
    .A2(_06908_));
 sg13g2_a221oi_1 _29221_ (.B2(\soc_I.div_reg[10] ),
    .C1(net8538),
    .B1(net8671),
    .A1(\soc_I.div_reg[9] ),
    .Y(_06910_),
    .A2(net8797));
 sg13g2_o21ai_1 _29222_ (.B1(net9303),
    .Y(_06911_),
    .A1(net5109),
    .A2(net8541));
 sg13g2_a21oi_1 _29223_ (.A1(_06909_),
    .A2(_06910_),
    .Y(_01851_),
    .B1(_06911_));
 sg13g2_xnor2_1 _29224_ (.Y(_06912_),
    .A(_00156_),
    .B(_06907_));
 sg13g2_nand2_1 _29225_ (.Y(_06913_),
    .A(net8799),
    .B(_06912_));
 sg13g2_a221oi_1 _29226_ (.B2(\soc_I.div_reg[11] ),
    .C1(net8538),
    .B1(net8671),
    .A1(\soc_I.div_reg[10] ),
    .Y(_06914_),
    .A2(net8797));
 sg13g2_o21ai_1 _29227_ (.B1(net9303),
    .Y(_06915_),
    .A1(net4759),
    .A2(net8541));
 sg13g2_a21oi_1 _29228_ (.A1(_06913_),
    .A2(_06914_),
    .Y(_01852_),
    .B1(_06915_));
 sg13g2_nand3_1 _29229_ (.B(_00156_),
    .C(_06907_),
    .A(\soc_I.rx_uart_i.wait_states[11] ),
    .Y(_06916_));
 sg13g2_a21oi_1 _29230_ (.A1(net8800),
    .A2(_06916_),
    .Y(_06917_),
    .B1(net8540));
 sg13g2_a21oi_1 _29231_ (.A1(_00156_),
    .A2(_06907_),
    .Y(_06918_),
    .B1(net5228));
 sg13g2_a22oi_1 _29232_ (.Y(_06919_),
    .B1(net8671),
    .B2(net5001),
    .A2(net8796),
    .A1(\soc_I.div_reg[11] ));
 sg13g2_o21ai_1 _29233_ (.B1(_06919_),
    .Y(_06920_),
    .A1(_06917_),
    .A2(_06918_));
 sg13g2_o21ai_1 _29234_ (.B1(_06920_),
    .Y(_06921_),
    .A1(net5228),
    .A2(net8541));
 sg13g2_nor2_1 _29235_ (.A(net9003),
    .B(net5229),
    .Y(_01853_));
 sg13g2_nand2_2 _29236_ (.Y(_06922_),
    .A(_06701_),
    .B(_06907_));
 sg13g2_xnor2_1 _29237_ (.Y(_06923_),
    .A(net5343),
    .B(_06922_));
 sg13g2_nand2_1 _29238_ (.Y(_06924_),
    .A(net8799),
    .B(_06923_));
 sg13g2_a221oi_1 _29239_ (.B2(net5313),
    .C1(net8538),
    .B1(net8672),
    .A1(net5001),
    .Y(_06925_),
    .A2(net8796));
 sg13g2_o21ai_1 _29240_ (.B1(net9305),
    .Y(_06926_),
    .A1(net5343),
    .A2(net8542));
 sg13g2_a21oi_1 _29241_ (.A1(_06924_),
    .A2(_06925_),
    .Y(_01854_),
    .B1(_06926_));
 sg13g2_nor3_2 _29242_ (.A(net5177),
    .B(\soc_I.rx_uart_i.wait_states[12] ),
    .C(_06922_),
    .Y(_06927_));
 sg13g2_o21ai_1 _29243_ (.B1(net5177),
    .Y(_06928_),
    .A1(\soc_I.rx_uart_i.wait_states[12] ),
    .A2(_06922_));
 sg13g2_inv_1 _29244_ (.Y(_06929_),
    .A(_06928_));
 sg13g2_o21ai_1 _29245_ (.B1(net8800),
    .Y(_06930_),
    .A1(_06927_),
    .A2(_06929_));
 sg13g2_a221oi_1 _29246_ (.B2(\soc_I.div_reg[14] ),
    .C1(net8538),
    .B1(net8672),
    .A1(\soc_I.div_reg[13] ),
    .Y(_06931_),
    .A2(net8796));
 sg13g2_o21ai_1 _29247_ (.B1(net9304),
    .Y(_06932_),
    .A1(net5177),
    .A2(net8542));
 sg13g2_a21oi_1 _29248_ (.A1(_06930_),
    .A2(_06931_),
    .Y(_01855_),
    .B1(_06932_));
 sg13g2_nand2_1 _29249_ (.Y(_06933_),
    .A(_00157_),
    .B(_06927_));
 sg13g2_or2_1 _29250_ (.X(_06934_),
    .B(_06927_),
    .A(_00157_));
 sg13g2_a21o_1 _29251_ (.A2(_06934_),
    .A1(_06933_),
    .B1(_06697_),
    .X(_06935_));
 sg13g2_a221oi_1 _29252_ (.B2(\soc_I.div_reg[15] ),
    .C1(net8538),
    .B1(net8672),
    .A1(\soc_I.div_reg[14] ),
    .Y(_06936_),
    .A2(net8796));
 sg13g2_o21ai_1 _29253_ (.B1(net9304),
    .Y(_06937_),
    .A1(net4866),
    .A2(net8542));
 sg13g2_a21oi_1 _29254_ (.A1(_06935_),
    .A2(_06936_),
    .Y(_01856_),
    .B1(_06937_));
 sg13g2_nor3_1 _29255_ (.A(\soc_I.rx_uart_i.wait_states[15] ),
    .B(_06697_),
    .C(_06933_),
    .Y(_06938_));
 sg13g2_a21oi_1 _29256_ (.A1(\soc_I.div_reg[15] ),
    .A2(net8796),
    .Y(_06939_),
    .B1(_06938_));
 sg13g2_a21oi_1 _29257_ (.A1(_00157_),
    .A2(_06927_),
    .Y(_06940_),
    .B1(_06697_));
 sg13g2_o21ai_1 _29258_ (.B1(net5368),
    .Y(_06941_),
    .A1(net8540),
    .A2(_06940_));
 sg13g2_o21ai_1 _29259_ (.B1(net5369),
    .Y(_06942_),
    .A1(net8540),
    .A2(_06939_));
 sg13g2_and2_1 _29260_ (.A(net9304),
    .B(_06942_),
    .X(_01857_));
 sg13g2_nand3_1 _29261_ (.B(_06701_),
    .C(_06907_),
    .A(_06700_),
    .Y(_06943_));
 sg13g2_nand3_1 _29262_ (.B(net8800),
    .C(_06846_),
    .A(net9303),
    .Y(_06944_));
 sg13g2_xnor2_1 _29263_ (.Y(_06945_),
    .A(_00290_),
    .B(_06943_));
 sg13g2_nand3_1 _29264_ (.B(net9303),
    .C(net8540),
    .A(net2633),
    .Y(_06946_));
 sg13g2_o21ai_1 _29265_ (.B1(_06946_),
    .Y(_01858_),
    .A1(_06944_),
    .A2(_06945_));
 sg13g2_o21ai_1 _29266_ (.B1(net9299),
    .Y(_06947_),
    .A1(\soc_I.rx_uart_i.fifo_i.wr_ptr[0] ),
    .A2(net8819));
 sg13g2_a21oi_1 _29267_ (.A1(_10392_),
    .A2(net8819),
    .Y(_01859_),
    .B1(_06947_));
 sg13g2_a21oi_1 _29268_ (.A1(\soc_I.rx_uart_i.fifo_i.wr_ptr[0] ),
    .A2(net8819),
    .Y(_06948_),
    .B1(net3953));
 sg13g2_nor3_1 _29269_ (.A(net9003),
    .B(_02805_),
    .C(net3954),
    .Y(_01860_));
 sg13g2_o21ai_1 _29270_ (.B1(net9299),
    .Y(_06949_),
    .A1(net9273),
    .A2(_02805_));
 sg13g2_a21oi_1 _29271_ (.A1(net9273),
    .A2(_02805_),
    .Y(_01861_),
    .B1(_06949_));
 sg13g2_a21oi_1 _29272_ (.A1(net9273),
    .A2(_02805_),
    .Y(_06950_),
    .B1(net5183));
 sg13g2_nand2_1 _29273_ (.Y(_06951_),
    .A(net9299),
    .B(net8591));
 sg13g2_nand2_1 _29274_ (.Y(_06952_),
    .A(_14123_),
    .B(_02805_));
 sg13g2_nor2_1 _29275_ (.A(net5184),
    .B(_06951_),
    .Y(_01862_));
 sg13g2_o21ai_1 _29276_ (.B1(net9298),
    .Y(_06953_),
    .A1(net3926),
    .A2(_06645_));
 sg13g2_a21oi_1 _29277_ (.A1(_10390_),
    .A2(_06645_),
    .Y(_01863_),
    .B1(_06953_));
 sg13g2_a21oi_1 _29278_ (.A1(\soc_I.rx_uart_i.fifo_i.rd_ptr[0] ),
    .A2(_06645_),
    .Y(_06954_),
    .B1(net3907));
 sg13g2_nand3_1 _29279_ (.B(net3926),
    .C(_06645_),
    .A(net3907),
    .Y(_06955_));
 sg13g2_nand2_1 _29280_ (.Y(_06956_),
    .A(net9298),
    .B(_06955_));
 sg13g2_nor2_1 _29281_ (.A(net3908),
    .B(_06956_),
    .Y(_01864_));
 sg13g2_nand2b_1 _29282_ (.Y(_06957_),
    .B(_06955_),
    .A_N(net3576));
 sg13g2_nand4_1 _29283_ (.B(\soc_I.rx_uart_i.fifo_i.rd_ptr[1] ),
    .C(\soc_I.rx_uart_i.fifo_i.rd_ptr[0] ),
    .A(net3576),
    .Y(_06958_),
    .D(_06645_));
 sg13g2_and3_1 _29284_ (.X(_01865_),
    .A(net9298),
    .B(_06957_),
    .C(net3577));
 sg13g2_o21ai_1 _29285_ (.B1(net9298),
    .Y(_06959_),
    .A1(_10389_),
    .A2(net3577));
 sg13g2_a21oi_1 _29286_ (.A1(_10389_),
    .A2(net3577),
    .Y(_01866_),
    .B1(_06959_));
 sg13g2_and2_1 _29287_ (.A(net9310),
    .B(net5),
    .X(_01867_));
 sg13g2_and2_1 _29288_ (.A(net9305),
    .B(net2728),
    .X(_01868_));
 sg13g2_and2_1 _29289_ (.A(net9299),
    .B(net4442),
    .X(_01869_));
 sg13g2_and2_1 _29290_ (.A(\soc_I.tx_uart_i.state[1] ),
    .B(\soc_I.tx_uart_i.state[0] ),
    .X(_06960_));
 sg13g2_nand2_1 _29291_ (.Y(_06961_),
    .A(\soc_I.tx_uart_i.state[1] ),
    .B(\soc_I.tx_uart_i.state[0] ));
 sg13g2_nor3_1 _29292_ (.A(\soc_I.tx_uart_i.return_state[1] ),
    .B(net3927),
    .C(net8935),
    .Y(_06962_));
 sg13g2_nor4_1 _29293_ (.A(net3615),
    .B(net4239),
    .C(net3107),
    .D(\soc_I.tx_uart_i.wait_states[6] ),
    .Y(_06963_));
 sg13g2_nor4_1 _29294_ (.A(_10589_),
    .B(\soc_I.tx_uart_i.wait_states[1] ),
    .C(net3239),
    .D(net3244),
    .Y(_06964_));
 sg13g2_nor4_1 _29295_ (.A(\soc_I.tx_uart_i.wait_states[9] ),
    .B(\soc_I.tx_uart_i.wait_states[8] ),
    .C(\soc_I.tx_uart_i.wait_states[11] ),
    .D(\soc_I.tx_uart_i.wait_states[10] ),
    .Y(_06965_));
 sg13g2_nor4_1 _29296_ (.A(\soc_I.tx_uart_i.wait_states[13] ),
    .B(\soc_I.tx_uart_i.wait_states[12] ),
    .C(\soc_I.tx_uart_i.wait_states[15] ),
    .D(\soc_I.tx_uart_i.wait_states[14] ),
    .Y(_06966_));
 sg13g2_and4_1 _29297_ (.A(_06963_),
    .B(_06964_),
    .C(_06965_),
    .D(_06966_),
    .X(_06967_));
 sg13g2_a21oi_1 _29298_ (.A1(_06962_),
    .A2(_06967_),
    .Y(_06968_),
    .B1(net4281));
 sg13g2_nor3_1 _29299_ (.A(net9005),
    .B(_13665_),
    .C(net4282),
    .Y(_01870_));
 sg13g2_o21ai_1 _29300_ (.B1(\soc_I.tx_uart_i.bit_idx[1] ),
    .Y(_06969_),
    .A1(_10386_),
    .A2(\soc_I.tx_uart_i.bit_idx[0] ));
 sg13g2_a21oi_1 _29301_ (.A1(\soc_I.tx_uart_i.tx_data_reg[7] ),
    .A2(net9272),
    .Y(_06970_),
    .B1(_06969_));
 sg13g2_mux2_1 _29302_ (.A0(\soc_I.tx_uart_i.tx_data_reg[4] ),
    .A1(\soc_I.tx_uart_i.tx_data_reg[5] ),
    .S(\soc_I.tx_uart_i.bit_idx[0] ),
    .X(_06971_));
 sg13g2_o21ai_1 _29303_ (.B1(\soc_I.tx_uart_i.bit_idx[2] ),
    .Y(_06972_),
    .A1(\soc_I.tx_uart_i.bit_idx[1] ),
    .A2(_06971_));
 sg13g2_nand2b_1 _29304_ (.Y(_06973_),
    .B(net9272),
    .A_N(\soc_I.tx_uart_i.tx_data_reg[3] ));
 sg13g2_o21ai_1 _29305_ (.B1(_06973_),
    .Y(_06974_),
    .A1(\soc_I.tx_uart_i.tx_data_reg[2] ),
    .A2(net9272));
 sg13g2_nand2b_1 _29306_ (.Y(_06975_),
    .B(net4646),
    .A_N(net9272));
 sg13g2_a21oi_1 _29307_ (.A1(\soc_I.tx_uart_i.tx_data_reg[1] ),
    .A2(net9272),
    .Y(_06976_),
    .B1(\soc_I.tx_uart_i.bit_idx[1] ));
 sg13g2_a221oi_1 _29308_ (.B2(_06976_),
    .C1(net4753),
    .B1(_06975_),
    .A1(\soc_I.tx_uart_i.bit_idx[1] ),
    .Y(_06977_),
    .A2(_06974_));
 sg13g2_nor2b_2 _29309_ (.A(\soc_I.tx_uart_i.state[1] ),
    .B_N(\soc_I.tx_uart_i.state[0] ),
    .Y(_06978_));
 sg13g2_o21ai_1 _29310_ (.B1(_06978_),
    .Y(_06979_),
    .A1(_06970_),
    .A2(_06972_));
 sg13g2_o21ai_1 _29311_ (.B1(net8935),
    .Y(_06980_),
    .A1(_06977_),
    .A2(_06979_));
 sg13g2_nand2_2 _29312_ (.Y(_06981_),
    .A(net8665),
    .B(_13169_));
 sg13g2_nor3_2 _29313_ (.A(net4281),
    .B(_13666_),
    .C(_06981_),
    .Y(_06982_));
 sg13g2_and3_2 _29314_ (.X(_06983_),
    .A(_10388_),
    .B(net8665),
    .C(_13280_));
 sg13g2_and2_1 _29315_ (.A(_13665_),
    .B(_06983_),
    .X(_06984_));
 sg13g2_a21oi_1 _29316_ (.A1(net5207),
    .A2(net8938),
    .Y(_06985_),
    .B1(net9007));
 sg13g2_o21ai_1 _29317_ (.B1(_06985_),
    .Y(_01871_),
    .A1(_06980_),
    .A2(net7396));
 sg13g2_and3_1 _29318_ (.X(_01872_),
    .A(net9333),
    .B(_12895_),
    .C(_13154_));
 sg13g2_o21ai_1 _29319_ (.B1(net9306),
    .Y(_06986_),
    .A1(net9272),
    .A2(_06978_));
 sg13g2_a21oi_1 _29320_ (.A1(_10387_),
    .A2(_06978_),
    .Y(_01873_),
    .B1(_06986_));
 sg13g2_a21oi_1 _29321_ (.A1(net9272),
    .A2(_06978_),
    .Y(_06987_),
    .B1(net4735));
 sg13g2_nand3_1 _29322_ (.B(net9272),
    .C(_06978_),
    .A(net4735),
    .Y(_06988_));
 sg13g2_nand2_1 _29323_ (.Y(_06989_),
    .A(net9306),
    .B(_06988_));
 sg13g2_nor2_1 _29324_ (.A(net4736),
    .B(_06989_),
    .Y(_01874_));
 sg13g2_xor2_1 _29325_ (.B(_06988_),
    .A(net4753),
    .X(_06990_));
 sg13g2_nor2_1 _29326_ (.A(net9006),
    .B(_06990_),
    .Y(_01875_));
 sg13g2_o21ai_1 _29327_ (.B1(net9313),
    .Y(_06991_),
    .A1(net4646),
    .A2(net7396));
 sg13g2_a21oi_1 _29328_ (.A1(_13978_),
    .A2(_06982_),
    .Y(_01876_),
    .B1(_06991_));
 sg13g2_o21ai_1 _29329_ (.B1(net9313),
    .Y(_06992_),
    .A1(net4289),
    .A2(net7396));
 sg13g2_a21oi_1 _29330_ (.A1(net8612),
    .A2(_06982_),
    .Y(_01877_),
    .B1(_06992_));
 sg13g2_o21ai_1 _29331_ (.B1(net9312),
    .Y(_06993_),
    .A1(net4513),
    .A2(_06984_));
 sg13g2_a21oi_1 _29332_ (.A1(net8610),
    .A2(_06982_),
    .Y(_01878_),
    .B1(_06993_));
 sg13g2_nand2_1 _29333_ (.Y(_06994_),
    .A(net8549),
    .B(net7396));
 sg13g2_o21ai_1 _29334_ (.B1(_06994_),
    .Y(_06995_),
    .A1(net4536),
    .A2(net7396));
 sg13g2_nor2_1 _29335_ (.A(net9005),
    .B(_06995_),
    .Y(_01879_));
 sg13g2_o21ai_1 _29336_ (.B1(net9312),
    .Y(_06996_),
    .A1(net4045),
    .A2(net7396));
 sg13g2_a21oi_1 _29337_ (.A1(net8608),
    .A2(_06982_),
    .Y(_01880_),
    .B1(_06996_));
 sg13g2_o21ai_1 _29338_ (.B1(net9312),
    .Y(_06997_),
    .A1(net4558),
    .A2(_06984_));
 sg13g2_a21oi_1 _29339_ (.A1(net8606),
    .A2(_06982_),
    .Y(_01881_),
    .B1(_06997_));
 sg13g2_o21ai_1 _29340_ (.B1(net9312),
    .Y(_06998_),
    .A1(net4419),
    .A2(_06984_));
 sg13g2_a21oi_1 _29341_ (.A1(net8604),
    .A2(_06982_),
    .Y(_01882_),
    .B1(_06998_));
 sg13g2_nand2_1 _29342_ (.Y(_06999_),
    .A(_14024_),
    .B(net7396));
 sg13g2_o21ai_1 _29343_ (.B1(_06999_),
    .Y(_07000_),
    .A1(net4657),
    .A2(net7396));
 sg13g2_nor2_1 _29344_ (.A(net9005),
    .B(_07000_),
    .Y(_01883_));
 sg13g2_nand2_1 _29345_ (.Y(_07001_),
    .A(_02802_),
    .B(_02810_));
 sg13g2_nand2_1 _29346_ (.Y(_07002_),
    .A(net2798),
    .B(_07001_));
 sg13g2_o21ai_1 _29347_ (.B1(net2799),
    .Y(_01884_),
    .A1(net9171),
    .A2(net8583));
 sg13g2_mux2_1 _29348_ (.A0(net9289),
    .A1(net4184),
    .S(net8583),
    .X(_01885_));
 sg13g2_mux2_1 _29349_ (.A0(net9286),
    .A1(net4199),
    .S(net8583),
    .X(_01886_));
 sg13g2_mux2_1 _29350_ (.A0(net9285),
    .A1(net4250),
    .S(net8583),
    .X(_01887_));
 sg13g2_mux2_1 _29351_ (.A0(net9282),
    .A1(net3939),
    .S(net8583),
    .X(_01888_));
 sg13g2_mux2_1 _29352_ (.A0(net9280),
    .A1(net4271),
    .S(net8583),
    .X(_01889_));
 sg13g2_mux2_1 _29353_ (.A0(net9278),
    .A1(net4150),
    .S(net8583),
    .X(_01890_));
 sg13g2_mux2_1 _29354_ (.A0(net9276),
    .A1(net4176),
    .S(net8583),
    .X(_01891_));
 sg13g2_nand2_1 _29355_ (.Y(_07003_),
    .A(_14126_),
    .B(_06463_));
 sg13g2_nand2_1 _29356_ (.Y(_07004_),
    .A(net2996),
    .B(net8094));
 sg13g2_o21ai_1 _29357_ (.B1(_07004_),
    .Y(_01892_),
    .A1(net7485),
    .A2(net8094));
 sg13g2_nand2_1 _29358_ (.Y(_07005_),
    .A(net3654),
    .B(net8092));
 sg13g2_o21ai_1 _29359_ (.B1(_07005_),
    .Y(_01893_),
    .A1(net7665),
    .A2(net8091));
 sg13g2_nand2_1 _29360_ (.Y(_07006_),
    .A(net3199),
    .B(net8092));
 sg13g2_o21ai_1 _29361_ (.B1(_07006_),
    .Y(_01894_),
    .A1(net7614),
    .A2(net8092));
 sg13g2_nand2_1 _29362_ (.Y(_07007_),
    .A(net3716),
    .B(net8091));
 sg13g2_o21ai_1 _29363_ (.B1(_07007_),
    .Y(_01895_),
    .A1(net7607),
    .A2(net8091));
 sg13g2_nand2_1 _29364_ (.Y(_07008_),
    .A(net3066),
    .B(net8095));
 sg13g2_o21ai_1 _29365_ (.B1(_07008_),
    .Y(_01896_),
    .A1(net7587),
    .A2(net8095));
 sg13g2_nand2_1 _29366_ (.Y(_07009_),
    .A(net3241),
    .B(net8090));
 sg13g2_o21ai_1 _29367_ (.B1(_07009_),
    .Y(_01897_),
    .A1(net7598),
    .A2(net8090));
 sg13g2_nand2_1 _29368_ (.Y(_07010_),
    .A(net3351),
    .B(net8093));
 sg13g2_o21ai_1 _29369_ (.B1(_07010_),
    .Y(_01898_),
    .A1(net7593),
    .A2(net8093));
 sg13g2_nand2_1 _29370_ (.Y(_07011_),
    .A(net2804),
    .B(net8088));
 sg13g2_o21ai_1 _29371_ (.B1(_07011_),
    .Y(_01899_),
    .A1(net7604),
    .A2(net8088));
 sg13g2_nand2_1 _29372_ (.Y(_07012_),
    .A(net2786),
    .B(net8095));
 sg13g2_o21ai_1 _29373_ (.B1(_07012_),
    .Y(_01900_),
    .A1(net7561),
    .A2(net8090));
 sg13g2_nand2_1 _29374_ (.Y(_07013_),
    .A(net2862),
    .B(net8091));
 sg13g2_o21ai_1 _29375_ (.B1(_07013_),
    .Y(_01901_),
    .A1(net7576),
    .A2(net8092));
 sg13g2_nand2_1 _29376_ (.Y(_07014_),
    .A(net3698),
    .B(net8093));
 sg13g2_o21ai_1 _29377_ (.B1(_07014_),
    .Y(_01902_),
    .A1(net7547),
    .A2(net8093));
 sg13g2_nand2_1 _29378_ (.Y(_07015_),
    .A(net2887),
    .B(net8086));
 sg13g2_o21ai_1 _29379_ (.B1(_07015_),
    .Y(_01903_),
    .A1(net7570),
    .A2(net8086));
 sg13g2_nand2_1 _29380_ (.Y(_07016_),
    .A(net2941),
    .B(net8093));
 sg13g2_o21ai_1 _29381_ (.B1(_07016_),
    .Y(_01904_),
    .A1(net7540),
    .A2(net8093));
 sg13g2_nand2_1 _29382_ (.Y(_07017_),
    .A(net3227),
    .B(net8093));
 sg13g2_o21ai_1 _29383_ (.B1(_07017_),
    .Y(_01905_),
    .A1(net7551),
    .A2(net8093));
 sg13g2_nand2_1 _29384_ (.Y(_07018_),
    .A(net2729),
    .B(net8089));
 sg13g2_o21ai_1 _29385_ (.B1(_07018_),
    .Y(_01906_),
    .A1(net7580),
    .A2(net8089));
 sg13g2_nand2_1 _29386_ (.Y(_07019_),
    .A(net3284),
    .B(net8087));
 sg13g2_o21ai_1 _29387_ (.B1(_07019_),
    .Y(_01907_),
    .A1(net7566),
    .A2(net8087));
 sg13g2_nand2_1 _29388_ (.Y(_07020_),
    .A(net3583),
    .B(net8086));
 sg13g2_o21ai_1 _29389_ (.B1(_07020_),
    .Y(_01908_),
    .A1(net7524),
    .A2(net8086));
 sg13g2_nand2_1 _29390_ (.Y(_07021_),
    .A(net3513),
    .B(net8086));
 sg13g2_o21ai_1 _29391_ (.B1(_07021_),
    .Y(_01909_),
    .A1(net7537),
    .A2(net8086));
 sg13g2_nand2_1 _29392_ (.Y(_07022_),
    .A(net3224),
    .B(net8087));
 sg13g2_o21ai_1 _29393_ (.B1(_07022_),
    .Y(_01910_),
    .A1(net7530),
    .A2(net8087));
 sg13g2_nand2_1 _29394_ (.Y(_07023_),
    .A(net3717),
    .B(net8088));
 sg13g2_o21ai_1 _29395_ (.B1(_07023_),
    .Y(_01911_),
    .A1(net7516),
    .A2(net8088));
 sg13g2_nand2_1 _29396_ (.Y(_07024_),
    .A(net2871),
    .B(net8094));
 sg13g2_o21ai_1 _29397_ (.B1(_07024_),
    .Y(_01912_),
    .A1(net7504),
    .A2(net8094));
 sg13g2_nand2_1 _29398_ (.Y(_07025_),
    .A(net3080),
    .B(net8090));
 sg13g2_o21ai_1 _29399_ (.B1(_07025_),
    .Y(_01913_),
    .A1(net7515),
    .A2(net8089));
 sg13g2_nand2_1 _29400_ (.Y(_07026_),
    .A(net3213),
    .B(net8091));
 sg13g2_o21ai_1 _29401_ (.B1(_07026_),
    .Y(_01914_),
    .A1(net7498),
    .A2(net8091));
 sg13g2_nand2_1 _29402_ (.Y(_07027_),
    .A(net2993),
    .B(net8086));
 sg13g2_o21ai_1 _29403_ (.B1(_07027_),
    .Y(_01915_),
    .A1(net7502),
    .A2(net8086));
 sg13g2_nand2_1 _29404_ (.Y(_07028_),
    .A(net2718),
    .B(net8090));
 sg13g2_o21ai_1 _29405_ (.B1(_07028_),
    .Y(_01916_),
    .A1(net7646),
    .A2(net8090));
 sg13g2_nand2_1 _29406_ (.Y(_07029_),
    .A(net3743),
    .B(net8094));
 sg13g2_o21ai_1 _29407_ (.B1(_07029_),
    .Y(_01917_),
    .A1(net7649),
    .A2(net8094));
 sg13g2_nand2_1 _29408_ (.Y(_07030_),
    .A(net3572),
    .B(net8091));
 sg13g2_o21ai_1 _29409_ (.B1(_07030_),
    .Y(_01918_),
    .A1(net7657),
    .A2(net8091));
 sg13g2_nand2_1 _29410_ (.Y(_07031_),
    .A(net3151),
    .B(net8089));
 sg13g2_o21ai_1 _29411_ (.B1(_07031_),
    .Y(_01919_),
    .A1(net7658),
    .A2(net8096));
 sg13g2_nand2_1 _29412_ (.Y(_07032_),
    .A(net2976),
    .B(net8089));
 sg13g2_o21ai_1 _29413_ (.B1(_07032_),
    .Y(_01920_),
    .A1(net7637),
    .A2(net8089));
 sg13g2_nand2_1 _29414_ (.Y(_07033_),
    .A(net3139),
    .B(net8090));
 sg13g2_o21ai_1 _29415_ (.B1(_07033_),
    .Y(_01921_),
    .A1(net7626),
    .A2(net8090));
 sg13g2_nand2_1 _29416_ (.Y(_07034_),
    .A(net2682),
    .B(net8089));
 sg13g2_o21ai_1 _29417_ (.B1(_07034_),
    .Y(_01922_),
    .A1(net7623),
    .A2(net8089));
 sg13g2_nand2_1 _29418_ (.Y(_07035_),
    .A(net3598),
    .B(net8088));
 sg13g2_o21ai_1 _29419_ (.B1(_07035_),
    .Y(_01923_),
    .A1(net7633),
    .A2(net8088));
 sg13g2_nand2b_1 _29420_ (.Y(_07036_),
    .B(_13665_),
    .A_N(_06983_));
 sg13g2_nand2_1 _29421_ (.Y(_07037_),
    .A(net9306),
    .B(_07036_));
 sg13g2_nor2b_1 _29422_ (.A(\soc_I.tx_uart_i.state[0] ),
    .B_N(\soc_I.tx_uart_i.state[1] ),
    .Y(_07038_));
 sg13g2_nand2b_1 _29423_ (.Y(_07039_),
    .B(\soc_I.tx_uart_i.state[1] ),
    .A_N(\soc_I.tx_uart_i.state[0] ));
 sg13g2_mux2_1 _29424_ (.A0(\soc_I.div_reg[1] ),
    .A1(\soc_I.tx_uart_i.wait_states[1] ),
    .S(net8937),
    .X(_07040_));
 sg13g2_nand2_1 _29425_ (.Y(_07041_),
    .A(\soc_I.div_reg[0] ),
    .B(net8934));
 sg13g2_o21ai_1 _29426_ (.B1(_07041_),
    .Y(_07042_),
    .A1(_10589_),
    .A2(net8934));
 sg13g2_or2_1 _29427_ (.X(_07043_),
    .B(_07042_),
    .A(_07040_));
 sg13g2_xor2_1 _29428_ (.B(_07042_),
    .A(_07040_),
    .X(_07044_));
 sg13g2_nand2_1 _29429_ (.Y(_07045_),
    .A(net8930),
    .B(_07044_));
 sg13g2_o21ai_1 _29430_ (.B1(_07045_),
    .Y(_07046_),
    .A1(_00106_),
    .A2(net8930));
 sg13g2_nand2_1 _29431_ (.Y(_07047_),
    .A(net4020),
    .B(net7394));
 sg13g2_o21ai_1 _29432_ (.B1(_07047_),
    .Y(_01924_),
    .A1(net7394),
    .A2(_07046_));
 sg13g2_nand2_1 _29433_ (.Y(_07048_),
    .A(net8933),
    .B(_07044_));
 sg13g2_mux2_1 _29434_ (.A0(\soc_I.div_reg[2] ),
    .A1(\soc_I.tx_uart_i.wait_states[2] ),
    .S(net8936),
    .X(_07049_));
 sg13g2_or2_1 _29435_ (.X(_07050_),
    .B(_07049_),
    .A(_07043_));
 sg13g2_xnor2_1 _29436_ (.Y(_07051_),
    .A(_07043_),
    .B(_07049_));
 sg13g2_o21ai_1 _29437_ (.B1(_07048_),
    .Y(_07052_),
    .A1(net8933),
    .A2(_07051_));
 sg13g2_nand2_1 _29438_ (.Y(_07053_),
    .A(net3244),
    .B(net7393));
 sg13g2_o21ai_1 _29439_ (.B1(_07053_),
    .Y(_01925_),
    .A1(net7393),
    .A2(_07052_));
 sg13g2_mux2_1 _29440_ (.A0(\soc_I.div_reg[3] ),
    .A1(\soc_I.tx_uart_i.wait_states[3] ),
    .S(net8937),
    .X(_07054_));
 sg13g2_xor2_1 _29441_ (.B(_07054_),
    .A(_07050_),
    .X(_07055_));
 sg13g2_nand2_1 _29442_ (.Y(_07056_),
    .A(net8930),
    .B(_07055_));
 sg13g2_o21ai_1 _29443_ (.B1(_07056_),
    .Y(_07057_),
    .A1(net8930),
    .A2(_07051_));
 sg13g2_nand2_1 _29444_ (.Y(_07058_),
    .A(net3239),
    .B(net7393));
 sg13g2_o21ai_1 _29445_ (.B1(_07058_),
    .Y(_01926_),
    .A1(net7393),
    .A2(_07057_));
 sg13g2_mux2_1 _29446_ (.A0(\soc_I.div_reg[4] ),
    .A1(\soc_I.tx_uart_i.wait_states[4] ),
    .S(net8937),
    .X(_07059_));
 sg13g2_o21ai_1 _29447_ (.B1(_07059_),
    .Y(_07060_),
    .A1(_07050_),
    .A2(_07054_));
 sg13g2_or3_1 _29448_ (.A(_07050_),
    .B(_07054_),
    .C(_07059_),
    .X(_07061_));
 sg13g2_and2_1 _29449_ (.A(net8929),
    .B(_07060_),
    .X(_07062_));
 sg13g2_a221oi_1 _29450_ (.B2(_07062_),
    .C1(net7393),
    .B1(_07061_),
    .A1(net8933),
    .Y(_07063_),
    .A2(_07055_));
 sg13g2_a21o_1 _29451_ (.A2(net7393),
    .A1(net4239),
    .B1(_07063_),
    .X(_01927_));
 sg13g2_nor4_2 _29452_ (.A(\soc_I.div_reg[3] ),
    .B(\soc_I.div_reg[2] ),
    .C(\soc_I.div_reg[1] ),
    .Y(_07064_),
    .D(\soc_I.div_reg[0] ));
 sg13g2_nand2_1 _29453_ (.Y(_07065_),
    .A(_00128_),
    .B(_07064_));
 sg13g2_o21ai_1 _29454_ (.B1(net8931),
    .Y(_07066_),
    .A1(_00128_),
    .A2(_07064_));
 sg13g2_nand2b_1 _29455_ (.Y(_07067_),
    .B(_07065_),
    .A_N(_07066_));
 sg13g2_mux2_1 _29456_ (.A0(\soc_I.div_reg[5] ),
    .A1(\soc_I.tx_uart_i.wait_states[5] ),
    .S(net8937),
    .X(_07068_));
 sg13g2_nor2_1 _29457_ (.A(_07061_),
    .B(_07068_),
    .Y(_07069_));
 sg13g2_a21o_1 _29458_ (.A2(_07068_),
    .A1(_07061_),
    .B1(net8932),
    .X(_07070_));
 sg13g2_o21ai_1 _29459_ (.B1(_07067_),
    .Y(_07071_),
    .A1(_07069_),
    .A2(_07070_));
 sg13g2_nand2_1 _29460_ (.Y(_07072_),
    .A(net3615),
    .B(net7393));
 sg13g2_o21ai_1 _29461_ (.B1(_07072_),
    .Y(_01928_),
    .A1(net7390),
    .A2(_07071_));
 sg13g2_mux2_1 _29462_ (.A0(\soc_I.div_reg[6] ),
    .A1(\soc_I.tx_uart_i.wait_states[6] ),
    .S(net8936),
    .X(_07073_));
 sg13g2_nor3_1 _29463_ (.A(_07061_),
    .B(_07068_),
    .C(_07073_),
    .Y(_07074_));
 sg13g2_xnor2_1 _29464_ (.Y(_07075_),
    .A(_07069_),
    .B(_07073_));
 sg13g2_nand2_1 _29465_ (.Y(_07076_),
    .A(net8929),
    .B(_07075_));
 sg13g2_xor2_1 _29466_ (.B(_07065_),
    .A(\soc_I.div_reg[5] ),
    .X(_07077_));
 sg13g2_a21oi_1 _29467_ (.A1(net8931),
    .A2(_07077_),
    .Y(_07078_),
    .B1(net7391));
 sg13g2_a22oi_1 _29468_ (.Y(_07079_),
    .B1(_07076_),
    .B2(_07078_),
    .A2(net7391),
    .A1(net4716));
 sg13g2_inv_1 _29469_ (.Y(_01929_),
    .A(_07079_));
 sg13g2_nand2_1 _29470_ (.Y(_07080_),
    .A(net8932),
    .B(_07075_));
 sg13g2_mux2_1 _29471_ (.A0(\soc_I.div_reg[7] ),
    .A1(\soc_I.tx_uart_i.wait_states[7] ),
    .S(net8936),
    .X(_07081_));
 sg13g2_nor2b_1 _29472_ (.A(_07081_),
    .B_N(_07074_),
    .Y(_07082_));
 sg13g2_xor2_1 _29473_ (.B(_07081_),
    .A(_07074_),
    .X(_07083_));
 sg13g2_o21ai_1 _29474_ (.B1(_07080_),
    .Y(_07084_),
    .A1(net8932),
    .A2(_07083_));
 sg13g2_nand2_1 _29475_ (.Y(_07085_),
    .A(net3107),
    .B(net7390));
 sg13g2_o21ai_1 _29476_ (.B1(_07085_),
    .Y(_01930_),
    .A1(net7392),
    .A2(_07084_));
 sg13g2_mux2_1 _29477_ (.A0(\soc_I.div_reg[8] ),
    .A1(\soc_I.tx_uart_i.wait_states[8] ),
    .S(net8936),
    .X(_07086_));
 sg13g2_nand2b_1 _29478_ (.Y(_07087_),
    .B(_07082_),
    .A_N(_07086_));
 sg13g2_xnor2_1 _29479_ (.Y(_07088_),
    .A(_07082_),
    .B(_07086_));
 sg13g2_nor2_1 _29480_ (.A(net8932),
    .B(_07088_),
    .Y(_07089_));
 sg13g2_a21oi_1 _29481_ (.A1(net8932),
    .A2(_07083_),
    .Y(_07090_),
    .B1(_07089_));
 sg13g2_nand2_1 _29482_ (.Y(_07091_),
    .A(net3016),
    .B(net7392));
 sg13g2_o21ai_1 _29483_ (.B1(_07091_),
    .Y(_01931_),
    .A1(net7392),
    .A2(_07090_));
 sg13g2_nor4_1 _29484_ (.A(\soc_I.div_reg[7] ),
    .B(\soc_I.div_reg[6] ),
    .C(\soc_I.div_reg[5] ),
    .D(\soc_I.div_reg[4] ),
    .Y(_07092_));
 sg13g2_and2_1 _29485_ (.A(_07064_),
    .B(_07092_),
    .X(_07093_));
 sg13g2_nand2_1 _29486_ (.Y(_07094_),
    .A(_00074_),
    .B(_07093_));
 sg13g2_o21ai_1 _29487_ (.B1(net8931),
    .Y(_07095_),
    .A1(_00074_),
    .A2(_07093_));
 sg13g2_nand2b_1 _29488_ (.Y(_07096_),
    .B(_07094_),
    .A_N(_07095_));
 sg13g2_mux2_1 _29489_ (.A0(\soc_I.div_reg[9] ),
    .A1(\soc_I.tx_uart_i.wait_states[9] ),
    .S(net8936),
    .X(_07097_));
 sg13g2_nor2_1 _29490_ (.A(_07087_),
    .B(_07097_),
    .Y(_07098_));
 sg13g2_a21o_1 _29491_ (.A2(_07097_),
    .A1(_07087_),
    .B1(net8932),
    .X(_07099_));
 sg13g2_o21ai_1 _29492_ (.B1(_07096_),
    .Y(_07100_),
    .A1(_07098_),
    .A2(_07099_));
 sg13g2_nand2_1 _29493_ (.Y(_07101_),
    .A(net3930),
    .B(net7390));
 sg13g2_o21ai_1 _29494_ (.B1(_07101_),
    .Y(_01932_),
    .A1(net7390),
    .A2(_07100_));
 sg13g2_nand2_1 _29495_ (.Y(_07102_),
    .A(net3527),
    .B(net7390));
 sg13g2_mux2_1 _29496_ (.A0(\soc_I.div_reg[10] ),
    .A1(\soc_I.tx_uart_i.wait_states[10] ),
    .S(net8936),
    .X(_07103_));
 sg13g2_nor3_1 _29497_ (.A(_07087_),
    .B(_07097_),
    .C(_07103_),
    .Y(_07104_));
 sg13g2_xor2_1 _29498_ (.B(_07103_),
    .A(_07098_),
    .X(_07105_));
 sg13g2_a21oi_1 _29499_ (.A1(\soc_I.div_reg[9] ),
    .A2(_07094_),
    .Y(_07106_),
    .B1(net8929));
 sg13g2_o21ai_1 _29500_ (.B1(_07106_),
    .Y(_07107_),
    .A1(\soc_I.div_reg[9] ),
    .A2(_07094_));
 sg13g2_o21ai_1 _29501_ (.B1(_07107_),
    .Y(_07108_),
    .A1(net8932),
    .A2(_07105_));
 sg13g2_o21ai_1 _29502_ (.B1(_07102_),
    .Y(_01933_),
    .A1(net7390),
    .A2(_07108_));
 sg13g2_mux2_1 _29503_ (.A0(\soc_I.div_reg[11] ),
    .A1(\soc_I.tx_uart_i.wait_states[11] ),
    .S(net8936),
    .X(_07109_));
 sg13g2_nand2b_1 _29504_ (.Y(_07110_),
    .B(_07104_),
    .A_N(_07109_));
 sg13g2_xnor2_1 _29505_ (.Y(_07111_),
    .A(_07104_),
    .B(_07109_));
 sg13g2_nand2_1 _29506_ (.Y(_07112_),
    .A(net8929),
    .B(_07111_));
 sg13g2_o21ai_1 _29507_ (.B1(_07112_),
    .Y(_07113_),
    .A1(net8929),
    .A2(_07105_));
 sg13g2_nand2_1 _29508_ (.Y(_07114_),
    .A(net3522),
    .B(net7390));
 sg13g2_o21ai_1 _29509_ (.B1(_07114_),
    .Y(_01934_),
    .A1(net7390),
    .A2(_07113_));
 sg13g2_nand2_1 _29510_ (.Y(_07115_),
    .A(net8931),
    .B(_07111_));
 sg13g2_mux2_1 _29511_ (.A0(\soc_I.div_reg[12] ),
    .A1(\soc_I.tx_uart_i.wait_states[12] ),
    .S(net8936),
    .X(_07116_));
 sg13g2_nor2_1 _29512_ (.A(_07110_),
    .B(_07116_),
    .Y(_07117_));
 sg13g2_a21o_1 _29513_ (.A2(_07116_),
    .A1(_07110_),
    .B1(net8931),
    .X(_07118_));
 sg13g2_o21ai_1 _29514_ (.B1(_07115_),
    .Y(_07119_),
    .A1(_07117_),
    .A2(_07118_));
 sg13g2_nand2_1 _29515_ (.Y(_07120_),
    .A(net3687),
    .B(net7391));
 sg13g2_o21ai_1 _29516_ (.B1(_07120_),
    .Y(_01935_),
    .A1(net7391),
    .A2(_07119_));
 sg13g2_nand2b_1 _29517_ (.Y(_07121_),
    .B(net8934),
    .A_N(\soc_I.div_reg[13] ));
 sg13g2_o21ai_1 _29518_ (.B1(_07121_),
    .Y(_07122_),
    .A1(\soc_I.tx_uart_i.wait_states[13] ),
    .A2(net8934));
 sg13g2_nand2_1 _29519_ (.Y(_07123_),
    .A(_07117_),
    .B(_07122_));
 sg13g2_nor2_1 _29520_ (.A(_07117_),
    .B(_07122_),
    .Y(_07124_));
 sg13g2_nor2_1 _29521_ (.A(net8931),
    .B(_07124_),
    .Y(_07125_));
 sg13g2_nor4_1 _29522_ (.A(\soc_I.div_reg[11] ),
    .B(\soc_I.div_reg[10] ),
    .C(\soc_I.div_reg[9] ),
    .D(\soc_I.div_reg[8] ),
    .Y(_07126_));
 sg13g2_nand3_1 _29523_ (.B(_07093_),
    .C(_07126_),
    .A(_00090_),
    .Y(_07127_));
 sg13g2_a21oi_1 _29524_ (.A1(_07093_),
    .A2(_07126_),
    .Y(_07128_),
    .B1(_00090_));
 sg13g2_nor2_1 _29525_ (.A(net8929),
    .B(_07128_),
    .Y(_07129_));
 sg13g2_a221oi_1 _29526_ (.B2(_07129_),
    .C1(net7391),
    .B1(_07127_),
    .A1(_07123_),
    .Y(_07130_),
    .A2(_07125_));
 sg13g2_a21o_1 _29527_ (.A2(net7391),
    .A1(net4195),
    .B1(_07130_),
    .X(_01936_));
 sg13g2_nand2_1 _29528_ (.Y(_07131_),
    .A(\soc_I.div_reg[14] ),
    .B(net8934));
 sg13g2_o21ai_1 _29529_ (.B1(_07131_),
    .Y(_07132_),
    .A1(_10649_),
    .A2(net8934));
 sg13g2_nor2_1 _29530_ (.A(_07123_),
    .B(_07132_),
    .Y(_07133_));
 sg13g2_xor2_1 _29531_ (.B(_07132_),
    .A(_07123_),
    .X(_07134_));
 sg13g2_or2_1 _29532_ (.X(_07135_),
    .B(_07134_),
    .A(net8933));
 sg13g2_xnor2_1 _29533_ (.Y(_07136_),
    .A(\soc_I.div_reg[13] ),
    .B(_07127_));
 sg13g2_a21oi_1 _29534_ (.A1(net8931),
    .A2(_07136_),
    .Y(_07137_),
    .B1(net7391));
 sg13g2_a22oi_1 _29535_ (.Y(_01937_),
    .B1(_07135_),
    .B2(_07137_),
    .A2(net7391),
    .A1(_10649_));
 sg13g2_nand2b_1 _29536_ (.Y(_07138_),
    .B(net8931),
    .A_N(_07134_));
 sg13g2_nand2_1 _29537_ (.Y(_07139_),
    .A(\soc_I.div_reg[15] ),
    .B(net8934));
 sg13g2_o21ai_1 _29538_ (.B1(_07139_),
    .Y(_07140_),
    .A1(_10648_),
    .A2(net8934));
 sg13g2_xor2_1 _29539_ (.B(_07140_),
    .A(_07133_),
    .X(_07141_));
 sg13g2_a21oi_1 _29540_ (.A1(net8929),
    .A2(_07141_),
    .Y(_07142_),
    .B1(net7392));
 sg13g2_a22oi_1 _29541_ (.Y(_01938_),
    .B1(_07138_),
    .B2(_07142_),
    .A2(net7392),
    .A1(_10648_));
 sg13g2_nand2_2 _29542_ (.Y(_07143_),
    .A(_14301_),
    .B(_06463_));
 sg13g2_nand2_1 _29543_ (.Y(_07144_),
    .A(net3122),
    .B(net8084));
 sg13g2_o21ai_1 _29544_ (.B1(_07144_),
    .Y(_01939_),
    .A1(net7485),
    .A2(net8084));
 sg13g2_nand2_1 _29545_ (.Y(_07145_),
    .A(net3827),
    .B(net8081));
 sg13g2_o21ai_1 _29546_ (.B1(_07145_),
    .Y(_01940_),
    .A1(net7665),
    .A2(net8081));
 sg13g2_nand2_1 _29547_ (.Y(_07146_),
    .A(net3725),
    .B(net8083));
 sg13g2_o21ai_1 _29548_ (.B1(_07146_),
    .Y(_01941_),
    .A1(net7616),
    .A2(net8083));
 sg13g2_nand2_1 _29549_ (.Y(_07147_),
    .A(net3090),
    .B(net8082));
 sg13g2_o21ai_1 _29550_ (.B1(_07147_),
    .Y(_01942_),
    .A1(net7607),
    .A2(net8081));
 sg13g2_nand2_1 _29551_ (.Y(_07148_),
    .A(net3457),
    .B(net8084));
 sg13g2_o21ai_1 _29552_ (.B1(_07148_),
    .Y(_01943_),
    .A1(net7586),
    .A2(net8084));
 sg13g2_nand2_1 _29553_ (.Y(_07149_),
    .A(net3395),
    .B(net8080));
 sg13g2_o21ai_1 _29554_ (.B1(_07149_),
    .Y(_01944_),
    .A1(net7598),
    .A2(net8080));
 sg13g2_nand2_1 _29555_ (.Y(_07150_),
    .A(net3187),
    .B(net8082));
 sg13g2_o21ai_1 _29556_ (.B1(_07150_),
    .Y(_01945_),
    .A1(net7593),
    .A2(net8082));
 sg13g2_nand2_1 _29557_ (.Y(_07151_),
    .A(net3378),
    .B(net8077));
 sg13g2_o21ai_1 _29558_ (.B1(_07151_),
    .Y(_01946_),
    .A1(net7604),
    .A2(net8077));
 sg13g2_nand2_1 _29559_ (.Y(_07152_),
    .A(net3048),
    .B(net8085));
 sg13g2_o21ai_1 _29560_ (.B1(_07152_),
    .Y(_01947_),
    .A1(net7560),
    .A2(net8085));
 sg13g2_nand2_1 _29561_ (.Y(_07153_),
    .A(net3249),
    .B(net8081));
 sg13g2_o21ai_1 _29562_ (.B1(_07153_),
    .Y(_01948_),
    .A1(net7576),
    .A2(net8083));
 sg13g2_nand2_1 _29563_ (.Y(_07154_),
    .A(net2954),
    .B(net8082));
 sg13g2_o21ai_1 _29564_ (.B1(_07154_),
    .Y(_01949_),
    .A1(net7547),
    .A2(net8082));
 sg13g2_nand2_1 _29565_ (.Y(_07155_),
    .A(net3606),
    .B(net8076));
 sg13g2_o21ai_1 _29566_ (.B1(_07155_),
    .Y(_01950_),
    .A1(net7570),
    .A2(net8076));
 sg13g2_nand2_1 _29567_ (.Y(_07156_),
    .A(net3315),
    .B(net8083));
 sg13g2_o21ai_1 _29568_ (.B1(_07156_),
    .Y(_01951_),
    .A1(net7541),
    .A2(net8083));
 sg13g2_nand2_1 _29569_ (.Y(_07157_),
    .A(net3468),
    .B(net8082));
 sg13g2_o21ai_1 _29570_ (.B1(_07157_),
    .Y(_01952_),
    .A1(net7554),
    .A2(net8082));
 sg13g2_nand2_1 _29571_ (.Y(_07158_),
    .A(net2822),
    .B(_07143_));
 sg13g2_o21ai_1 _29572_ (.B1(_07158_),
    .Y(_01953_),
    .A1(net7580),
    .A2(net8079));
 sg13g2_nand2_1 _29573_ (.Y(_07159_),
    .A(net3676),
    .B(net8077));
 sg13g2_o21ai_1 _29574_ (.B1(_07159_),
    .Y(_01954_),
    .A1(net7566),
    .A2(net8076));
 sg13g2_nand2_1 _29575_ (.Y(_07160_),
    .A(net3388),
    .B(net8076));
 sg13g2_o21ai_1 _29576_ (.B1(_07160_),
    .Y(_01955_),
    .A1(net7524),
    .A2(net8076));
 sg13g2_nand2_1 _29577_ (.Y(_07161_),
    .A(net2866),
    .B(net8076));
 sg13g2_o21ai_1 _29578_ (.B1(_07161_),
    .Y(_01956_),
    .A1(net7537),
    .A2(net8076));
 sg13g2_nand2_1 _29579_ (.Y(_07162_),
    .A(net3862),
    .B(net8077));
 sg13g2_o21ai_1 _29580_ (.B1(_07162_),
    .Y(_01957_),
    .A1(net7531),
    .A2(net8077));
 sg13g2_nand2_1 _29581_ (.Y(_07163_),
    .A(net3441),
    .B(net8077));
 sg13g2_o21ai_1 _29582_ (.B1(_07163_),
    .Y(_01958_),
    .A1(net7516),
    .A2(net8078));
 sg13g2_nand2_1 _29583_ (.Y(_07164_),
    .A(net3306),
    .B(net8084));
 sg13g2_o21ai_1 _29584_ (.B1(_07164_),
    .Y(_01959_),
    .A1(net7504),
    .A2(net8084));
 sg13g2_nand2_1 _29585_ (.Y(_07165_),
    .A(net3632),
    .B(net8080));
 sg13g2_o21ai_1 _29586_ (.B1(_07165_),
    .Y(_01960_),
    .A1(net7511),
    .A2(net8080));
 sg13g2_nand2_1 _29587_ (.Y(_07166_),
    .A(net2920),
    .B(net8081));
 sg13g2_o21ai_1 _29588_ (.B1(_07166_),
    .Y(_01961_),
    .A1(net7494),
    .A2(net8081));
 sg13g2_nand2_1 _29589_ (.Y(_07167_),
    .A(net3252),
    .B(net8078));
 sg13g2_o21ai_1 _29590_ (.B1(_07167_),
    .Y(_01962_),
    .A1(net7501),
    .A2(net8076));
 sg13g2_nand2_1 _29591_ (.Y(_07168_),
    .A(net3160),
    .B(net8080));
 sg13g2_o21ai_1 _29592_ (.B1(_07168_),
    .Y(_01963_),
    .A1(net7642),
    .A2(net8080));
 sg13g2_nand2_1 _29593_ (.Y(_07169_),
    .A(net3143),
    .B(net8084));
 sg13g2_o21ai_1 _29594_ (.B1(_07169_),
    .Y(_01964_),
    .A1(net7649),
    .A2(net8084));
 sg13g2_nand2_1 _29595_ (.Y(_07170_),
    .A(net3937),
    .B(net8081));
 sg13g2_o21ai_1 _29596_ (.B1(_07170_),
    .Y(_01965_),
    .A1(net7657),
    .A2(net8081));
 sg13g2_nand2_1 _29597_ (.Y(_07171_),
    .A(net3323),
    .B(net8079));
 sg13g2_o21ai_1 _29598_ (.B1(_07171_),
    .Y(_01966_),
    .A1(net7662),
    .A2(net8079));
 sg13g2_nand2_1 _29599_ (.Y(_07172_),
    .A(net2991),
    .B(net8079));
 sg13g2_o21ai_1 _29600_ (.B1(_07172_),
    .Y(_01967_),
    .A1(net7636),
    .A2(net8079));
 sg13g2_nand2_1 _29601_ (.Y(_07173_),
    .A(net3875),
    .B(net8080));
 sg13g2_o21ai_1 _29602_ (.B1(_07173_),
    .Y(_01968_),
    .A1(net7626),
    .A2(net8080));
 sg13g2_nand2_1 _29603_ (.Y(_07174_),
    .A(net3149),
    .B(net8079));
 sg13g2_o21ai_1 _29604_ (.B1(_07174_),
    .Y(_01969_),
    .A1(net7623),
    .A2(net8079));
 sg13g2_nand2_1 _29605_ (.Y(_07175_),
    .A(net3548),
    .B(net8077));
 sg13g2_o21ai_1 _29606_ (.B1(_07175_),
    .Y(_01970_),
    .A1(net7630),
    .A2(net8077));
 sg13g2_nor2_1 _29607_ (.A(_00286_),
    .B(net8830),
    .Y(_07176_));
 sg13g2_o21ai_1 _29608_ (.B1(net9333),
    .Y(_07177_),
    .A1(net3866),
    .A2(net8670));
 sg13g2_a21oi_1 _29609_ (.A1(_10385_),
    .A2(net8670),
    .Y(_01971_),
    .B1(net3867));
 sg13g2_o21ai_1 _29610_ (.B1(net9325),
    .Y(_07178_),
    .A1(\soc_I.spi0_I.rx_data[1] ),
    .A2(net8669));
 sg13g2_a21oi_1 _29611_ (.A1(_10384_),
    .A2(net8668),
    .Y(_01972_),
    .B1(_07178_));
 sg13g2_o21ai_1 _29612_ (.B1(net9325),
    .Y(_07179_),
    .A1(\soc_I.spi0_I.rx_data[2] ),
    .A2(net8669));
 sg13g2_a21oi_1 _29613_ (.A1(_10383_),
    .A2(net8668),
    .Y(_01973_),
    .B1(_07179_));
 sg13g2_o21ai_1 _29614_ (.B1(net9324),
    .Y(_07180_),
    .A1(\soc_I.spi0_I.rx_data[3] ),
    .A2(net8668));
 sg13g2_a21oi_1 _29615_ (.A1(_10382_),
    .A2(net8668),
    .Y(_01974_),
    .B1(_07180_));
 sg13g2_o21ai_1 _29616_ (.B1(net9324),
    .Y(_07181_),
    .A1(\soc_I.spi0_I.rx_data[4] ),
    .A2(net8668));
 sg13g2_a21oi_1 _29617_ (.A1(_10381_),
    .A2(net8668),
    .Y(_01975_),
    .B1(_07181_));
 sg13g2_o21ai_1 _29618_ (.B1(net9323),
    .Y(_07182_),
    .A1(\soc_I.spi0_I.rx_data[5] ),
    .A2(net8668));
 sg13g2_a21oi_1 _29619_ (.A1(_10380_),
    .A2(net8668),
    .Y(_01976_),
    .B1(_07182_));
 sg13g2_o21ai_1 _29620_ (.B1(net9325),
    .Y(_07183_),
    .A1(net4627),
    .A2(net8669));
 sg13g2_a21oi_1 _29621_ (.A1(_10379_),
    .A2(net8669),
    .Y(_01977_),
    .B1(_07183_));
 sg13g2_o21ai_1 _29622_ (.B1(net9333),
    .Y(_07184_),
    .A1(\soc_I.spi0_I.rx_data[7] ),
    .A2(net8670));
 sg13g2_a21oi_1 _29623_ (.A1(_10378_),
    .A2(net8670),
    .Y(_01978_),
    .B1(_07184_));
 sg13g2_nor2_2 _29624_ (.A(net9195),
    .B(\soc_I.qqspi_I.state[6] ),
    .Y(_07185_));
 sg13g2_nor2_2 _29625_ (.A(_10594_),
    .B(net8682),
    .Y(_07186_));
 sg13g2_nand2_2 _29626_ (.Y(_07187_),
    .A(net9195),
    .B(net8688));
 sg13g2_nor2_2 _29627_ (.A(net8681),
    .B(_07185_),
    .Y(_07188_));
 sg13g2_a21oi_2 _29628_ (.B1(net8681),
    .Y(_07189_),
    .A2(_07185_),
    .A1(_14272_));
 sg13g2_nand2_1 _29629_ (.Y(_07190_),
    .A(net5381),
    .B(_07189_));
 sg13g2_inv_1 _29630_ (.Y(_07191_),
    .A(_07190_));
 sg13g2_nor2_1 _29631_ (.A(net5534),
    .B(_10856_),
    .Y(_07192_));
 sg13g2_nor3_1 _29632_ (.A(_14284_),
    .B(_07190_),
    .C(_07192_),
    .Y(_07193_));
 sg13g2_o21ai_1 _29633_ (.B1(net9342),
    .Y(_07194_),
    .A1(uio_oe[1]),
    .A2(_07189_));
 sg13g2_nor2_1 _29634_ (.A(_07193_),
    .B(_07194_),
    .Y(_01979_));
 sg13g2_nand2b_1 _29635_ (.Y(_07195_),
    .B(_07192_),
    .A_N(_14284_));
 sg13g2_o21ai_1 _29636_ (.B1(net9341),
    .Y(_07196_),
    .A1(uio_oe[5]),
    .A2(_07189_));
 sg13g2_a21oi_1 _29637_ (.A1(_07191_),
    .A2(_07195_),
    .Y(_01980_),
    .B1(_07196_));
 sg13g2_nor2_1 _29638_ (.A(\soc_I.qqspi_I.state[0] ),
    .B(\soc_I.qqspi_I.state[4] ),
    .Y(_07197_));
 sg13g2_o21ai_1 _29639_ (.B1(net8683),
    .Y(_07198_),
    .A1(_00243_),
    .A2(_12558_));
 sg13g2_nor2_1 _29640_ (.A(_07197_),
    .B(_07198_),
    .Y(_07199_));
 sg13g2_or2_2 _29641_ (.X(_07200_),
    .B(_07198_),
    .A(_07197_));
 sg13g2_nor4_2 _29642_ (.A(net5394),
    .B(_12469_),
    .C(_12522_),
    .Y(_07201_),
    .D(_12552_));
 sg13g2_a21oi_1 _29643_ (.A1(uio_out[0]),
    .A2(_07200_),
    .Y(_07202_),
    .B1(net9016));
 sg13g2_o21ai_1 _29644_ (.B1(_07202_),
    .Y(_01981_),
    .A1(_07200_),
    .A2(_07201_));
 sg13g2_or4_1 _29645_ (.A(_00150_),
    .B(_12469_),
    .C(_12531_),
    .D(_12550_),
    .X(_07203_));
 sg13g2_o21ai_1 _29646_ (.B1(_07199_),
    .Y(_07204_),
    .A1(_13134_),
    .A2(_07203_));
 sg13g2_a21oi_1 _29647_ (.A1(net5513),
    .A2(_07200_),
    .Y(_07205_),
    .B1(net9016));
 sg13g2_nand2_1 _29648_ (.Y(_01982_),
    .A(_07204_),
    .B(_07205_));
 sg13g2_o21ai_1 _29649_ (.B1(_07199_),
    .Y(_07206_),
    .A1(_13135_),
    .A2(_07203_));
 sg13g2_a21oi_1 _29650_ (.A1(net5508),
    .A2(_07200_),
    .Y(_07207_),
    .B1(net9016));
 sg13g2_nand2_1 _29651_ (.Y(_01983_),
    .A(_07206_),
    .B(_07207_));
 sg13g2_nor2_1 _29652_ (.A(net3052),
    .B(net8684),
    .Y(_07208_));
 sg13g2_a22oi_1 _29653_ (.Y(_01984_),
    .B1(_07208_),
    .B2(net9341),
    .A2(_12560_),
    .A1(_10377_));
 sg13g2_nor2_1 _29654_ (.A(net3558),
    .B(net8466),
    .Y(_07209_));
 sg13g2_a21oi_1 _29655_ (.A1(net8383),
    .A2(net8466),
    .Y(_01985_),
    .B1(_07209_));
 sg13g2_nor2_1 _29656_ (.A(net3622),
    .B(net8469),
    .Y(_07210_));
 sg13g2_nor3_2 _29657_ (.A(_10925_),
    .B(_11022_),
    .C(_13289_),
    .Y(_07211_));
 sg13g2_nand3b_1 _29658_ (.B(_11021_),
    .C(_10924_),
    .Y(_07212_),
    .A_N(_13289_));
 sg13g2_nor2_1 _29659_ (.A(_00209_),
    .B(net8323),
    .Y(_07213_));
 sg13g2_xnor2_1 _29660_ (.Y(_07214_),
    .A(net8403),
    .B(_07213_));
 sg13g2_a21oi_1 _29661_ (.A1(net8469),
    .A2(_07214_),
    .Y(_01986_),
    .B1(_07210_));
 sg13g2_nor2_1 _29662_ (.A(net3313),
    .B(net8469),
    .Y(_07215_));
 sg13g2_nor2_1 _29663_ (.A(_11649_),
    .B(net8324),
    .Y(_07216_));
 sg13g2_xnor2_1 _29664_ (.Y(_07217_),
    .A(net8425),
    .B(_07216_));
 sg13g2_a21oi_1 _29665_ (.A1(net8469),
    .A2(_07217_),
    .Y(_01987_),
    .B1(_07215_));
 sg13g2_nor2_1 _29666_ (.A(net3381),
    .B(net8472),
    .Y(_07218_));
 sg13g2_nor2_1 _29667_ (.A(_11651_),
    .B(net8324),
    .Y(_07219_));
 sg13g2_xnor2_1 _29668_ (.Y(_07220_),
    .A(net8441),
    .B(_07219_));
 sg13g2_a21oi_1 _29669_ (.A1(net8472),
    .A2(_07220_),
    .Y(_01988_),
    .B1(_07218_));
 sg13g2_a21oi_1 _29670_ (.A1(net8437),
    .A2(_11651_),
    .Y(_07221_),
    .B1(net8323));
 sg13g2_xnor2_1 _29671_ (.Y(_07222_),
    .A(net8451),
    .B(_07221_));
 sg13g2_nand2_1 _29672_ (.Y(_07223_),
    .A(net2631),
    .B(net8458));
 sg13g2_o21ai_1 _29673_ (.B1(_07223_),
    .Y(_01989_),
    .A1(net8458),
    .A2(_07222_));
 sg13g2_o21ai_1 _29674_ (.B1(net8471),
    .Y(_07224_),
    .A1(net8520),
    .A2(net8328));
 sg13g2_a21oi_1 _29675_ (.A1(_04875_),
    .A2(net8329),
    .Y(_07225_),
    .B1(_07224_));
 sg13g2_a21o_1 _29676_ (.A2(net8458),
    .A1(net3772),
    .B1(_07225_),
    .X(_01990_));
 sg13g2_o21ai_1 _29677_ (.B1(net8472),
    .Y(_07226_),
    .A1(net8521),
    .A2(net8330));
 sg13g2_a21o_1 _29678_ (.A2(net8330),
    .A1(_04872_),
    .B1(_07226_),
    .X(_07227_));
 sg13g2_o21ai_1 _29679_ (.B1(_07227_),
    .Y(_01991_),
    .A1(_10609_),
    .A2(net8472));
 sg13g2_o21ai_1 _29680_ (.B1(net8472),
    .Y(_07228_),
    .A1(net8522),
    .A2(net8330));
 sg13g2_a21o_1 _29681_ (.A2(net8330),
    .A1(_04867_),
    .B1(_07228_),
    .X(_07229_));
 sg13g2_o21ai_1 _29682_ (.B1(_07229_),
    .Y(_01992_),
    .A1(_10610_),
    .A2(net8472));
 sg13g2_o21ai_1 _29683_ (.B1(net8472),
    .Y(_07230_),
    .A1(net8507),
    .A2(net8333));
 sg13g2_a21oi_1 _29684_ (.A1(_04911_),
    .A2(net8333),
    .Y(_07231_),
    .B1(_07230_));
 sg13g2_a21o_1 _29685_ (.A2(net8463),
    .A1(net3966),
    .B1(_07231_),
    .X(_01993_));
 sg13g2_o21ai_1 _29686_ (.B1(net8472),
    .Y(_07232_),
    .A1(net8505),
    .A2(net8330));
 sg13g2_a21oi_1 _29687_ (.A1(_04917_),
    .A2(net8330),
    .Y(_07233_),
    .B1(_07232_));
 sg13g2_a21o_1 _29688_ (.A2(net8463),
    .A1(net3514),
    .B1(_07233_),
    .X(_01994_));
 sg13g2_o21ai_1 _29689_ (.B1(net8474),
    .Y(_07234_),
    .A1(net8506),
    .A2(net8330));
 sg13g2_a21oi_1 _29690_ (.A1(_04923_),
    .A2(net8330),
    .Y(_07235_),
    .B1(_07234_));
 sg13g2_a21o_1 _29691_ (.A2(net8463),
    .A1(net3607),
    .B1(_07235_),
    .X(_01995_));
 sg13g2_o21ai_1 _29692_ (.B1(net8474),
    .Y(_07236_),
    .A1(net8382),
    .A2(net8331));
 sg13g2_a21oi_1 _29693_ (.A1(_04929_),
    .A2(net8331),
    .Y(_07237_),
    .B1(_07236_));
 sg13g2_a21o_1 _29694_ (.A2(net8463),
    .A1(net3967),
    .B1(_07237_),
    .X(_01996_));
 sg13g2_o21ai_1 _29695_ (.B1(net8474),
    .Y(_07238_),
    .A1(net8380),
    .A2(net8331));
 sg13g2_a21oi_1 _29696_ (.A1(_04935_),
    .A2(net8331),
    .Y(_07239_),
    .B1(_07238_));
 sg13g2_a21o_1 _29697_ (.A2(net8462),
    .A1(net3852),
    .B1(_07239_),
    .X(_01997_));
 sg13g2_nand2_1 _29698_ (.Y(_07240_),
    .A(net4871),
    .B(net8462));
 sg13g2_a21oi_1 _29699_ (.A1(net8290),
    .A2(net8326),
    .Y(_07241_),
    .B1(net8463));
 sg13g2_o21ai_1 _29700_ (.B1(_07241_),
    .Y(_07242_),
    .A1(_04942_),
    .A2(net8326));
 sg13g2_and2_1 _29701_ (.A(_07240_),
    .B(_07242_),
    .X(_07243_));
 sg13g2_inv_1 _29702_ (.Y(_01998_),
    .A(_07243_));
 sg13g2_a21oi_1 _29703_ (.A1(_11273_),
    .A2(net8326),
    .Y(_07244_),
    .B1(net8463));
 sg13g2_o21ai_1 _29704_ (.B1(_07244_),
    .Y(_07245_),
    .A1(_04947_),
    .A2(net8325));
 sg13g2_o21ai_1 _29705_ (.B1(_07245_),
    .Y(_01999_),
    .A1(_10611_),
    .A2(net8475));
 sg13g2_o21ai_1 _29706_ (.B1(net8473),
    .Y(_07246_),
    .A1(net8381),
    .A2(net8332));
 sg13g2_a21oi_1 _29707_ (.A1(_04863_),
    .A2(net8332),
    .Y(_07247_),
    .B1(_07246_));
 sg13g2_a21o_1 _29708_ (.A2(net8462),
    .A1(net3585),
    .B1(_07247_),
    .X(_02000_));
 sg13g2_a21oi_1 _29709_ (.A1(_11383_),
    .A2(net8325),
    .Y(_07248_),
    .B1(net8461));
 sg13g2_o21ai_1 _29710_ (.B1(_07248_),
    .Y(_07249_),
    .A1(_04955_),
    .A2(net8326));
 sg13g2_o21ai_1 _29711_ (.B1(_07249_),
    .Y(_02001_),
    .A1(_10612_),
    .A2(net8473));
 sg13g2_a21oi_1 _29712_ (.A1(_11416_),
    .A2(net8325),
    .Y(_07250_),
    .B1(net8459));
 sg13g2_o21ai_1 _29713_ (.B1(_07250_),
    .Y(_07251_),
    .A1(_04961_),
    .A2(net8325));
 sg13g2_o21ai_1 _29714_ (.B1(_07251_),
    .Y(_02002_),
    .A1(_10613_),
    .A2(net8473));
 sg13g2_nand2_1 _29715_ (.Y(_07252_),
    .A(net2759),
    .B(net8459));
 sg13g2_nor2_1 _29716_ (.A(_04968_),
    .B(net8325),
    .Y(_07253_));
 sg13g2_o21ai_1 _29717_ (.B1(net8469),
    .Y(_07254_),
    .A1(net8379),
    .A2(net8333));
 sg13g2_o21ai_1 _29718_ (.B1(_07252_),
    .Y(_02003_),
    .A1(_07253_),
    .A2(_07254_));
 sg13g2_o21ai_1 _29719_ (.B1(net8469),
    .Y(_07255_),
    .A1(_11404_),
    .A2(net8333));
 sg13g2_a21oi_1 _29720_ (.A1(_04974_),
    .A2(net8333),
    .Y(_07256_),
    .B1(_07255_));
 sg13g2_a21o_1 _29721_ (.A2(net8459),
    .A1(net3996),
    .B1(_07256_),
    .X(_02004_));
 sg13g2_a21oi_1 _29722_ (.A1(_11354_),
    .A2(net8325),
    .Y(_07257_),
    .B1(net8461));
 sg13g2_o21ai_1 _29723_ (.B1(_07257_),
    .Y(_07258_),
    .A1(_04860_),
    .A2(net8325));
 sg13g2_o21ai_1 _29724_ (.B1(_07258_),
    .Y(_02005_),
    .A1(_10614_),
    .A2(net8473));
 sg13g2_o21ai_1 _29725_ (.B1(net8470),
    .Y(_07259_),
    .A1(_11365_),
    .A2(net8333));
 sg13g2_a21oi_1 _29726_ (.A1(_04855_),
    .A2(net8333),
    .Y(_07260_),
    .B1(_07259_));
 sg13g2_a21o_1 _29727_ (.A2(net8459),
    .A1(net3646),
    .B1(_07260_),
    .X(_02006_));
 sg13g2_nor2_1 _29728_ (.A(_10615_),
    .B(net8473),
    .Y(_07261_));
 sg13g2_nor2_1 _29729_ (.A(_04851_),
    .B(net8324),
    .Y(_07262_));
 sg13g2_a21oi_1 _29730_ (.A1(_11326_),
    .A2(net8325),
    .Y(_07263_),
    .B1(_07262_));
 sg13g2_a21oi_1 _29731_ (.A1(net8473),
    .A2(_07263_),
    .Y(_07264_),
    .B1(_07261_));
 sg13g2_inv_1 _29732_ (.Y(_02007_),
    .A(_07264_));
 sg13g2_nor2_1 _29733_ (.A(_10616_),
    .B(net8473),
    .Y(_07265_));
 sg13g2_nor2_1 _29734_ (.A(_04847_),
    .B(net8324),
    .Y(_07266_));
 sg13g2_a21oi_2 _29735_ (.B1(_07266_),
    .Y(_07267_),
    .A2(net8324),
    .A1(_11339_));
 sg13g2_a21oi_1 _29736_ (.A1(net8473),
    .A2(_07267_),
    .Y(_07268_),
    .B1(_07265_));
 sg13g2_inv_1 _29737_ (.Y(_02008_),
    .A(_07268_));
 sg13g2_o21ai_1 _29738_ (.B1(net8470),
    .Y(_07269_),
    .A1(_11465_),
    .A2(net8329));
 sg13g2_a21oi_2 _29739_ (.B1(_07269_),
    .Y(_07270_),
    .A2(net8329),
    .A1(_04987_));
 sg13g2_a21o_1 _29740_ (.A2(net8465),
    .A1(net3854),
    .B1(_07270_),
    .X(_02009_));
 sg13g2_a21oi_1 _29741_ (.A1(_11477_),
    .A2(net8323),
    .Y(_07271_),
    .B1(net8460));
 sg13g2_o21ai_1 _29742_ (.B1(_07271_),
    .Y(_07272_),
    .A1(_04844_),
    .A2(net8323));
 sg13g2_o21ai_1 _29743_ (.B1(_07272_),
    .Y(_02010_),
    .A1(_10617_),
    .A2(_05647_));
 sg13g2_o21ai_1 _29744_ (.B1(net8470),
    .Y(_07273_),
    .A1(net8006),
    .A2(net8328));
 sg13g2_a21oi_2 _29745_ (.B1(_07273_),
    .Y(_07274_),
    .A2(net8329),
    .A1(_04995_));
 sg13g2_a21o_1 _29746_ (.A2(net8462),
    .A1(net3869),
    .B1(_07274_),
    .X(_02011_));
 sg13g2_nand2_1 _29747_ (.Y(_07275_),
    .A(net4909),
    .B(net8464));
 sg13g2_a21oi_1 _29748_ (.A1(_11453_),
    .A2(net8323),
    .Y(_07276_),
    .B1(net8455));
 sg13g2_o21ai_1 _29749_ (.B1(_07276_),
    .Y(_07277_),
    .A1(_04841_),
    .A2(net8323));
 sg13g2_and2_1 _29750_ (.A(_07275_),
    .B(_07277_),
    .X(_07278_));
 sg13g2_inv_1 _29751_ (.Y(_02012_),
    .A(_07278_));
 sg13g2_nand2_1 _29752_ (.Y(_07279_),
    .A(net4913),
    .B(net8458));
 sg13g2_a21oi_1 _29753_ (.A1(_11495_),
    .A2(net8323),
    .Y(_07280_),
    .B1(net8456));
 sg13g2_o21ai_1 _29754_ (.B1(_07280_),
    .Y(_07281_),
    .A1(_05003_),
    .A2(net8323));
 sg13g2_and2_1 _29755_ (.A(_07279_),
    .B(_07281_),
    .X(_07282_));
 sg13g2_inv_1 _29756_ (.Y(_02013_),
    .A(_07282_));
 sg13g2_o21ai_1 _29757_ (.B1(net8468),
    .Y(_07283_),
    .A1(net8007),
    .A2(net8328));
 sg13g2_a21oi_1 _29758_ (.A1(_04838_),
    .A2(net8328),
    .Y(_07284_),
    .B1(_07283_));
 sg13g2_a21o_1 _29759_ (.A2(net8458),
    .A1(net4079),
    .B1(_07284_),
    .X(_02014_));
 sg13g2_o21ai_1 _29760_ (.B1(net8468),
    .Y(_07285_),
    .A1(net8008),
    .A2(net8328));
 sg13g2_a21oi_1 _29761_ (.A1(_05012_),
    .A2(net8328),
    .Y(_07286_),
    .B1(_07285_));
 sg13g2_a21o_1 _29762_ (.A2(net8458),
    .A1(net3859),
    .B1(_07286_),
    .X(_02015_));
 sg13g2_nor3_1 _29763_ (.A(_10925_),
    .B(_13289_),
    .C(_04834_),
    .Y(_07287_));
 sg13g2_nor3_2 _29764_ (.A(_11022_),
    .B(net8457),
    .C(_07287_),
    .Y(_07288_));
 sg13g2_a21o_1 _29765_ (.A2(net8458),
    .A1(net3938),
    .B1(_07288_),
    .X(_02016_));
 sg13g2_nor2_1 _29766_ (.A(_00244_),
    .B(_12556_),
    .Y(_07289_));
 sg13g2_nor2_1 _29767_ (.A(_00243_),
    .B(_07289_),
    .Y(_07290_));
 sg13g2_nor2_1 _29768_ (.A(net8678),
    .B(_07290_),
    .Y(_07291_));
 sg13g2_nand2_1 _29769_ (.Y(_07292_),
    .A(\soc_I.qqspi_I.state[0] ),
    .B(_07291_));
 sg13g2_a22oi_1 _29770_ (.Y(_07293_),
    .B1(_07292_),
    .B2(net9268),
    .A2(_07291_),
    .A1(net4673));
 sg13g2_nor2_1 _29771_ (.A(net9019),
    .B(net4818),
    .Y(_02017_));
 sg13g2_nor2b_1 _29772_ (.A(net9256),
    .B_N(\soc_I.qqspi_I.spi_buf[31] ),
    .Y(_07294_));
 sg13g2_a21oi_1 _29773_ (.A1(net9256),
    .A2(net5578),
    .Y(_07295_),
    .B1(_07294_));
 sg13g2_o21ai_1 _29774_ (.B1(net9340),
    .Y(_07296_),
    .A1(net4584),
    .A2(net8678));
 sg13g2_a21oi_1 _29775_ (.A1(net8678),
    .A2(_07295_),
    .Y(_02018_),
    .B1(_07296_));
 sg13g2_and3_1 _29776_ (.X(_07297_),
    .A(net9256),
    .B(net9340),
    .C(net8677));
 sg13g2_a22oi_1 _29777_ (.Y(_07298_),
    .B1(_07297_),
    .B2(\soc_I.qqspi_I.spi_buf[29] ),
    .A2(_12560_),
    .A1(net3587));
 sg13g2_inv_1 _29778_ (.Y(_02019_),
    .A(net3588));
 sg13g2_a22oi_1 _29779_ (.Y(_07299_),
    .B1(_07297_),
    .B2(\soc_I.qqspi_I.spi_buf[30] ),
    .A2(net8626),
    .A1(net3102));
 sg13g2_inv_1 _29780_ (.Y(_02020_),
    .A(net3103));
 sg13g2_a22oi_1 _29781_ (.Y(_07300_),
    .B1(_07297_),
    .B2(\soc_I.qqspi_I.spi_buf[31] ),
    .A2(net8626),
    .A1(net3072));
 sg13g2_inv_1 _29782_ (.Y(_02021_),
    .A(net3073));
 sg13g2_or3_1 _29783_ (.A(_00291_),
    .B(net8665),
    .C(net8678),
    .X(_07301_));
 sg13g2_nand3b_1 _29784_ (.B(_14275_),
    .C(_07301_),
    .Y(_07302_),
    .A_N(_14271_));
 sg13g2_inv_1 _29785_ (.Y(_07303_),
    .A(net8452));
 sg13g2_nor2_1 _29786_ (.A(_00242_),
    .B(_07185_),
    .Y(_07304_));
 sg13g2_a21oi_2 _29787_ (.B1(_07188_),
    .Y(_07305_),
    .A2(net8689),
    .A1(net8666));
 sg13g2_a21oi_1 _29788_ (.A1(_13086_),
    .A2(_07304_),
    .Y(_07306_),
    .B1(_07305_));
 sg13g2_o21ai_1 _29789_ (.B1(_07306_),
    .Y(_07307_),
    .A1(_10594_),
    .A2(_14076_));
 sg13g2_a21oi_1 _29790_ (.A1(\soc_I.qqspi_I.spi_buf[20] ),
    .A2(net9264),
    .Y(_07308_),
    .B1(net8689));
 sg13g2_o21ai_1 _29791_ (.B1(_07308_),
    .Y(_07309_),
    .A1(_10375_),
    .A2(net9263));
 sg13g2_nor2b_1 _29792_ (.A(net8453),
    .B_N(_07309_),
    .Y(_07310_));
 sg13g2_a22oi_1 _29793_ (.Y(_07311_),
    .B1(_07307_),
    .B2(_07310_),
    .A2(net8453),
    .A1(net4975));
 sg13g2_nor2_1 _29794_ (.A(net9029),
    .B(net4976),
    .Y(_02022_));
 sg13g2_a21oi_1 _29795_ (.A1(_13064_),
    .A2(_07304_),
    .Y(_07312_),
    .B1(_07305_));
 sg13g2_o21ai_1 _29796_ (.B1(_07312_),
    .Y(_07313_),
    .A1(_10594_),
    .A2(_14082_));
 sg13g2_a21oi_1 _29797_ (.A1(\soc_I.qqspi_I.spi_buf[21] ),
    .A2(net9259),
    .Y(_07314_),
    .B1(net8689));
 sg13g2_o21ai_1 _29798_ (.B1(_07314_),
    .Y(_07315_),
    .A1(net9258),
    .A2(_10376_));
 sg13g2_nor2b_1 _29799_ (.A(net8452),
    .B_N(_07315_),
    .Y(_07316_));
 sg13g2_a22oi_1 _29800_ (.Y(_07317_),
    .B1(_07313_),
    .B2(_07316_),
    .A2(net8453),
    .A1(net5130));
 sg13g2_nor2_1 _29801_ (.A(net9019),
    .B(net5131),
    .Y(_02023_));
 sg13g2_nand2_1 _29802_ (.Y(_07318_),
    .A(_10595_),
    .B(_13075_));
 sg13g2_o21ai_1 _29803_ (.B1(_07318_),
    .Y(_07319_),
    .A1(_00291_),
    .A2(_14088_));
 sg13g2_mux2_1 _29804_ (.A0(\soc_I.qqspi_I.spi_buf[25] ),
    .A1(\soc_I.qqspi_I.spi_buf[22] ),
    .S(net9259),
    .X(_07320_));
 sg13g2_a22oi_1 _29805_ (.Y(_07321_),
    .B1(_07320_),
    .B2(net8680),
    .A2(_07319_),
    .A1(_07188_));
 sg13g2_o21ai_1 _29806_ (.B1(net9344),
    .Y(_07322_),
    .A1(net5417),
    .A2(_07303_));
 sg13g2_a21oi_1 _29807_ (.A1(_07303_),
    .A2(_07321_),
    .Y(_02024_),
    .B1(_07322_));
 sg13g2_nor2_1 _29808_ (.A(\soc_I.clint_I.addr[1] ),
    .B(_14297_),
    .Y(_07323_));
 sg13g2_or2_1 _29809_ (.X(_07324_),
    .B(_14092_),
    .A(_10594_));
 sg13g2_nand2_1 _29810_ (.Y(_07325_),
    .A(_10595_),
    .B(_13097_));
 sg13g2_nand3_1 _29811_ (.B(_07324_),
    .C(_07325_),
    .A(_07188_),
    .Y(_07326_));
 sg13g2_nor2b_1 _29812_ (.A(net9258),
    .B_N(\soc_I.qqspi_I.spi_buf[26] ),
    .Y(_07327_));
 sg13g2_a21oi_1 _29813_ (.A1(\soc_I.qqspi_I.spi_buf[23] ),
    .A2(net9258),
    .Y(_07328_),
    .B1(_07327_));
 sg13g2_a21oi_1 _29814_ (.A1(net8680),
    .A2(_07328_),
    .Y(_07329_),
    .B1(net8452));
 sg13g2_a22oi_1 _29815_ (.Y(_07330_),
    .B1(_07326_),
    .B2(_07329_),
    .A2(net8452),
    .A1(net5180));
 sg13g2_nor2_1 _29816_ (.A(net9019),
    .B(net5181),
    .Y(_02025_));
 sg13g2_a21oi_1 _29817_ (.A1(_10595_),
    .A2(_13120_),
    .Y(_07331_),
    .B1(_07185_));
 sg13g2_o21ai_1 _29818_ (.B1(_07331_),
    .Y(_07332_),
    .A1(_10594_),
    .A2(_14099_));
 sg13g2_nand2b_1 _29819_ (.Y(_07333_),
    .B(_07332_),
    .A_N(_07305_));
 sg13g2_nor2_1 _29820_ (.A(net9259),
    .B(net5180),
    .Y(_07334_));
 sg13g2_a21oi_1 _29821_ (.A1(net9258),
    .A2(_10376_),
    .Y(_07335_),
    .B1(_07334_));
 sg13g2_a21oi_1 _29822_ (.A1(net8680),
    .A2(_07335_),
    .Y(_07336_),
    .B1(net8453));
 sg13g2_o21ai_1 _29823_ (.B1(net9344),
    .Y(_07337_),
    .A1(net5530),
    .A2(_07303_));
 sg13g2_a21oi_1 _29824_ (.A1(_07333_),
    .A2(_07336_),
    .Y(_02026_),
    .B1(_07337_));
 sg13g2_a22oi_1 _29825_ (.Y(_07338_),
    .B1(_14105_),
    .B2(net9195),
    .A2(_13109_),
    .A1(_10595_));
 sg13g2_nor2b_1 _29826_ (.A(\soc_I.qqspi_I.is_quad ),
    .B_N(\soc_I.qqspi_I.spi_buf[28] ),
    .Y(_07339_));
 sg13g2_a21oi_1 _29827_ (.A1(net9265),
    .A2(\soc_I.qqspi_I.spi_buf[25] ),
    .Y(_07340_),
    .B1(_07339_));
 sg13g2_a221oi_1 _29828_ (.B2(net8681),
    .C1(net8453),
    .B1(_07340_),
    .A1(_07188_),
    .Y(_07341_),
    .A2(_07338_));
 sg13g2_a21oi_1 _29829_ (.A1(net5454),
    .A2(net8452),
    .Y(_07342_),
    .B1(_07341_));
 sg13g2_nor2_1 _29830_ (.A(net9019),
    .B(net5455),
    .Y(_02027_));
 sg13g2_nor2b_1 _29831_ (.A(net9258),
    .B_N(\soc_I.qqspi_I.spi_buf[29] ),
    .Y(_07343_));
 sg13g2_a21oi_1 _29832_ (.A1(net9258),
    .A2(\soc_I.qqspi_I.spi_buf[26] ),
    .Y(_07344_),
    .B1(_07343_));
 sg13g2_a21oi_1 _29833_ (.A1(net8680),
    .A2(_07344_),
    .Y(_07345_),
    .B1(net8452));
 sg13g2_a21oi_1 _29834_ (.A1(_13146_),
    .A2(_07304_),
    .Y(_07346_),
    .B1(_07305_));
 sg13g2_o21ai_1 _29835_ (.B1(_07346_),
    .Y(_07347_),
    .A1(_10594_),
    .A2(_14111_));
 sg13g2_a22oi_1 _29836_ (.Y(_07348_),
    .B1(_07345_),
    .B2(_07347_),
    .A2(net8453),
    .A1(net5442));
 sg13g2_nor2_1 _29837_ (.A(net9019),
    .B(net5443),
    .Y(_02028_));
 sg13g2_nor2b_1 _29838_ (.A(net9258),
    .B_N(\soc_I.qqspi_I.spi_buf[30] ),
    .Y(_07349_));
 sg13g2_a21oi_1 _29839_ (.A1(net9265),
    .A2(\soc_I.qqspi_I.spi_buf[27] ),
    .Y(_07350_),
    .B1(_07349_));
 sg13g2_a21oi_1 _29840_ (.A1(net8680),
    .A2(_07350_),
    .Y(_07351_),
    .B1(net8452));
 sg13g2_and2_1 _29841_ (.A(\soc_I.qqspi_I.state[6] ),
    .B(_13134_),
    .X(_07352_));
 sg13g2_a21oi_1 _29842_ (.A1(net7458),
    .A2(_07352_),
    .Y(_07353_),
    .B1(_07305_));
 sg13g2_o21ai_1 _29843_ (.B1(_07353_),
    .Y(_07354_),
    .A1(_10594_),
    .A2(_14116_));
 sg13g2_a22oi_1 _29844_ (.Y(_07355_),
    .B1(_07351_),
    .B2(_07354_),
    .A2(net8452),
    .A1(\soc_I.qqspi_I.spi_buf[31] ));
 sg13g2_nor2_1 _29845_ (.A(net9018),
    .B(_07355_),
    .Y(_02029_));
 sg13g2_o21ai_1 _29846_ (.B1(net9265),
    .Y(_07356_),
    .A1(net8681),
    .A2(_14272_));
 sg13g2_nor2b_1 _29847_ (.A(_07188_),
    .B_N(_07356_),
    .Y(_07357_));
 sg13g2_nor2_1 _29848_ (.A(net9018),
    .B(_07357_),
    .Y(_02030_));
 sg13g2_nor2_1 _29849_ (.A(net9006),
    .B(_13163_),
    .Y(_02031_));
 sg13g2_and2_1 _29850_ (.A(net9323),
    .B(_13170_),
    .X(_02032_));
 sg13g2_nor2_2 _29851_ (.A(_10856_),
    .B(_13163_),
    .Y(_07358_));
 sg13g2_nor4_2 _29852_ (.A(net9254),
    .B(_10856_),
    .C(_13157_),
    .Y(_07359_),
    .D(_13264_));
 sg13g2_and2_2 _29853_ (.A(net8665),
    .B(_13279_),
    .X(_07360_));
 sg13g2_o21ai_1 _29854_ (.B1(net9312),
    .Y(_07361_),
    .A1(net5398),
    .A2(net7426));
 sg13g2_a21oi_1 _29855_ (.A1(_13978_),
    .A2(net7426),
    .Y(_02033_),
    .B1(_07361_));
 sg13g2_o21ai_1 _29856_ (.B1(net9312),
    .Y(_07362_),
    .A1(net5359),
    .A2(net7426));
 sg13g2_a21oi_1 _29857_ (.A1(net8612),
    .A2(net7426),
    .Y(_02034_),
    .B1(_07362_));
 sg13g2_o21ai_1 _29858_ (.B1(net9307),
    .Y(_07363_),
    .A1(net5436),
    .A2(net7428));
 sg13g2_a21oi_1 _29859_ (.A1(net8610),
    .A2(net7428),
    .Y(_02035_),
    .B1(_07363_));
 sg13g2_o21ai_1 _29860_ (.B1(net9312),
    .Y(_07364_),
    .A1(net5434),
    .A2(net7426));
 sg13g2_a21oi_1 _29861_ (.A1(net8549),
    .A2(net7427),
    .Y(_02036_),
    .B1(_07364_));
 sg13g2_o21ai_1 _29862_ (.B1(net9312),
    .Y(_07365_),
    .A1(net5421),
    .A2(net7426));
 sg13g2_a21oi_1 _29863_ (.A1(net8608),
    .A2(net7395),
    .Y(_02037_),
    .B1(_07365_));
 sg13g2_o21ai_1 _29864_ (.B1(net9310),
    .Y(_07366_),
    .A1(net5467),
    .A2(net7430));
 sg13g2_a21oi_1 _29865_ (.A1(net8606),
    .A2(net7430),
    .Y(_02038_),
    .B1(_07366_));
 sg13g2_o21ai_1 _29866_ (.B1(net9307),
    .Y(_07367_),
    .A1(net5327),
    .A2(net7428));
 sg13g2_a21oi_1 _29867_ (.A1(net8604),
    .A2(net7428),
    .Y(_02039_),
    .B1(_07367_));
 sg13g2_o21ai_1 _29868_ (.B1(net9307),
    .Y(_07368_),
    .A1(net5319),
    .A2(net7426));
 sg13g2_a21oi_1 _29869_ (.A1(_14024_),
    .A2(net7426),
    .Y(_02040_),
    .B1(_07368_));
 sg13g2_o21ai_1 _29870_ (.B1(net9307),
    .Y(_07369_),
    .A1(net5271),
    .A2(net7427));
 sg13g2_a21oi_1 _29871_ (.A1(_13979_),
    .A2(net7395),
    .Y(_02041_),
    .B1(_07369_));
 sg13g2_o21ai_1 _29872_ (.B1(net9307),
    .Y(_07370_),
    .A1(net5384),
    .A2(net7429));
 sg13g2_a21oi_1 _29873_ (.A1(_13988_),
    .A2(net7429),
    .Y(_02042_),
    .B1(_07370_));
 sg13g2_o21ai_1 _29874_ (.B1(net9307),
    .Y(_07371_),
    .A1(net5253),
    .A2(net7427));
 sg13g2_a21oi_1 _29875_ (.A1(_13995_),
    .A2(net7427),
    .Y(_02043_),
    .B1(_07371_));
 sg13g2_o21ai_1 _29876_ (.B1(net9307),
    .Y(_07372_),
    .A1(net5232),
    .A2(net7429));
 sg13g2_a21oi_1 _29877_ (.A1(_14001_),
    .A2(net7429),
    .Y(_02044_),
    .B1(_07372_));
 sg13g2_o21ai_1 _29878_ (.B1(net9307),
    .Y(_07373_),
    .A1(net5001),
    .A2(net7427));
 sg13g2_a21oi_1 _29879_ (.A1(_14007_),
    .A2(net7427),
    .Y(_02045_),
    .B1(_07373_));
 sg13g2_o21ai_1 _29880_ (.B1(net9309),
    .Y(_07374_),
    .A1(net5313),
    .A2(net7427));
 sg13g2_a21oi_1 _29881_ (.A1(_14014_),
    .A2(net7395),
    .Y(_02046_),
    .B1(_07374_));
 sg13g2_o21ai_1 _29882_ (.B1(net9309),
    .Y(_07375_),
    .A1(net5250),
    .A2(net7429));
 sg13g2_a21oi_1 _29883_ (.A1(_14020_),
    .A2(net7429),
    .Y(_02047_),
    .B1(_07375_));
 sg13g2_o21ai_1 _29884_ (.B1(net9322),
    .Y(_07376_),
    .A1(net5367),
    .A2(net7430));
 sg13g2_a21oi_1 _29885_ (.A1(_14029_),
    .A2(net7418),
    .Y(_02048_),
    .B1(_07376_));
 sg13g2_o21ai_1 _29886_ (.B1(net9327),
    .Y(_07377_),
    .A1(net5457),
    .A2(net7433));
 sg13g2_a21oi_1 _29887_ (.A1(_14037_),
    .A2(net7418),
    .Y(_02049_),
    .B1(_07377_));
 sg13g2_o21ai_1 _29888_ (.B1(net9327),
    .Y(_07378_),
    .A1(net5375),
    .A2(net7433));
 sg13g2_a21oi_1 _29889_ (.A1(_14041_),
    .A2(net7418),
    .Y(_02050_),
    .B1(_07378_));
 sg13g2_nand2_1 _29890_ (.Y(_07379_),
    .A(_14046_),
    .B(net7418));
 sg13g2_o21ai_1 _29891_ (.B1(_07379_),
    .Y(_07380_),
    .A1(net5146),
    .A2(_07358_));
 sg13g2_nor2_1 _29892_ (.A(net9013),
    .B(_07380_),
    .Y(_02051_));
 sg13g2_o21ai_1 _29893_ (.B1(net9328),
    .Y(_07381_),
    .A1(net5292),
    .A2(net7431));
 sg13g2_a21oi_1 _29894_ (.A1(_14051_),
    .A2(_07360_),
    .Y(_02052_),
    .B1(_07381_));
 sg13g2_o21ai_1 _29895_ (.B1(net9339),
    .Y(_07382_),
    .A1(net4420),
    .A2(net7432));
 sg13g2_a21oi_1 _29896_ (.A1(_14056_),
    .A2(net7418),
    .Y(_02053_),
    .B1(_07382_));
 sg13g2_nand2_1 _29897_ (.Y(_07383_),
    .A(_14060_),
    .B(_07360_));
 sg13g2_o21ai_1 _29898_ (.B1(_07383_),
    .Y(_07384_),
    .A1(net5416),
    .A2(net7395));
 sg13g2_nor2_1 _29899_ (.A(net9013),
    .B(_07384_),
    .Y(_02054_));
 sg13g2_o21ai_1 _29900_ (.B1(net9339),
    .Y(_07385_),
    .A1(net5185),
    .A2(net7431));
 sg13g2_a21oi_1 _29901_ (.A1(_14065_),
    .A2(net7431),
    .Y(_02055_),
    .B1(_07385_));
 sg13g2_o21ai_1 _29902_ (.B1(net9339),
    .Y(_07386_),
    .A1(net5074),
    .A2(net7431));
 sg13g2_a21oi_1 _29903_ (.A1(_14070_),
    .A2(_07360_),
    .Y(_02056_),
    .B1(_07386_));
 sg13g2_o21ai_1 _29904_ (.B1(net9328),
    .Y(_07387_),
    .A1(net4454),
    .A2(net7432));
 sg13g2_a21oi_1 _29905_ (.A1(_14076_),
    .A2(net7418),
    .Y(_02057_),
    .B1(_07387_));
 sg13g2_o21ai_1 _29906_ (.B1(net9333),
    .Y(_07388_),
    .A1(net5252),
    .A2(net7432));
 sg13g2_a21oi_1 _29907_ (.A1(_14082_),
    .A2(net7395),
    .Y(_02058_),
    .B1(_07388_));
 sg13g2_o21ai_1 _29908_ (.B1(net9328),
    .Y(_07389_),
    .A1(net5033),
    .A2(net7432));
 sg13g2_a21oi_1 _29909_ (.A1(_14088_),
    .A2(net7432),
    .Y(_02059_),
    .B1(_07389_));
 sg13g2_o21ai_1 _29910_ (.B1(net9328),
    .Y(_07390_),
    .A1(net5047),
    .A2(net7431));
 sg13g2_a21oi_1 _29911_ (.A1(_14092_),
    .A2(net7418),
    .Y(_02060_),
    .B1(_07390_));
 sg13g2_o21ai_1 _29912_ (.B1(net9329),
    .Y(_07391_),
    .A1(net4418),
    .A2(net7431));
 sg13g2_a21oi_1 _29913_ (.A1(_14099_),
    .A2(net7395),
    .Y(_02061_),
    .B1(_07391_));
 sg13g2_o21ai_1 _29914_ (.B1(net9327),
    .Y(_07392_),
    .A1(net5260),
    .A2(net7433));
 sg13g2_a21oi_1 _29915_ (.A1(_14104_),
    .A2(net7395),
    .Y(_02062_),
    .B1(_07392_));
 sg13g2_o21ai_1 _29916_ (.B1(net9327),
    .Y(_07393_),
    .A1(net5017),
    .A2(net7431));
 sg13g2_a21oi_1 _29917_ (.A1(_14111_),
    .A2(net7418),
    .Y(_02063_),
    .B1(_07393_));
 sg13g2_o21ai_1 _29918_ (.B1(net9328),
    .Y(_07394_),
    .A1(net5148),
    .A2(net7431));
 sg13g2_a21oi_1 _29919_ (.A1(_14116_),
    .A2(net7395),
    .Y(_02064_),
    .B1(_07394_));
 sg13g2_nor2_1 _29920_ (.A(net9014),
    .B(_06981_),
    .Y(_02065_));
 sg13g2_and2_2 _29921_ (.A(net8665),
    .B(_13170_),
    .X(_07395_));
 sg13g2_nor2_1 _29922_ (.A(_10856_),
    .B(_13276_),
    .Y(_07396_));
 sg13g2_o21ai_1 _29923_ (.B1(net9333),
    .Y(_07397_),
    .A1(net5550),
    .A2(net7416));
 sg13g2_a21oi_1 _29924_ (.A1(_13978_),
    .A2(net7416),
    .Y(_02066_),
    .B1(_07397_));
 sg13g2_o21ai_1 _29925_ (.B1(net9323),
    .Y(_07398_),
    .A1(net5210),
    .A2(net7408));
 sg13g2_a21oi_1 _29926_ (.A1(net8612),
    .A2(net7408),
    .Y(_02067_),
    .B1(_07398_));
 sg13g2_o21ai_1 _29927_ (.B1(net9323),
    .Y(_07399_),
    .A1(net5153),
    .A2(net7409));
 sg13g2_a21oi_1 _29928_ (.A1(net8610),
    .A2(_07395_),
    .Y(_02068_),
    .B1(_07399_));
 sg13g2_o21ai_1 _29929_ (.B1(net9323),
    .Y(_07400_),
    .A1(net5037),
    .A2(net7408));
 sg13g2_a21oi_1 _29930_ (.A1(net8549),
    .A2(net7408),
    .Y(_02069_),
    .B1(_07400_));
 sg13g2_o21ai_1 _29931_ (.B1(net9313),
    .Y(_07401_),
    .A1(net4939),
    .A2(net7408));
 sg13g2_a21oi_1 _29932_ (.A1(net8608),
    .A2(_07395_),
    .Y(_02070_),
    .B1(_07401_));
 sg13g2_o21ai_1 _29933_ (.B1(net9313),
    .Y(_07402_),
    .A1(net4890),
    .A2(net7408));
 sg13g2_a21oi_1 _29934_ (.A1(net8606),
    .A2(net7408),
    .Y(_02071_),
    .B1(_07402_));
 sg13g2_o21ai_1 _29935_ (.B1(net9313),
    .Y(_07403_),
    .A1(net5108),
    .A2(net7408));
 sg13g2_a21oi_1 _29936_ (.A1(net8604),
    .A2(_07395_),
    .Y(_02072_),
    .B1(_07403_));
 sg13g2_o21ai_1 _29937_ (.B1(net9323),
    .Y(_07404_),
    .A1(net5009),
    .A2(net7409));
 sg13g2_a21oi_1 _29938_ (.A1(_14024_),
    .A2(net7409),
    .Y(_02073_),
    .B1(_07404_));
 sg13g2_o21ai_1 _29939_ (.B1(net9313),
    .Y(_07405_),
    .A1(net4767),
    .A2(net7410));
 sg13g2_a21oi_1 _29940_ (.A1(_13979_),
    .A2(net7410),
    .Y(_02074_),
    .B1(_07405_));
 sg13g2_nand2_1 _29941_ (.Y(_07406_),
    .A(_13988_),
    .B(net7407));
 sg13g2_o21ai_1 _29942_ (.B1(_07406_),
    .Y(_07407_),
    .A1(net5282),
    .A2(net7407));
 sg13g2_nor2_1 _29943_ (.A(net9006),
    .B(_07407_),
    .Y(_02075_));
 sg13g2_o21ai_1 _29944_ (.B1(net9323),
    .Y(_07408_),
    .A1(net5234),
    .A2(net7409));
 sg13g2_a21oi_1 _29945_ (.A1(_13995_),
    .A2(_07395_),
    .Y(_02076_),
    .B1(_07408_));
 sg13g2_o21ai_1 _29946_ (.B1(net9310),
    .Y(_07409_),
    .A1(net5358),
    .A2(net7407));
 sg13g2_a21oi_1 _29947_ (.A1(_14001_),
    .A2(net7407),
    .Y(_02077_),
    .B1(_07409_));
 sg13g2_o21ai_1 _29948_ (.B1(net9313),
    .Y(_07410_),
    .A1(net5123),
    .A2(net7410));
 sg13g2_a21oi_1 _29949_ (.A1(_14007_),
    .A2(net7410),
    .Y(_02078_),
    .B1(_07410_));
 sg13g2_o21ai_1 _29950_ (.B1(net9310),
    .Y(_07411_),
    .A1(net5304),
    .A2(net7407));
 sg13g2_a21oi_1 _29951_ (.A1(_14014_),
    .A2(net7407),
    .Y(_02079_),
    .B1(_07411_));
 sg13g2_nand2_1 _29952_ (.Y(_07412_),
    .A(_14020_),
    .B(net7407));
 sg13g2_o21ai_1 _29953_ (.B1(_07412_),
    .Y(_07413_),
    .A1(net5276),
    .A2(net7407));
 sg13g2_nor2_1 _29954_ (.A(net9006),
    .B(_07413_),
    .Y(_02080_));
 sg13g2_nand2_1 _29955_ (.Y(_07414_),
    .A(_14029_),
    .B(net7411));
 sg13g2_o21ai_1 _29956_ (.B1(_07414_),
    .Y(_07415_),
    .A1(net5364),
    .A2(net7411));
 sg13g2_nor2_1 _29957_ (.A(net9014),
    .B(_07415_),
    .Y(_02081_));
 sg13g2_o21ai_1 _29958_ (.B1(net9337),
    .Y(_07416_),
    .A1(net4438),
    .A2(net7412));
 sg13g2_a21oi_1 _29959_ (.A1(_14037_),
    .A2(net7412),
    .Y(_02082_),
    .B1(_07416_));
 sg13g2_o21ai_1 _29960_ (.B1(net9337),
    .Y(_07417_),
    .A1(net4341),
    .A2(net7412));
 sg13g2_a21oi_1 _29961_ (.A1(_14041_),
    .A2(net7412),
    .Y(_02083_),
    .B1(_07417_));
 sg13g2_o21ai_1 _29962_ (.B1(net9315),
    .Y(_07418_),
    .A1(net4523),
    .A2(net7417));
 sg13g2_a21oi_1 _29963_ (.A1(_14046_),
    .A2(net7417),
    .Y(_02084_),
    .B1(_07418_));
 sg13g2_o21ai_1 _29964_ (.B1(net9339),
    .Y(_07419_),
    .A1(net4563),
    .A2(net7413));
 sg13g2_a21oi_1 _29965_ (.A1(_14051_),
    .A2(net7413),
    .Y(_02085_),
    .B1(_07419_));
 sg13g2_o21ai_1 _29966_ (.B1(net9329),
    .Y(_07420_),
    .A1(net4701),
    .A2(net7415));
 sg13g2_a21oi_1 _29967_ (.A1(_14056_),
    .A2(net7415),
    .Y(_02086_),
    .B1(_07420_));
 sg13g2_o21ai_1 _29968_ (.B1(net9337),
    .Y(_07421_),
    .A1(net4369),
    .A2(net7413));
 sg13g2_a21oi_1 _29969_ (.A1(_14060_),
    .A2(net7412),
    .Y(_02087_),
    .B1(_07421_));
 sg13g2_o21ai_1 _29970_ (.B1(net9339),
    .Y(_07422_),
    .A1(net4639),
    .A2(net7413));
 sg13g2_a21oi_1 _29971_ (.A1(_14065_),
    .A2(net7412),
    .Y(_02088_),
    .B1(_07422_));
 sg13g2_o21ai_1 _29972_ (.B1(net9337),
    .Y(_07423_),
    .A1(net4632),
    .A2(net7412));
 sg13g2_a21oi_1 _29973_ (.A1(_14070_),
    .A2(net7412),
    .Y(_02089_),
    .B1(_07423_));
 sg13g2_o21ai_1 _29974_ (.B1(net9339),
    .Y(_07424_),
    .A1(net4593),
    .A2(net7415));
 sg13g2_a21oi_1 _29975_ (.A1(_14076_),
    .A2(net7415),
    .Y(_02090_),
    .B1(_07424_));
 sg13g2_o21ai_1 _29976_ (.B1(net9340),
    .Y(_07425_),
    .A1(net4444),
    .A2(net7415));
 sg13g2_a21oi_1 _29977_ (.A1(_14082_),
    .A2(net7415),
    .Y(_02091_),
    .B1(_07425_));
 sg13g2_o21ai_1 _29978_ (.B1(net9329),
    .Y(_07426_),
    .A1(net4815),
    .A2(net7415));
 sg13g2_a21oi_1 _29979_ (.A1(_14088_),
    .A2(net7415),
    .Y(_02092_),
    .B1(_07426_));
 sg13g2_o21ai_1 _29980_ (.B1(net9329),
    .Y(_07427_),
    .A1(net4507),
    .A2(net7413));
 sg13g2_a21oi_1 _29981_ (.A1(_14092_),
    .A2(net7413),
    .Y(_02093_),
    .B1(_07427_));
 sg13g2_o21ai_1 _29982_ (.B1(net9330),
    .Y(_07428_),
    .A1(net4392),
    .A2(net7414));
 sg13g2_a21oi_1 _29983_ (.A1(_14099_),
    .A2(net7414),
    .Y(_02094_),
    .B1(_07428_));
 sg13g2_o21ai_1 _29984_ (.B1(net9327),
    .Y(_07429_),
    .A1(net4312),
    .A2(net7416));
 sg13g2_a21oi_1 _29985_ (.A1(_14104_),
    .A2(net7416),
    .Y(_02095_),
    .B1(_07429_));
 sg13g2_o21ai_1 _29986_ (.B1(net9330),
    .Y(_07430_),
    .A1(net4688),
    .A2(net7414));
 sg13g2_a21oi_1 _29987_ (.A1(_14111_),
    .A2(net7414),
    .Y(_02096_),
    .B1(_07430_));
 sg13g2_o21ai_1 _29988_ (.B1(net9340),
    .Y(_07431_),
    .A1(net4361),
    .A2(net7416));
 sg13g2_a21oi_1 _29989_ (.A1(_14116_),
    .A2(net7416),
    .Y(_02097_),
    .B1(_07431_));
 sg13g2_nor2_1 _29990_ (.A(net9016),
    .B(_13166_),
    .Y(_02098_));
 sg13g2_nor4_2 _29991_ (.A(net9016),
    .B(net9245),
    .C(net8665),
    .Y(_02099_),
    .D(_13168_));
 sg13g2_nand2_1 _29992_ (.Y(_07432_),
    .A(_14122_),
    .B(_02802_));
 sg13g2_nand2_1 _29993_ (.Y(_07433_),
    .A(net2620),
    .B(_07432_));
 sg13g2_o21ai_1 _29994_ (.B1(net2621),
    .Y(_02100_),
    .A1(net9171),
    .A2(net8537));
 sg13g2_mux2_1 _29995_ (.A0(net9289),
    .A1(net4146),
    .S(net8537),
    .X(_02101_));
 sg13g2_mux2_1 _29996_ (.A0(net9286),
    .A1(net4006),
    .S(net8537),
    .X(_02102_));
 sg13g2_mux2_1 _29997_ (.A0(net9285),
    .A1(net3691),
    .S(net8537),
    .X(_02103_));
 sg13g2_mux2_1 _29998_ (.A0(net9282),
    .A1(net4209),
    .S(net8537),
    .X(_02104_));
 sg13g2_mux2_1 _29999_ (.A0(net9280),
    .A1(net3806),
    .S(net8537),
    .X(_02105_));
 sg13g2_mux2_1 _30000_ (.A0(net9278),
    .A1(net3620),
    .S(net8537),
    .X(_02106_));
 sg13g2_mux2_1 _30001_ (.A0(net9276),
    .A1(net3532),
    .S(net8537),
    .X(_02107_));
 sg13g2_o21ai_1 _30002_ (.B1(net9363),
    .Y(_07434_),
    .A1(net4377),
    .A2(net7765));
 sg13g2_a21oi_1 _30003_ (.A1(_04070_),
    .A2(net7765),
    .Y(_02108_),
    .B1(_07434_));
 sg13g2_o21ai_1 _30004_ (.B1(net9382),
    .Y(_07435_),
    .A1(net4448),
    .A2(net7762));
 sg13g2_a21oi_1 _30005_ (.A1(_03841_),
    .A2(net7762),
    .Y(_02109_),
    .B1(_07435_));
 sg13g2_o21ai_1 _30006_ (.B1(net9373),
    .Y(_07436_),
    .A1(net4310),
    .A2(net7767));
 sg13g2_a21oi_1 _30007_ (.A1(_03862_),
    .A2(net7767),
    .Y(_02110_),
    .B1(_07436_));
 sg13g2_o21ai_1 _30008_ (.B1(net9379),
    .Y(_07437_),
    .A1(net4443),
    .A2(net7767));
 sg13g2_a21oi_1 _30009_ (.A1(_03871_),
    .A2(net7767),
    .Y(_02111_),
    .B1(_07437_));
 sg13g2_o21ai_1 _30010_ (.B1(net9379),
    .Y(_07438_),
    .A1(net4504),
    .A2(net7767));
 sg13g2_a21oi_1 _30011_ (.A1(_03889_),
    .A2(net7767),
    .Y(_02112_),
    .B1(_07438_));
 sg13g2_o21ai_1 _30012_ (.B1(net9370),
    .Y(_07439_),
    .A1(net4520),
    .A2(net7767));
 sg13g2_a21oi_1 _30013_ (.A1(_03896_),
    .A2(net7767),
    .Y(_02113_),
    .B1(_07439_));
 sg13g2_o21ai_1 _30014_ (.B1(net9395),
    .Y(_07440_),
    .A1(net4638),
    .A2(net7770));
 sg13g2_a21oi_1 _30015_ (.A1(_03904_),
    .A2(net7770),
    .Y(_02114_),
    .B1(_07440_));
 sg13g2_o21ai_1 _30016_ (.B1(net9370),
    .Y(_07441_),
    .A1(net4630),
    .A2(net7771));
 sg13g2_a21oi_1 _30017_ (.A1(_03921_),
    .A2(net7762),
    .Y(_02115_),
    .B1(_07441_));
 sg13g2_o21ai_1 _30018_ (.B1(net9352),
    .Y(_07442_),
    .A1(net4430),
    .A2(net7762));
 sg13g2_a21oi_1 _30019_ (.A1(_03927_),
    .A2(net7762),
    .Y(_02116_),
    .B1(_07442_));
 sg13g2_o21ai_1 _30020_ (.B1(net9346),
    .Y(_07443_),
    .A1(net4435),
    .A2(net7762));
 sg13g2_a21oi_1 _30021_ (.A1(_03933_),
    .A2(net7762),
    .Y(_02117_),
    .B1(_07443_));
 sg13g2_o21ai_1 _30022_ (.B1(net9355),
    .Y(_07444_),
    .A1(net4356),
    .A2(net7763));
 sg13g2_a21oi_1 _30023_ (.A1(_03952_),
    .A2(net7763),
    .Y(_02118_),
    .B1(_07444_));
 sg13g2_o21ai_1 _30024_ (.B1(net9357),
    .Y(_07445_),
    .A1(net4351),
    .A2(net7763));
 sg13g2_a21oi_1 _30025_ (.A1(_03958_),
    .A2(net7763),
    .Y(_02119_),
    .B1(_07445_));
 sg13g2_o21ai_1 _30026_ (.B1(net9354),
    .Y(_07446_),
    .A1(net4294),
    .A2(net7763));
 sg13g2_a21oi_1 _30027_ (.A1(_03964_),
    .A2(net7763),
    .Y(_02120_),
    .B1(_07446_));
 sg13g2_o21ai_1 _30028_ (.B1(net9357),
    .Y(_07447_),
    .A1(net4633),
    .A2(net7763));
 sg13g2_a21oi_1 _30029_ (.A1(_03971_),
    .A2(net7763),
    .Y(_02121_),
    .B1(_07447_));
 sg13g2_nor2_1 _30030_ (.A(net8350),
    .B(_04595_),
    .Y(_07448_));
 sg13g2_nand2_1 _30031_ (.Y(_07449_),
    .A(net5397),
    .B(net5266));
 sg13g2_o21ai_1 _30032_ (.B1(_07448_),
    .Y(_07450_),
    .A1(_04607_),
    .A2(_07449_));
 sg13g2_a21oi_1 _30033_ (.A1(_03979_),
    .A2(net8120),
    .Y(_07451_),
    .B1(_07450_));
 sg13g2_o21ai_1 _30034_ (.B1(net9350),
    .Y(_07452_),
    .A1(net5397),
    .A2(_07448_));
 sg13g2_nor2_1 _30035_ (.A(_07451_),
    .B(_07452_),
    .Y(_02122_));
 sg13g2_o21ai_1 _30036_ (.B1(net9358),
    .Y(_07453_),
    .A1(net4366),
    .A2(net7764));
 sg13g2_a21oi_1 _30037_ (.A1(_03987_),
    .A2(net7764),
    .Y(_02123_),
    .B1(_07453_));
 sg13g2_o21ai_1 _30038_ (.B1(net9359),
    .Y(_07454_),
    .A1(net4752),
    .A2(net7764));
 sg13g2_a21oi_1 _30039_ (.A1(_03995_),
    .A2(net7764),
    .Y(_02124_),
    .B1(_07454_));
 sg13g2_o21ai_1 _30040_ (.B1(net9367),
    .Y(_07455_),
    .A1(net4479),
    .A2(net7766));
 sg13g2_a21oi_1 _30041_ (.A1(_04002_),
    .A2(net7766),
    .Y(_02125_),
    .B1(_07455_));
 sg13g2_o21ai_1 _30042_ (.B1(net9401),
    .Y(_07456_),
    .A1(net4661),
    .A2(net7769));
 sg13g2_a21oi_1 _30043_ (.A1(_04008_),
    .A2(net7769),
    .Y(_02126_),
    .B1(_07456_));
 sg13g2_o21ai_1 _30044_ (.B1(net9400),
    .Y(_07457_),
    .A1(net4465),
    .A2(net7769));
 sg13g2_a21oi_1 _30045_ (.A1(_04014_),
    .A2(net7769),
    .Y(_02127_),
    .B1(_07457_));
 sg13g2_o21ai_1 _30046_ (.B1(net9388),
    .Y(_07458_),
    .A1(net4378),
    .A2(net7768));
 sg13g2_a21oi_1 _30047_ (.A1(_04020_),
    .A2(net7768),
    .Y(_02128_),
    .B1(_07458_));
 sg13g2_o21ai_1 _30048_ (.B1(net9388),
    .Y(_07459_),
    .A1(net4514),
    .A2(net7768));
 sg13g2_a21oi_1 _30049_ (.A1(_04027_),
    .A2(net7768),
    .Y(_02129_),
    .B1(_07459_));
 sg13g2_o21ai_1 _30050_ (.B1(net9388),
    .Y(_07460_),
    .A1(net4864),
    .A2(net7768));
 sg13g2_a21oi_1 _30051_ (.A1(_04033_),
    .A2(net7768),
    .Y(_02130_),
    .B1(_07460_));
 sg13g2_o21ai_1 _30052_ (.B1(net9402),
    .Y(_07461_),
    .A1(net5060),
    .A2(net7769));
 sg13g2_a21oi_1 _30053_ (.A1(_04039_),
    .A2(net7769),
    .Y(_02131_),
    .B1(_07461_));
 sg13g2_o21ai_1 _30054_ (.B1(net9383),
    .Y(_07462_),
    .A1(net4412),
    .A2(net7768));
 sg13g2_a21oi_1 _30055_ (.A1(_04045_),
    .A2(net7768),
    .Y(_02132_),
    .B1(_07462_));
 sg13g2_o21ai_1 _30056_ (.B1(net9384),
    .Y(_07463_),
    .A1(net4311),
    .A2(net7765));
 sg13g2_a21oi_1 _30057_ (.A1(_04052_),
    .A2(net7765),
    .Y(_02133_),
    .B1(_07463_));
 sg13g2_o21ai_1 _30058_ (.B1(net9383),
    .Y(_07464_),
    .A1(net4557),
    .A2(net7765));
 sg13g2_a21oi_1 _30059_ (.A1(_04058_),
    .A2(net7765),
    .Y(_02134_),
    .B1(_07464_));
 sg13g2_o21ai_1 _30060_ (.B1(net9364),
    .Y(_07465_),
    .A1(net4401),
    .A2(net7765));
 sg13g2_a21oi_1 _30061_ (.A1(_04064_),
    .A2(net7765),
    .Y(_02135_),
    .B1(_07465_));
 sg13g2_nand2_1 _30062_ (.Y(_07466_),
    .A(net8929),
    .B(_07042_));
 sg13g2_mux2_1 _30063_ (.A0(_07466_),
    .A1(net4117),
    .S(net7393),
    .X(_02136_));
 sg13g2_nor2_1 _30064_ (.A(net8938),
    .B(net7394),
    .Y(_07467_));
 sg13g2_o21ai_1 _30065_ (.B1(_07467_),
    .Y(_07468_),
    .A1(net4032),
    .A2(_06988_));
 sg13g2_o21ai_1 _30066_ (.B1(_07468_),
    .Y(_07469_),
    .A1(\soc_I.tx_uart_i.return_state[1] ),
    .A2(_07467_));
 sg13g2_inv_1 _30067_ (.Y(_02137_),
    .A(net4033));
 sg13g2_o21ai_1 _30068_ (.B1(net3927),
    .Y(_07470_),
    .A1(net8938),
    .A2(net7394));
 sg13g2_o21ai_1 _30069_ (.B1(_07470_),
    .Y(_02138_),
    .A1(net8933),
    .A2(_07468_));
 sg13g2_nand2_1 _30070_ (.Y(_07471_),
    .A(net3009),
    .B(_06847_));
 sg13g2_nand2_1 _30071_ (.Y(_07472_),
    .A(\soc_I.rx_uart_i.state[1] ),
    .B(\soc_I.rx_uart_i.state[0] ));
 sg13g2_nand2_1 _30072_ (.Y(_07473_),
    .A(net8798),
    .B(_07472_));
 sg13g2_o21ai_1 _30073_ (.B1(_07471_),
    .Y(_02139_),
    .A1(_06847_),
    .A2(_07473_));
 sg13g2_nand2_1 _30074_ (.Y(_07474_),
    .A(_06852_),
    .B(net8798));
 sg13g2_mux2_1 _30075_ (.A0(_07474_),
    .A1(net2611),
    .S(_06847_),
    .X(_02140_));
 sg13g2_nand2_1 _30076_ (.Y(_07475_),
    .A(net9411),
    .B(net9226));
 sg13g2_nor3_1 _30077_ (.A(net2601),
    .B(_05641_),
    .C(_07475_),
    .Y(_02141_));
 sg13g2_or2_1 _30078_ (.X(_07476_),
    .B(_05023_),
    .A(net2616));
 sg13g2_a221oi_1 _30079_ (.B2(_07476_),
    .C1(net9054),
    .B1(_05642_),
    .A1(_10592_),
    .Y(_02142_),
    .A2(net8943));
 sg13g2_nor4_1 _30080_ (.A(net9060),
    .B(net8984),
    .C(net9718),
    .D(_05750_),
    .Y(_02143_));
 sg13g2_nor2b_1 _30081_ (.A(_05646_),
    .B_N(_05751_),
    .Y(_07477_));
 sg13g2_nor2_1 _30082_ (.A(net9060),
    .B(_07477_),
    .Y(_02144_));
 sg13g2_nand2b_1 _30083_ (.Y(_07478_),
    .B(net9078),
    .A_N(_05733_));
 sg13g2_nand3_1 _30084_ (.B(_05731_),
    .C(_07478_),
    .A(net9001),
    .Y(_07479_));
 sg13g2_nand2_1 _30085_ (.Y(_07480_),
    .A(_10993_),
    .B(net8328));
 sg13g2_o21ai_1 _30086_ (.B1(_07480_),
    .Y(_07481_),
    .A1(net7975),
    .A2(net8328));
 sg13g2_a21o_1 _30087_ (.A2(_07481_),
    .A1(net9217),
    .B1(_07479_),
    .X(_07482_));
 sg13g2_inv_2 _30088_ (.Y(_07483_),
    .A(net7755));
 sg13g2_nor2b_1 _30089_ (.A(net9769),
    .B_N(net9758),
    .Y(_07484_));
 sg13g2_mux4_1 _30090_ (.S0(net9769),
    .A0(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[0] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[1] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[2] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[3] ),
    .S1(net9758),
    .X(_07485_));
 sg13g2_a21oi_1 _30091_ (.A1(net9769),
    .A2(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[5] ),
    .Y(_07486_),
    .B1(net9758));
 sg13g2_o21ai_1 _30092_ (.B1(_07486_),
    .Y(_07487_),
    .A1(net9769),
    .A2(_10608_));
 sg13g2_a221oi_1 _30093_ (.B2(_10609_),
    .C1(net9070),
    .B1(_07484_),
    .A1(_10610_),
    .Y(_07488_),
    .A2(_05739_));
 sg13g2_a21o_1 _30094_ (.A2(_07485_),
    .A1(net9070),
    .B1(net9740),
    .X(_07489_));
 sg13g2_a21o_1 _30095_ (.A2(_07488_),
    .A1(_07487_),
    .B1(_07489_),
    .X(_07490_));
 sg13g2_mux4_1 _30096_ (.S0(net9768),
    .A0(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[12] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[13] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[14] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[15] ),
    .S1(net9752),
    .X(_07491_));
 sg13g2_nor2_1 _30097_ (.A(_05749_),
    .B(_07491_),
    .Y(_07492_));
 sg13g2_mux4_1 _30098_ (.S0(net9768),
    .A0(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[8] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[9] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[10] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[11] ),
    .S1(net9752),
    .X(_07493_));
 sg13g2_nand2b_1 _30099_ (.Y(_07494_),
    .B(net9740),
    .A_N(net9744));
 sg13g2_o21ai_1 _30100_ (.B1(net9076),
    .Y(_07495_),
    .A1(_07493_),
    .A2(_07494_));
 sg13g2_nor2_1 _30101_ (.A(_07492_),
    .B(_07495_),
    .Y(_07496_));
 sg13g2_nand2_1 _30102_ (.Y(_07497_),
    .A(_07490_),
    .B(_07496_));
 sg13g2_a21oi_1 _30103_ (.A1(net9769),
    .A2(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[21] ),
    .Y(_07498_),
    .B1(net9758));
 sg13g2_o21ai_1 _30104_ (.B1(_07498_),
    .Y(_07499_),
    .A1(net9769),
    .A2(_10614_));
 sg13g2_a221oi_1 _30105_ (.B2(_10615_),
    .C1(net9070),
    .B1(_07484_),
    .A1(_10616_),
    .Y(_07500_),
    .A2(_05739_));
 sg13g2_mux4_1 _30106_ (.S0(net9769),
    .A0(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[16] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[17] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[18] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[19] ),
    .S1(net9758),
    .X(_07501_));
 sg13g2_a21o_1 _30107_ (.A2(_07501_),
    .A1(net9070),
    .B1(net9740),
    .X(_07502_));
 sg13g2_a21o_1 _30108_ (.A2(_07500_),
    .A1(_07499_),
    .B1(_07502_),
    .X(_07503_));
 sg13g2_mux4_1 _30109_ (.S0(net9767),
    .A0(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[24] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[25] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[26] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[27] ),
    .S1(net9757),
    .X(_07504_));
 sg13g2_nor2_1 _30110_ (.A(_07494_),
    .B(_07504_),
    .Y(_07505_));
 sg13g2_mux4_1 _30111_ (.S0(net9769),
    .A0(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[28] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[29] ),
    .A2(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[30] ),
    .A3(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[31] ),
    .S1(net9758),
    .X(_07506_));
 sg13g2_o21ai_1 _30112_ (.B1(net9719),
    .Y(_07507_),
    .A1(_05749_),
    .A2(_07506_));
 sg13g2_nor2_1 _30113_ (.A(_07505_),
    .B(_07507_),
    .Y(_07508_));
 sg13g2_nand2_1 _30114_ (.Y(_07509_),
    .A(_07503_),
    .B(_07508_));
 sg13g2_a22oi_1 _30115_ (.Y(_07510_),
    .B1(_07503_),
    .B2(_07508_),
    .A2(_07496_),
    .A1(_07490_));
 sg13g2_nand2_1 _30116_ (.Y(_07511_),
    .A(_07497_),
    .B(_07509_));
 sg13g2_nand3_1 _30117_ (.B(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[31] ),
    .C(net8533),
    .A(net9766),
    .Y(_07512_));
 sg13g2_nor2_1 _30118_ (.A(_00256_),
    .B(_07512_),
    .Y(_07513_));
 sg13g2_nand2b_1 _30119_ (.Y(_07514_),
    .B(_07513_),
    .A_N(_00255_));
 sg13g2_nor2_2 _30120_ (.A(net9731),
    .B(_07514_),
    .Y(_07515_));
 sg13g2_nand3_1 _30121_ (.B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[62] ),
    .C(_07515_),
    .A(net9724),
    .Y(_07516_));
 sg13g2_nand2_1 _30122_ (.Y(_07517_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[29] ),
    .B(net8532));
 sg13g2_nand2_1 _30123_ (.Y(_07518_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[28] ),
    .B(net8534));
 sg13g2_mux2_1 _30124_ (.A0(_07517_),
    .A1(_07518_),
    .S(net9766),
    .X(_07519_));
 sg13g2_nand2_1 _30125_ (.Y(_07520_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[30] ),
    .B(net8533));
 sg13g2_a21oi_1 _30126_ (.A1(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[31] ),
    .A2(net8533),
    .Y(_07521_),
    .B1(net9764));
 sg13g2_a21o_1 _30127_ (.A2(_07520_),
    .A1(net9767),
    .B1(_07521_),
    .X(_07522_));
 sg13g2_mux2_1 _30128_ (.A0(_07519_),
    .A1(_07522_),
    .S(net9065),
    .X(_07523_));
 sg13g2_nor2_1 _30129_ (.A(_00255_),
    .B(_07523_),
    .Y(_07524_));
 sg13g2_nor3_2 _30130_ (.A(_00255_),
    .B(net9732),
    .C(_07523_),
    .Y(_07525_));
 sg13g2_and2_1 _30131_ (.A(net9724),
    .B(_07525_),
    .X(_07526_));
 sg13g2_and2_1 _30132_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[59] ),
    .B(_07526_),
    .X(_07527_));
 sg13g2_xor2_1 _30133_ (.B(_07526_),
    .A(_00280_),
    .X(_07528_));
 sg13g2_nor2_1 _30134_ (.A(_00256_),
    .B(_07522_),
    .Y(_07529_));
 sg13g2_nand2_1 _30135_ (.Y(_07530_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[27] ),
    .B(net8534));
 sg13g2_nand2_1 _30136_ (.Y(_07531_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[26] ),
    .B(net8533));
 sg13g2_mux2_1 _30137_ (.A0(_07530_),
    .A1(_07531_),
    .S(net9766),
    .X(_07532_));
 sg13g2_mux2_1 _30138_ (.A0(_07519_),
    .A1(_07532_),
    .S(net9755),
    .X(_07533_));
 sg13g2_nor2_1 _30139_ (.A(net9068),
    .B(_07533_),
    .Y(_07534_));
 sg13g2_a21oi_1 _30140_ (.A1(net9070),
    .A2(_07529_),
    .Y(_07535_),
    .B1(_07534_));
 sg13g2_nor2_2 _30141_ (.A(net9732),
    .B(_07535_),
    .Y(_07536_));
 sg13g2_nand2_1 _30142_ (.Y(_07537_),
    .A(net9724),
    .B(_07536_));
 sg13g2_nand2_1 _30143_ (.Y(_07538_),
    .A(_00278_),
    .B(_07537_));
 sg13g2_nor2_1 _30144_ (.A(_00278_),
    .B(_07537_),
    .Y(_07539_));
 sg13g2_mux2_1 _30145_ (.A0(_07520_),
    .A1(_07517_),
    .S(net9767),
    .X(_07540_));
 sg13g2_mux2_2 _30146_ (.A0(_07512_),
    .A1(_07540_),
    .S(net9754),
    .X(_07541_));
 sg13g2_nand2_1 _30147_ (.Y(_07542_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[25] ),
    .B(net8532));
 sg13g2_nand3_1 _30148_ (.B(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[25] ),
    .C(net8533),
    .A(net9764),
    .Y(_07543_));
 sg13g2_o21ai_1 _30149_ (.B1(_07543_),
    .Y(_07544_),
    .A1(net9766),
    .A2(_07531_));
 sg13g2_mux2_1 _30150_ (.A0(_07518_),
    .A1(_07530_),
    .S(net9766),
    .X(_07545_));
 sg13g2_nand2_1 _30151_ (.Y(_07546_),
    .A(net9065),
    .B(_07545_));
 sg13g2_o21ai_1 _30152_ (.B1(_07546_),
    .Y(_07547_),
    .A1(net9065),
    .A2(_07544_));
 sg13g2_mux2_2 _30153_ (.A0(_07541_),
    .A1(_07547_),
    .S(net9749),
    .X(_07548_));
 sg13g2_nor2_1 _30154_ (.A(net9731),
    .B(_07548_),
    .Y(_07549_));
 sg13g2_nor3_2 _30155_ (.A(net9076),
    .B(net9731),
    .C(_07548_),
    .Y(_07550_));
 sg13g2_xor2_1 _30156_ (.B(_07550_),
    .A(_00277_),
    .X(_07551_));
 sg13g2_nor2_1 _30157_ (.A(net9745),
    .B(_07523_),
    .Y(_07552_));
 sg13g2_nand3_1 _30158_ (.B(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[24] ),
    .C(net8532),
    .A(net9768),
    .Y(_07553_));
 sg13g2_o21ai_1 _30159_ (.B1(_07553_),
    .Y(_07554_),
    .A1(net9765),
    .A2(_07542_));
 sg13g2_nor2_1 _30160_ (.A(_10512_),
    .B(_07554_),
    .Y(_07555_));
 sg13g2_a21oi_1 _30161_ (.A1(net9065),
    .A2(_07532_),
    .Y(_07556_),
    .B1(_07555_));
 sg13g2_a21oi_2 _30162_ (.B1(_07552_),
    .Y(_07557_),
    .A2(_07556_),
    .A1(net9745));
 sg13g2_nor2_2 _30163_ (.A(net9731),
    .B(_07557_),
    .Y(_07558_));
 sg13g2_nand2_1 _30164_ (.Y(_07559_),
    .A(net9725),
    .B(_07558_));
 sg13g2_or2_1 _30165_ (.X(_07560_),
    .B(_07559_),
    .A(_00276_));
 sg13g2_nand2_1 _30166_ (.Y(_07561_),
    .A(_00276_),
    .B(_07559_));
 sg13g2_mux2_1 _30167_ (.A0(_07540_),
    .A1(_07545_),
    .S(net9755),
    .X(_07562_));
 sg13g2_nand2_1 _30168_ (.Y(_07563_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[23] ),
    .B(net8533));
 sg13g2_a21oi_1 _30169_ (.A1(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[24] ),
    .A2(net8532),
    .Y(_07564_),
    .B1(net9768));
 sg13g2_a21oi_1 _30170_ (.A1(net9765),
    .A2(_07563_),
    .Y(_07565_),
    .B1(_07564_));
 sg13g2_and2_1 _30171_ (.A(net9754),
    .B(_07565_),
    .X(_07566_));
 sg13g2_a21oi_1 _30172_ (.A1(net9065),
    .A2(_07544_),
    .Y(_07567_),
    .B1(_07566_));
 sg13g2_and2_1 _30173_ (.A(net9069),
    .B(_07562_),
    .X(_07568_));
 sg13g2_a21oi_1 _30174_ (.A1(net9746),
    .A2(_07567_),
    .Y(_07569_),
    .B1(_07568_));
 sg13g2_nand2_1 _30175_ (.Y(_07570_),
    .A(net9737),
    .B(_07569_));
 sg13g2_o21ai_1 _30176_ (.B1(_07570_),
    .Y(_07571_),
    .A1(net9737),
    .A2(_07514_));
 sg13g2_nand2_1 _30177_ (.Y(_07572_),
    .A(net9724),
    .B(_07571_));
 sg13g2_nand3_1 _30178_ (.B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[54] ),
    .C(_07571_),
    .A(net9724),
    .Y(_07573_));
 sg13g2_xor2_1 _30179_ (.B(_07572_),
    .A(_00275_),
    .X(_07574_));
 sg13g2_inv_1 _30180_ (.Y(_07575_),
    .A(_07574_));
 sg13g2_nand2b_1 _30181_ (.Y(_07576_),
    .B(_07529_),
    .A_N(_00255_));
 sg13g2_nand2_1 _30182_ (.Y(_07577_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[22] ),
    .B(net8533));
 sg13g2_mux2_1 _30183_ (.A0(_07563_),
    .A1(_07577_),
    .S(net9765),
    .X(_07578_));
 sg13g2_nor2_1 _30184_ (.A(net9754),
    .B(_07554_),
    .Y(_07579_));
 sg13g2_a21oi_1 _30185_ (.A1(net9754),
    .A2(_07578_),
    .Y(_07580_),
    .B1(_07579_));
 sg13g2_nand2_1 _30186_ (.Y(_07581_),
    .A(net9746),
    .B(_07580_));
 sg13g2_o21ai_1 _30187_ (.B1(_07581_),
    .Y(_07582_),
    .A1(net9745),
    .A2(_07533_));
 sg13g2_nand2_1 _30188_ (.Y(_07583_),
    .A(net9737),
    .B(_07582_));
 sg13g2_o21ai_1 _30189_ (.B1(_07583_),
    .Y(_07584_),
    .A1(net9738),
    .A2(_07576_));
 sg13g2_nand2_1 _30190_ (.Y(_07585_),
    .A(net9725),
    .B(_07584_));
 sg13g2_nor2_1 _30191_ (.A(_00274_),
    .B(_07585_),
    .Y(_07586_));
 sg13g2_nand2_1 _30192_ (.Y(_07587_),
    .A(_00274_),
    .B(_07585_));
 sg13g2_or3_1 _30193_ (.A(net9740),
    .B(_00255_),
    .C(_07541_),
    .X(_07588_));
 sg13g2_nor2_1 _30194_ (.A(net9749),
    .B(_07547_),
    .Y(_07589_));
 sg13g2_nand2_1 _30195_ (.Y(_07590_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[21] ),
    .B(net8534));
 sg13g2_nand3_1 _30196_ (.B(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[21] ),
    .C(net8534),
    .A(net9765),
    .Y(_07591_));
 sg13g2_o21ai_1 _30197_ (.B1(_07591_),
    .Y(_07592_),
    .A1(net9764),
    .A2(_07577_));
 sg13g2_mux2_1 _30198_ (.A0(_07565_),
    .A1(_07592_),
    .S(net9757),
    .X(_07593_));
 sg13g2_a21oi_1 _30199_ (.A1(net9745),
    .A2(_07593_),
    .Y(_07594_),
    .B1(_07589_));
 sg13g2_o21ai_1 _30200_ (.B1(_07588_),
    .Y(_07595_),
    .A1(net9072),
    .A2(_07594_));
 sg13g2_and2_1 _30201_ (.A(net9726),
    .B(_07595_),
    .X(_07596_));
 sg13g2_nand2_1 _30202_ (.Y(_07597_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[52] ),
    .B(_07596_));
 sg13g2_nand2_1 _30203_ (.Y(_07598_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[20] ),
    .B(net8532));
 sg13g2_mux2_1 _30204_ (.A0(_07590_),
    .A1(_07598_),
    .S(net9765),
    .X(_07599_));
 sg13g2_and2_1 _30205_ (.A(net9754),
    .B(_07599_),
    .X(_07600_));
 sg13g2_a21oi_1 _30206_ (.A1(_10512_),
    .A2(_07578_),
    .Y(_07601_),
    .B1(_07600_));
 sg13g2_mux2_1 _30207_ (.A0(_07556_),
    .A1(_07601_),
    .S(net9745),
    .X(_07602_));
 sg13g2_mux2_2 _30208_ (.A0(_07524_),
    .A1(_07602_),
    .S(net9737),
    .X(_07603_));
 sg13g2_a21oi_1 _30209_ (.A1(net9726),
    .A2(_07603_),
    .Y(_07604_),
    .B1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[51] ));
 sg13g2_nand3_1 _30210_ (.B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[51] ),
    .C(_07603_),
    .A(net9726),
    .Y(_07605_));
 sg13g2_nand2_1 _30211_ (.Y(_07606_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[19] ),
    .B(net8532));
 sg13g2_mux2_1 _30212_ (.A0(_07598_),
    .A1(_07606_),
    .S(net9764),
    .X(_07607_));
 sg13g2_nand2_1 _30213_ (.Y(_07608_),
    .A(net9754),
    .B(_07607_));
 sg13g2_o21ai_1 _30214_ (.B1(_07608_),
    .Y(_07609_),
    .A1(net9754),
    .A2(_07592_));
 sg13g2_or2_1 _30215_ (.X(_07610_),
    .B(_07609_),
    .A(net9068));
 sg13g2_o21ai_1 _30216_ (.B1(_07610_),
    .Y(_07611_),
    .A1(net9745),
    .A2(_07567_));
 sg13g2_nor2_1 _30217_ (.A(net9746),
    .B(_07513_),
    .Y(_07612_));
 sg13g2_a21oi_1 _30218_ (.A1(net9745),
    .A2(_07562_),
    .Y(_07613_),
    .B1(_07612_));
 sg13g2_mux2_2 _30219_ (.A0(_07611_),
    .A1(_07613_),
    .S(net9072),
    .X(_07614_));
 sg13g2_nand2_1 _30220_ (.Y(_07615_),
    .A(net9728),
    .B(_07614_));
 sg13g2_nand3_1 _30221_ (.B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[50] ),
    .C(_07614_),
    .A(net9728),
    .Y(_07616_));
 sg13g2_nand2_1 _30222_ (.Y(_07617_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[18] ),
    .B(net8532));
 sg13g2_mux2_1 _30223_ (.A0(_07606_),
    .A1(_07617_),
    .S(net9764),
    .X(_07618_));
 sg13g2_mux2_1 _30224_ (.A0(_07599_),
    .A1(_07618_),
    .S(net9754),
    .X(_07619_));
 sg13g2_nor2_1 _30225_ (.A(net9745),
    .B(_07580_),
    .Y(_07620_));
 sg13g2_a21oi_2 _30226_ (.B1(_07620_),
    .Y(_07621_),
    .A2(_07619_),
    .A1(net9746));
 sg13g2_nor2_1 _30227_ (.A(net9738),
    .B(_07535_),
    .Y(_07622_));
 sg13g2_a21oi_2 _30228_ (.B1(_07622_),
    .Y(_07623_),
    .A2(_07621_),
    .A1(net9739));
 sg13g2_nor3_1 _30229_ (.A(net9075),
    .B(_00271_),
    .C(_07623_),
    .Y(_07624_));
 sg13g2_o21ai_1 _30230_ (.B1(_00271_),
    .Y(_07625_),
    .A1(net9076),
    .A2(_07623_));
 sg13g2_nand2_1 _30231_ (.Y(_07626_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[16] ),
    .B(net8532));
 sg13g2_a21oi_1 _30232_ (.A1(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[17] ),
    .A2(net8535),
    .Y(_07627_),
    .B1(net9764));
 sg13g2_a21oi_1 _30233_ (.A1(net9766),
    .A2(_07626_),
    .Y(_07628_),
    .B1(_07627_));
 sg13g2_nand2_1 _30234_ (.Y(_07629_),
    .A(net9065),
    .B(_07618_));
 sg13g2_o21ai_1 _30235_ (.B1(_07629_),
    .Y(_07630_),
    .A1(net9065),
    .A2(_07628_));
 sg13g2_nor2_1 _30236_ (.A(net9747),
    .B(_07601_),
    .Y(_07631_));
 sg13g2_a21oi_1 _30237_ (.A1(net9747),
    .A2(_07630_),
    .Y(_07632_),
    .B1(_07631_));
 sg13g2_nor2_1 _30238_ (.A(net9072),
    .B(_07632_),
    .Y(_07633_));
 sg13g2_a21oi_2 _30239_ (.B1(_07633_),
    .Y(_07634_),
    .A2(_07557_),
    .A1(net9072));
 sg13g2_a21oi_1 _30240_ (.A1(net9729),
    .A2(_07634_),
    .Y(_07635_),
    .B1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[47] ));
 sg13g2_nand3_1 _30241_ (.B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[47] ),
    .C(_07634_),
    .A(net9729),
    .Y(_07636_));
 sg13g2_nand2b_1 _30242_ (.Y(_07637_),
    .B(_07636_),
    .A_N(_07635_));
 sg13g2_nor2_1 _30243_ (.A(net9749),
    .B(_07609_),
    .Y(_07638_));
 sg13g2_nand2_1 _30244_ (.Y(_07639_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[15] ),
    .B(net8535));
 sg13g2_mux2_1 _30245_ (.A0(_07626_),
    .A1(_07639_),
    .S(net9767),
    .X(_07640_));
 sg13g2_nand3_1 _30246_ (.B(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[17] ),
    .C(net8535),
    .A(net9764),
    .Y(_07641_));
 sg13g2_o21ai_1 _30247_ (.B1(_07641_),
    .Y(_07642_),
    .A1(net9764),
    .A2(_07617_));
 sg13g2_nor2_1 _30248_ (.A(net9755),
    .B(_07642_),
    .Y(_07643_));
 sg13g2_a21oi_1 _30249_ (.A1(net9756),
    .A2(_07640_),
    .Y(_07644_),
    .B1(_07643_));
 sg13g2_a21oi_2 _30250_ (.B1(_07638_),
    .Y(_07645_),
    .A2(_07644_),
    .A1(net9747));
 sg13g2_nand2_1 _30251_ (.Y(_07646_),
    .A(net9737),
    .B(_07645_));
 sg13g2_o21ai_1 _30252_ (.B1(_07646_),
    .Y(_07647_),
    .A1(net9737),
    .A2(_07569_));
 sg13g2_nor2_1 _30253_ (.A(net9727),
    .B(_07515_),
    .Y(_07648_));
 sg13g2_a21oi_2 _30254_ (.B1(_07648_),
    .Y(_07649_),
    .A2(_07647_),
    .A1(net9727));
 sg13g2_nand2_1 _30255_ (.Y(_07650_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[46] ),
    .B(_07649_));
 sg13g2_xor2_1 _30256_ (.B(_07649_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[46] ),
    .X(_07651_));
 sg13g2_inv_1 _30257_ (.Y(_07652_),
    .A(_07651_));
 sg13g2_nor2_1 _30258_ (.A(_07637_),
    .B(_07652_),
    .Y(_07653_));
 sg13g2_nor2_1 _30259_ (.A(net9731),
    .B(_07576_),
    .Y(_07654_));
 sg13g2_nand2_1 _30260_ (.Y(_07655_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[14] ),
    .B(net8536));
 sg13g2_mux2_1 _30261_ (.A0(_07639_),
    .A1(_07655_),
    .S(net9767),
    .X(_07656_));
 sg13g2_nor2_1 _30262_ (.A(net9755),
    .B(_07628_),
    .Y(_07657_));
 sg13g2_a21oi_2 _30263_ (.B1(_07657_),
    .Y(_07658_),
    .A2(_07656_),
    .A1(net9753));
 sg13g2_nand2_1 _30264_ (.Y(_07659_),
    .A(net9748),
    .B(_07658_));
 sg13g2_o21ai_1 _30265_ (.B1(_07659_),
    .Y(_07660_),
    .A1(net9747),
    .A2(_07619_));
 sg13g2_mux2_1 _30266_ (.A0(_07582_),
    .A1(_07660_),
    .S(net9738),
    .X(_07661_));
 sg13g2_mux2_1 _30267_ (.A0(_07654_),
    .A1(_07661_),
    .S(net9727),
    .X(_07662_));
 sg13g2_nor2_1 _30268_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[45] ),
    .B(_07662_),
    .Y(_07663_));
 sg13g2_inv_1 _30269_ (.Y(_07664_),
    .A(_07663_));
 sg13g2_nand2_1 _30270_ (.Y(_07665_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[45] ),
    .B(_07662_));
 sg13g2_nor3_2 _30271_ (.A(_00255_),
    .B(net9731),
    .C(_07541_),
    .Y(_07666_));
 sg13g2_nand2_1 _30272_ (.Y(_07667_),
    .A(_10512_),
    .B(_07607_));
 sg13g2_o21ai_1 _30273_ (.B1(_07667_),
    .Y(_07668_),
    .A1(net9065),
    .A2(_07642_));
 sg13g2_nand2_1 _30274_ (.Y(_07669_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[13] ),
    .B(net8536));
 sg13g2_mux2_1 _30275_ (.A0(_07655_),
    .A1(_07669_),
    .S(net9767),
    .X(_07670_));
 sg13g2_mux2_1 _30276_ (.A0(_07640_),
    .A1(_07670_),
    .S(net9753),
    .X(_07671_));
 sg13g2_or2_1 _30277_ (.X(_07672_),
    .B(_07671_),
    .A(net9067));
 sg13g2_o21ai_1 _30278_ (.B1(_07672_),
    .Y(_07673_),
    .A1(net9747),
    .A2(_07668_));
 sg13g2_nor2_1 _30279_ (.A(net9737),
    .B(_07594_),
    .Y(_07674_));
 sg13g2_a21oi_2 _30280_ (.B1(_07674_),
    .Y(_07675_),
    .A2(_07673_),
    .A1(net9737));
 sg13g2_nor2_1 _30281_ (.A(net9727),
    .B(_07666_),
    .Y(_07676_));
 sg13g2_a21oi_2 _30282_ (.B1(_07676_),
    .Y(_07677_),
    .A2(_07675_),
    .A1(net9720));
 sg13g2_nand2_1 _30283_ (.Y(_07678_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[44] ),
    .B(_07677_));
 sg13g2_nand2_1 _30284_ (.Y(_07679_),
    .A(_07665_),
    .B(_07678_));
 sg13g2_nand2_1 _30285_ (.Y(_07680_),
    .A(_07664_),
    .B(_07679_));
 sg13g2_nor2b_1 _30286_ (.A(_07663_),
    .B_N(_07665_),
    .Y(_07681_));
 sg13g2_xor2_1 _30287_ (.B(_07677_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[44] ),
    .X(_07682_));
 sg13g2_nand2_1 _30288_ (.Y(_07683_),
    .A(_07681_),
    .B(_07682_));
 sg13g2_nor2_1 _30289_ (.A(net9748),
    .B(_07630_),
    .Y(_07684_));
 sg13g2_nand2_1 _30290_ (.Y(_07685_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[12] ),
    .B(net8531));
 sg13g2_mux2_1 _30291_ (.A0(_07669_),
    .A1(_07685_),
    .S(net9762),
    .X(_07686_));
 sg13g2_and2_1 _30292_ (.A(net9753),
    .B(_07686_),
    .X(_07687_));
 sg13g2_a21oi_1 _30293_ (.A1(net9066),
    .A2(_07656_),
    .Y(_07688_),
    .B1(_07687_));
 sg13g2_a21oi_1 _30294_ (.A1(net9748),
    .A2(_07688_),
    .Y(_07689_),
    .B1(_07684_));
 sg13g2_nand2_1 _30295_ (.Y(_07690_),
    .A(net9735),
    .B(_07689_));
 sg13g2_o21ai_1 _30296_ (.B1(_07690_),
    .Y(_07691_),
    .A1(net9738),
    .A2(_07602_));
 sg13g2_nor2_1 _30297_ (.A(net9726),
    .B(_07525_),
    .Y(_07692_));
 sg13g2_a21oi_2 _30298_ (.B1(_07692_),
    .Y(_07693_),
    .A2(_07691_),
    .A1(net9727));
 sg13g2_nor2_1 _30299_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[43] ),
    .B(_07693_),
    .Y(_07694_));
 sg13g2_nor2b_2 _30300_ (.A(net9731),
    .B_N(_07613_),
    .Y(_07695_));
 sg13g2_and2_1 _30301_ (.A(net9067),
    .B(_07644_),
    .X(_07696_));
 sg13g2_nand3_1 _30302_ (.B(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[11] ),
    .C(net8531),
    .A(net9763),
    .Y(_07697_));
 sg13g2_o21ai_1 _30303_ (.B1(_07697_),
    .Y(_07698_),
    .A1(net9762),
    .A2(_07685_));
 sg13g2_nand2_1 _30304_ (.Y(_07699_),
    .A(net9753),
    .B(_07698_));
 sg13g2_o21ai_1 _30305_ (.B1(_07699_),
    .Y(_07700_),
    .A1(net9753),
    .A2(_07670_));
 sg13g2_a21oi_2 _30306_ (.B1(_07696_),
    .Y(_07701_),
    .A2(_07700_),
    .A1(net9748));
 sg13g2_nand2_1 _30307_ (.Y(_07702_),
    .A(net9736),
    .B(_07701_));
 sg13g2_o21ai_1 _30308_ (.B1(_07702_),
    .Y(_07703_),
    .A1(net9738),
    .A2(_07611_));
 sg13g2_nor2_1 _30309_ (.A(net9726),
    .B(_07695_),
    .Y(_07704_));
 sg13g2_a21oi_2 _30310_ (.B1(_07704_),
    .Y(_07705_),
    .A2(_07703_),
    .A1(net9721));
 sg13g2_nand2_1 _30311_ (.Y(_07706_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[42] ),
    .B(_07705_));
 sg13g2_nand2_1 _30312_ (.Y(_07707_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[43] ),
    .B(_07693_));
 sg13g2_and2_1 _30313_ (.A(_07706_),
    .B(_07707_),
    .X(_07708_));
 sg13g2_nor2_1 _30314_ (.A(_07694_),
    .B(_07708_),
    .Y(_07709_));
 sg13g2_xor2_1 _30315_ (.B(_07705_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[42] ),
    .X(_07710_));
 sg13g2_nor2b_1 _30316_ (.A(_07694_),
    .B_N(_07707_),
    .Y(_07711_));
 sg13g2_and2_1 _30317_ (.A(_07710_),
    .B(_07711_),
    .X(_07712_));
 sg13g2_nand2_1 _30318_ (.Y(_07713_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[10] ),
    .B(net8531));
 sg13g2_a21oi_1 _30319_ (.A1(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[11] ),
    .A2(net8531),
    .Y(_07714_),
    .B1(net9763));
 sg13g2_a21oi_1 _30320_ (.A1(net9761),
    .A2(_07713_),
    .Y(_07715_),
    .B1(_07714_));
 sg13g2_nor2_1 _30321_ (.A(net9753),
    .B(_07686_),
    .Y(_07716_));
 sg13g2_a21oi_1 _30322_ (.A1(net9750),
    .A2(_07715_),
    .Y(_07717_),
    .B1(_07716_));
 sg13g2_nor2_1 _30323_ (.A(net9067),
    .B(_07717_),
    .Y(_07718_));
 sg13g2_a21oi_2 _30324_ (.B1(_07718_),
    .Y(_07719_),
    .A2(_07658_),
    .A1(net9068));
 sg13g2_nor2_1 _30325_ (.A(net9738),
    .B(_07621_),
    .Y(_07720_));
 sg13g2_a21oi_1 _30326_ (.A1(net9738),
    .A2(_07719_),
    .Y(_07721_),
    .B1(_07720_));
 sg13g2_mux2_1 _30327_ (.A0(_07536_),
    .A1(_07721_),
    .S(net9727),
    .X(_07722_));
 sg13g2_nor2_1 _30328_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[41] ),
    .B(_07722_),
    .Y(_07723_));
 sg13g2_nand2_1 _30329_ (.Y(_07724_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[41] ),
    .B(_07722_));
 sg13g2_nor2_1 _30330_ (.A(net9748),
    .B(_07671_),
    .Y(_07725_));
 sg13g2_nand2_1 _30331_ (.Y(_07726_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[9] ),
    .B(net8531));
 sg13g2_mux2_1 _30332_ (.A0(_07713_),
    .A1(_07726_),
    .S(net9761),
    .X(_07727_));
 sg13g2_nor2_1 _30333_ (.A(net9753),
    .B(_07698_),
    .Y(_07728_));
 sg13g2_a21oi_1 _30334_ (.A1(net9753),
    .A2(_07727_),
    .Y(_07729_),
    .B1(_07728_));
 sg13g2_a21oi_1 _30335_ (.A1(net9748),
    .A2(_07729_),
    .Y(_07730_),
    .B1(_07725_));
 sg13g2_nand2_1 _30336_ (.Y(_07731_),
    .A(net9068),
    .B(_07593_));
 sg13g2_o21ai_1 _30337_ (.B1(_07731_),
    .Y(_07732_),
    .A1(net9068),
    .A2(_07668_));
 sg13g2_nor2_1 _30338_ (.A(net9739),
    .B(_07732_),
    .Y(_07733_));
 sg13g2_a21oi_1 _30339_ (.A1(net9736),
    .A2(_07730_),
    .Y(_07734_),
    .B1(_07733_));
 sg13g2_mux2_1 _30340_ (.A0(_07549_),
    .A1(_07734_),
    .S(net9720),
    .X(_07735_));
 sg13g2_and2_1 _30341_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[40] ),
    .B(_07735_),
    .X(_07736_));
 sg13g2_inv_1 _30342_ (.Y(_07737_),
    .A(_07736_));
 sg13g2_o21ai_1 _30343_ (.B1(_07724_),
    .Y(_07738_),
    .A1(_07723_),
    .A2(_07737_));
 sg13g2_a21oi_1 _30344_ (.A1(_07712_),
    .A2(_07738_),
    .Y(_07739_),
    .B1(_07709_));
 sg13g2_o21ai_1 _30345_ (.B1(_07680_),
    .Y(_07740_),
    .A1(_07683_),
    .A2(_07739_));
 sg13g2_o21ai_1 _30346_ (.B1(_07636_),
    .Y(_07741_),
    .A1(_07635_),
    .A2(_07650_));
 sg13g2_nor3_1 _30347_ (.A(_07637_),
    .B(_07652_),
    .C(_07683_),
    .Y(_07742_));
 sg13g2_nor2b_1 _30348_ (.A(_07723_),
    .B_N(_07724_),
    .Y(_07743_));
 sg13g2_and2_1 _30349_ (.A(net9067),
    .B(_07688_),
    .X(_07744_));
 sg13g2_nand2_1 _30350_ (.Y(_07745_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[8] ),
    .B(net8531));
 sg13g2_mux2_1 _30351_ (.A0(_07726_),
    .A1(_07745_),
    .S(net9761),
    .X(_07746_));
 sg13g2_nor2_1 _30352_ (.A(net9750),
    .B(_07715_),
    .Y(_07747_));
 sg13g2_a21oi_1 _30353_ (.A1(net9750),
    .A2(_07746_),
    .Y(_07748_),
    .B1(_07747_));
 sg13g2_a21oi_1 _30354_ (.A1(net9741),
    .A2(_07748_),
    .Y(_07749_),
    .B1(_07744_));
 sg13g2_nor2_1 _30355_ (.A(net9735),
    .B(_07632_),
    .Y(_07750_));
 sg13g2_a21oi_1 _30356_ (.A1(net9735),
    .A2(_07749_),
    .Y(_07751_),
    .B1(_07750_));
 sg13g2_mux2_2 _30357_ (.A0(_07558_),
    .A1(_07751_),
    .S(net9723),
    .X(_07752_));
 sg13g2_nor2_1 _30358_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[39] ),
    .B(_07752_),
    .Y(_07753_));
 sg13g2_nand2_1 _30359_ (.Y(_07754_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[7] ),
    .B(net8531));
 sg13g2_mux2_1 _30360_ (.A0(_07745_),
    .A1(_07754_),
    .S(net9761),
    .X(_07755_));
 sg13g2_mux2_1 _30361_ (.A0(_07727_),
    .A1(_07755_),
    .S(net9750),
    .X(_07756_));
 sg13g2_nor2_1 _30362_ (.A(net9067),
    .B(_07756_),
    .Y(_07757_));
 sg13g2_a21oi_2 _30363_ (.B1(_07757_),
    .Y(_07758_),
    .A2(_07700_),
    .A1(net9067));
 sg13g2_mux2_1 _30364_ (.A0(_07645_),
    .A1(_07758_),
    .S(net9735),
    .X(_07759_));
 sg13g2_nor2_1 _30365_ (.A(net9726),
    .B(_07571_),
    .Y(_07760_));
 sg13g2_a21oi_2 _30366_ (.B1(_07760_),
    .Y(_07761_),
    .A2(_07759_),
    .A1(net9723));
 sg13g2_nand2_1 _30367_ (.Y(_07762_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[38] ),
    .B(_07761_));
 sg13g2_nor2_1 _30368_ (.A(_07753_),
    .B(_07762_),
    .Y(_07763_));
 sg13g2_a21oi_1 _30369_ (.A1(net9206),
    .A2(_07752_),
    .Y(_07764_),
    .B1(_07763_));
 sg13g2_xor2_1 _30370_ (.B(_07752_),
    .A(net9206),
    .X(_07765_));
 sg13g2_xor2_1 _30371_ (.B(_07761_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[38] ),
    .X(_07766_));
 sg13g2_nand2_1 _30372_ (.Y(_07767_),
    .A(_07765_),
    .B(_07766_));
 sg13g2_nand3_1 _30373_ (.B(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[6] ),
    .C(net8531),
    .A(net9760),
    .Y(_07768_));
 sg13g2_o21ai_1 _30374_ (.B1(_07768_),
    .Y(_07769_),
    .A1(net9761),
    .A2(_07754_));
 sg13g2_nor2_1 _30375_ (.A(net9066),
    .B(_07769_),
    .Y(_07770_));
 sg13g2_a21oi_1 _30376_ (.A1(net9066),
    .A2(_07746_),
    .Y(_07771_),
    .B1(_07770_));
 sg13g2_nand2_1 _30377_ (.Y(_07772_),
    .A(net9742),
    .B(_07771_));
 sg13g2_o21ai_1 _30378_ (.B1(_07772_),
    .Y(_07773_),
    .A1(net9742),
    .A2(_07717_));
 sg13g2_nand2b_1 _30379_ (.Y(_07774_),
    .B(net9072),
    .A_N(_07660_));
 sg13g2_o21ai_1 _30380_ (.B1(_07774_),
    .Y(_07775_),
    .A1(net9071),
    .A2(_07773_));
 sg13g2_nand2_1 _30381_ (.Y(_07776_),
    .A(net9723),
    .B(_07775_));
 sg13g2_nand2b_2 _30382_ (.Y(_07777_),
    .B(net9075),
    .A_N(_07584_));
 sg13g2_a21o_1 _30383_ (.A2(_07777_),
    .A1(_07776_),
    .B1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[37] ),
    .X(_07778_));
 sg13g2_nand2_1 _30384_ (.Y(_07779_),
    .A(net9074),
    .B(_07595_));
 sg13g2_nor3_1 _30385_ (.A(net9759),
    .B(_10624_),
    .C(net8581),
    .Y(_07780_));
 sg13g2_nor2b_1 _30386_ (.A(net8581),
    .B_N(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[5] ),
    .Y(_07781_));
 sg13g2_a21oi_1 _30387_ (.A1(net9759),
    .A2(_07781_),
    .Y(_07782_),
    .B1(_07780_));
 sg13g2_mux2_1 _30388_ (.A0(_07755_),
    .A1(_07782_),
    .S(net9750),
    .X(_07783_));
 sg13g2_nor2_1 _30389_ (.A(net9067),
    .B(_07783_),
    .Y(_07784_));
 sg13g2_a21oi_1 _30390_ (.A1(net9067),
    .A2(_07729_),
    .Y(_07785_),
    .B1(_07784_));
 sg13g2_nand2_1 _30391_ (.Y(_07786_),
    .A(net9735),
    .B(_07785_));
 sg13g2_o21ai_1 _30392_ (.B1(_07786_),
    .Y(_07787_),
    .A1(net9735),
    .A2(_07673_));
 sg13g2_o21ai_1 _30393_ (.B1(_07779_),
    .Y(_07788_),
    .A1(net9074),
    .A2(_07787_));
 sg13g2_nand2_1 _30394_ (.Y(_07789_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[36] ),
    .B(_07788_));
 sg13g2_nand3_1 _30395_ (.B(_07776_),
    .C(_07777_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[37] ),
    .Y(_07790_));
 sg13g2_nand2_1 _30396_ (.Y(_07791_),
    .A(_07789_),
    .B(_07790_));
 sg13g2_nand2_1 _30397_ (.Y(_07792_),
    .A(_07778_),
    .B(_07791_));
 sg13g2_and2_1 _30398_ (.A(_07778_),
    .B(_07790_),
    .X(_07793_));
 sg13g2_inv_1 _30399_ (.Y(_07794_),
    .A(_07793_));
 sg13g2_nor2_1 _30400_ (.A(_10623_),
    .B(net8580),
    .Y(_07795_));
 sg13g2_mux2_1 _30401_ (.A0(_07781_),
    .A1(_07795_),
    .S(net9761),
    .X(_07796_));
 sg13g2_mux2_1 _30402_ (.A0(_07769_),
    .A1(_07796_),
    .S(net9750),
    .X(_07797_));
 sg13g2_and2_1 _30403_ (.A(net9741),
    .B(_07797_),
    .X(_07798_));
 sg13g2_a21oi_1 _30404_ (.A1(net9069),
    .A2(_07748_),
    .Y(_07799_),
    .B1(_07798_));
 sg13g2_mux2_1 _30405_ (.A0(_07689_),
    .A1(_07799_),
    .S(net9733),
    .X(_07800_));
 sg13g2_nor2_1 _30406_ (.A(net9075),
    .B(_07800_),
    .Y(_07801_));
 sg13g2_a21oi_2 _30407_ (.B1(_07801_),
    .Y(_07802_),
    .A2(_07603_),
    .A1(net9075));
 sg13g2_and2_1 _30408_ (.A(_10637_),
    .B(_07802_),
    .X(_07803_));
 sg13g2_nand2b_1 _30409_ (.Y(_07804_),
    .B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[35] ),
    .A_N(_07802_));
 sg13g2_nor2_1 _30410_ (.A(net9741),
    .B(_07756_),
    .Y(_07805_));
 sg13g2_nor2b_1 _30411_ (.A(net8580),
    .B_N(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[3] ),
    .Y(_07806_));
 sg13g2_nand2b_1 _30412_ (.Y(_07807_),
    .B(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[3] ),
    .A_N(net8580));
 sg13g2_mux2_1 _30413_ (.A0(_07795_),
    .A1(_07806_),
    .S(net9762),
    .X(_07808_));
 sg13g2_nor2_1 _30414_ (.A(net9066),
    .B(_07808_),
    .Y(_07809_));
 sg13g2_a21oi_1 _30415_ (.A1(net9066),
    .A2(_07782_),
    .Y(_07810_),
    .B1(_07809_));
 sg13g2_a21oi_2 _30416_ (.B1(_07805_),
    .Y(_07811_),
    .A2(_07810_),
    .A1(net9741));
 sg13g2_mux2_1 _30417_ (.A0(_07701_),
    .A1(_07811_),
    .S(net9736),
    .X(_07812_));
 sg13g2_nor2_1 _30418_ (.A(net9075),
    .B(_07812_),
    .Y(_07813_));
 sg13g2_a21oi_2 _30419_ (.B1(_07813_),
    .Y(_07814_),
    .A2(_07614_),
    .A1(net9075));
 sg13g2_nand2b_1 _30420_ (.Y(_07815_),
    .B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[34] ),
    .A_N(_07814_));
 sg13g2_nor2_1 _30421_ (.A(net9728),
    .B(_07623_),
    .Y(_07816_));
 sg13g2_nand2b_1 _30422_ (.Y(_07817_),
    .B(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[2] ),
    .A_N(net8581));
 sg13g2_mux2_1 _30423_ (.A0(_07807_),
    .A1(_07817_),
    .S(net9760),
    .X(_07818_));
 sg13g2_nor2_1 _30424_ (.A(net9751),
    .B(_07796_),
    .Y(_07819_));
 sg13g2_a21oi_1 _30425_ (.A1(net9750),
    .A2(_07818_),
    .Y(_07820_),
    .B1(_07819_));
 sg13g2_mux2_1 _30426_ (.A0(_07771_),
    .A1(_07820_),
    .S(net9742),
    .X(_07821_));
 sg13g2_nor2_1 _30427_ (.A(net9073),
    .B(_07821_),
    .Y(_07822_));
 sg13g2_a21oi_2 _30428_ (.B1(_07822_),
    .Y(_07823_),
    .A2(_07719_),
    .A1(net9073));
 sg13g2_a21oi_2 _30429_ (.B1(_07816_),
    .Y(_07824_),
    .A2(_07823_),
    .A1(net9728));
 sg13g2_inv_1 _30430_ (.Y(_07825_),
    .A(_07824_));
 sg13g2_nor2_1 _30431_ (.A(net9072),
    .B(_07732_),
    .Y(_07826_));
 sg13g2_a21oi_2 _30432_ (.B1(_07826_),
    .Y(_07827_),
    .A2(_07548_),
    .A1(net9073));
 sg13g2_nor2_1 _30433_ (.A(net9741),
    .B(_07783_),
    .Y(_07828_));
 sg13g2_nor2b_1 _30434_ (.A(net8580),
    .B_N(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[1] ),
    .Y(_07829_));
 sg13g2_nand3b_1 _30435_ (.B(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[1] ),
    .C(net9760),
    .Y(_07830_),
    .A_N(net8580));
 sg13g2_o21ai_1 _30436_ (.B1(_07830_),
    .Y(_07831_),
    .A1(net9760),
    .A2(_07817_));
 sg13g2_mux2_1 _30437_ (.A0(_07808_),
    .A1(_07831_),
    .S(net9751),
    .X(_07832_));
 sg13g2_a21oi_2 _30438_ (.B1(_07828_),
    .Y(_07833_),
    .A2(_07832_),
    .A1(net9741));
 sg13g2_mux2_1 _30439_ (.A0(_07730_),
    .A1(_07833_),
    .S(net9735),
    .X(_07834_));
 sg13g2_nor2_1 _30440_ (.A(net9074),
    .B(_07834_),
    .Y(_07835_));
 sg13g2_a21oi_2 _30441_ (.B1(_07835_),
    .Y(_07836_),
    .A2(_07827_),
    .A1(net9074));
 sg13g2_nor2_1 _30442_ (.A(_10635_),
    .B(_07836_),
    .Y(_07837_));
 sg13g2_and2_1 _30443_ (.A(net9074),
    .B(_07634_),
    .X(_07838_));
 sg13g2_o21ai_1 _30444_ (.B1(net9759),
    .Y(_07839_),
    .A1(_10618_),
    .A2(net8580));
 sg13g2_o21ai_1 _30445_ (.B1(_07839_),
    .Y(_07840_),
    .A1(net9760),
    .A2(_07829_));
 sg13g2_mux2_1 _30446_ (.A0(_07818_),
    .A1(_07840_),
    .S(net9751),
    .X(_07841_));
 sg13g2_nor2_1 _30447_ (.A(net9069),
    .B(_07841_),
    .Y(_07842_));
 sg13g2_a21oi_1 _30448_ (.A1(net9069),
    .A2(_07797_),
    .Y(_07843_),
    .B1(_07842_));
 sg13g2_and2_1 _30449_ (.A(net9733),
    .B(_07843_),
    .X(_07844_));
 sg13g2_a21oi_2 _30450_ (.B1(_07844_),
    .Y(_07845_),
    .A2(_07749_),
    .A1(net9071));
 sg13g2_a21oi_2 _30451_ (.B1(_07838_),
    .Y(_07846_),
    .A2(_07845_),
    .A1(net9729));
 sg13g2_and2_1 _30452_ (.A(_10634_),
    .B(_07846_),
    .X(_07847_));
 sg13g2_nand2b_1 _30453_ (.Y(_07848_),
    .B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[31] ),
    .A_N(_07846_));
 sg13g2_nor2_1 _30454_ (.A(net9728),
    .B(_07647_),
    .Y(_07849_));
 sg13g2_nand2_1 _30455_ (.Y(_07850_),
    .A(net9068),
    .B(_07810_));
 sg13g2_nor4_1 _30456_ (.A(net9066),
    .B(net9761),
    .C(_10618_),
    .D(net8580),
    .Y(_07851_));
 sg13g2_a21oi_2 _30457_ (.B1(_07851_),
    .Y(_07852_),
    .A2(_07831_),
    .A1(net9066));
 sg13g2_o21ai_1 _30458_ (.B1(_07850_),
    .Y(_07853_),
    .A1(net9068),
    .A2(_07852_));
 sg13g2_nor2_1 _30459_ (.A(net9073),
    .B(_07853_),
    .Y(_07854_));
 sg13g2_a21oi_2 _30460_ (.B1(_07854_),
    .Y(_07855_),
    .A2(_07758_),
    .A1(net9072));
 sg13g2_a21oi_2 _30461_ (.B1(_07849_),
    .Y(_07856_),
    .A2(_07855_),
    .A1(net9727));
 sg13g2_nand2b_1 _30462_ (.Y(_07857_),
    .B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[30] ),
    .A_N(_07856_));
 sg13g2_o21ai_1 _30463_ (.B1(_07848_),
    .Y(_07858_),
    .A1(_07847_),
    .A2(_07857_));
 sg13g2_nor2b_1 _30464_ (.A(_07847_),
    .B_N(_07848_),
    .Y(_07859_));
 sg13g2_xnor2_1 _30465_ (.Y(_07860_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[30] ),
    .B(_07856_));
 sg13g2_and2_1 _30466_ (.A(_07859_),
    .B(_07860_),
    .X(_07861_));
 sg13g2_nor3_1 _30467_ (.A(net9069),
    .B(net9751),
    .C(_07840_),
    .Y(_07862_));
 sg13g2_a21oi_1 _30468_ (.A1(net9069),
    .A2(_07820_),
    .Y(_07863_),
    .B1(_07862_));
 sg13g2_nand2_1 _30469_ (.Y(_07864_),
    .A(net9733),
    .B(_07863_));
 sg13g2_o21ai_1 _30470_ (.B1(_07864_),
    .Y(_07865_),
    .A1(net9734),
    .A2(_07773_));
 sg13g2_nor2_1 _30471_ (.A(net9075),
    .B(_07865_),
    .Y(_07866_));
 sg13g2_a21oi_2 _30472_ (.B1(_07866_),
    .Y(_07867_),
    .A2(_07661_),
    .A1(net9074));
 sg13g2_and2_1 _30473_ (.A(_10632_),
    .B(_07867_),
    .X(_07868_));
 sg13g2_inv_1 _30474_ (.Y(_07869_),
    .A(_07868_));
 sg13g2_or4_2 _30475_ (.A(net9750),
    .B(net9761),
    .C(_10618_),
    .D(net8580),
    .X(_07870_));
 sg13g2_nor2_1 _30476_ (.A(net9069),
    .B(_07870_),
    .Y(_07871_));
 sg13g2_a21oi_2 _30477_ (.B1(_07871_),
    .Y(_07872_),
    .A2(_07832_),
    .A1(net9069));
 sg13g2_and2_1 _30478_ (.A(net9735),
    .B(_07872_),
    .X(_07873_));
 sg13g2_a21oi_1 _30479_ (.A1(net9073),
    .A2(_07785_),
    .Y(_07874_),
    .B1(_07873_));
 sg13g2_nand2_1 _30480_ (.Y(_07875_),
    .A(net9721),
    .B(_07874_));
 sg13g2_o21ai_1 _30481_ (.B1(_07875_),
    .Y(_07876_),
    .A1(net9721),
    .A2(_07675_));
 sg13g2_nand2_1 _30482_ (.Y(_07877_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[28] ),
    .B(_07876_));
 sg13g2_o21ai_1 _30483_ (.B1(_07877_),
    .Y(_07878_),
    .A1(_10632_),
    .A2(_07867_));
 sg13g2_nand2_1 _30484_ (.Y(_07879_),
    .A(_07869_),
    .B(_07878_));
 sg13g2_xnor2_1 _30485_ (.Y(_07880_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[29] ),
    .B(_07867_));
 sg13g2_xor2_1 _30486_ (.B(_07876_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[28] ),
    .X(_07881_));
 sg13g2_and2_1 _30487_ (.A(_07880_),
    .B(_07881_),
    .X(_07882_));
 sg13g2_inv_1 _30488_ (.Y(_07883_),
    .A(_07882_));
 sg13g2_or3_1 _30489_ (.A(net9071),
    .B(net9741),
    .C(_07841_),
    .X(_07884_));
 sg13g2_o21ai_1 _30490_ (.B1(_07884_),
    .Y(_07885_),
    .A1(net9733),
    .A2(_07799_));
 sg13g2_inv_2 _30491_ (.Y(_07886_),
    .A(_07885_));
 sg13g2_nand2_2 _30492_ (.Y(_07887_),
    .A(net9730),
    .B(_07886_));
 sg13g2_nand2_2 _30493_ (.Y(_07888_),
    .A(net9074),
    .B(_07691_));
 sg13g2_and3_1 _30494_ (.X(_07889_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[27] ),
    .B(_07887_),
    .C(_07888_));
 sg13g2_nand3_1 _30495_ (.B(_07887_),
    .C(_07888_),
    .A(net9205),
    .Y(_07890_));
 sg13g2_a21oi_1 _30496_ (.A1(_07887_),
    .A2(_07888_),
    .Y(_07891_),
    .B1(net9205));
 sg13g2_nor2_1 _30497_ (.A(net9720),
    .B(_07703_),
    .Y(_07892_));
 sg13g2_nor2_1 _30498_ (.A(net9748),
    .B(_07852_),
    .Y(_07893_));
 sg13g2_nand2_1 _30499_ (.Y(_07894_),
    .A(net9736),
    .B(_07893_));
 sg13g2_o21ai_1 _30500_ (.B1(_07894_),
    .Y(_07895_),
    .A1(net9736),
    .A2(_07811_));
 sg13g2_a21oi_2 _30501_ (.B1(_07892_),
    .Y(_07896_),
    .A2(_07895_),
    .A1(net9720));
 sg13g2_nand2b_1 _30502_ (.Y(_07897_),
    .B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[26] ),
    .A_N(_07896_));
 sg13g2_a21oi_1 _30503_ (.A1(_07890_),
    .A2(_07897_),
    .Y(_07898_),
    .B1(_07891_));
 sg13g2_xnor2_1 _30504_ (.Y(_07899_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[26] ),
    .B(_07896_));
 sg13g2_nor2_2 _30505_ (.A(_07889_),
    .B(_07891_),
    .Y(_07900_));
 sg13g2_or3_1 _30506_ (.A(net9071),
    .B(net9742),
    .C(_07870_),
    .X(_07901_));
 sg13g2_o21ai_1 _30507_ (.B1(_07901_),
    .Y(_07902_),
    .A1(net9733),
    .A2(_07833_));
 sg13g2_mux2_2 _30508_ (.A0(_07734_),
    .A1(_07902_),
    .S(net9720),
    .X(_07903_));
 sg13g2_nand2_1 _30509_ (.Y(_07904_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[24] ),
    .B(_07903_));
 sg13g2_nor4_1 _30510_ (.A(net9071),
    .B(net9741),
    .C(net9751),
    .D(_07840_),
    .Y(_07905_));
 sg13g2_a21oi_2 _30511_ (.B1(_07905_),
    .Y(_07906_),
    .A2(_07821_),
    .A1(net9071));
 sg13g2_nand2_2 _30512_ (.Y(_07907_),
    .A(net9722),
    .B(_07906_));
 sg13g2_or2_1 _30513_ (.X(_07908_),
    .B(_07721_),
    .A(net9730));
 sg13g2_nand3_1 _30514_ (.B(_07907_),
    .C(_07908_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[25] ),
    .Y(_07909_));
 sg13g2_nand2_1 _30515_ (.Y(_07910_),
    .A(_07904_),
    .B(_07909_));
 sg13g2_a21o_1 _30516_ (.A2(_07908_),
    .A1(_07907_),
    .B1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[25] ),
    .X(_07911_));
 sg13g2_nand2_1 _30517_ (.Y(_07912_),
    .A(_07910_),
    .B(_07911_));
 sg13g2_nand2_1 _30518_ (.Y(_07913_),
    .A(_07909_),
    .B(_07911_));
 sg13g2_nor2_1 _30519_ (.A(net9733),
    .B(_07843_),
    .Y(_07914_));
 sg13g2_mux2_2 _30520_ (.A0(_07751_),
    .A1(_07914_),
    .S(net9719),
    .X(_07915_));
 sg13g2_nand2_1 _30521_ (.Y(_07916_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[23] ),
    .B(_07915_));
 sg13g2_inv_1 _30522_ (.Y(_07917_),
    .A(_07916_));
 sg13g2_nor2_1 _30523_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[23] ),
    .B(_07915_),
    .Y(_07918_));
 sg13g2_and2_1 _30524_ (.A(net9071),
    .B(_07853_),
    .X(_07919_));
 sg13g2_nand2_1 _30525_ (.Y(_07920_),
    .A(net9720),
    .B(_07919_));
 sg13g2_o21ai_1 _30526_ (.B1(_07920_),
    .Y(_07921_),
    .A1(net9719),
    .A2(_07759_));
 sg13g2_nand2_1 _30527_ (.Y(_07922_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[22] ),
    .B(_07921_));
 sg13g2_xor2_1 _30528_ (.B(_07921_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[22] ),
    .X(_07923_));
 sg13g2_nor2_1 _30529_ (.A(net9733),
    .B(_07863_),
    .Y(_07924_));
 sg13g2_nand2_1 _30530_ (.Y(_07925_),
    .A(net9722),
    .B(_07924_));
 sg13g2_o21ai_1 _30531_ (.B1(_07925_),
    .Y(_07926_),
    .A1(net9722),
    .A2(_07775_));
 sg13g2_nor2_1 _30532_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[21] ),
    .B(_07926_),
    .Y(_07927_));
 sg13g2_nor3_1 _30533_ (.A(net9734),
    .B(net9743),
    .C(_07841_),
    .Y(_07928_));
 sg13g2_nand2_1 _30534_ (.Y(_07929_),
    .A(net9719),
    .B(_07928_));
 sg13g2_o21ai_1 _30535_ (.B1(_07929_),
    .Y(_07930_),
    .A1(net9719),
    .A2(_07800_));
 sg13g2_or2_1 _30536_ (.X(_07931_),
    .B(_07930_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[19] ));
 sg13g2_inv_1 _30537_ (.Y(_07932_),
    .A(_07931_));
 sg13g2_nand2_1 _30538_ (.Y(_07933_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[19] ),
    .B(_07930_));
 sg13g2_nand3_1 _30539_ (.B(net9071),
    .C(_07893_),
    .A(net9720),
    .Y(_07934_));
 sg13g2_o21ai_1 _30540_ (.B1(_07934_),
    .Y(_07935_),
    .A1(net9720),
    .A2(_07812_));
 sg13g2_and2_1 _30541_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[18] ),
    .B(_07935_),
    .X(_07936_));
 sg13g2_or4_2 _30542_ (.A(net9734),
    .B(net9743),
    .C(net9751),
    .D(_07840_),
    .X(_07937_));
 sg13g2_nor2_1 _30543_ (.A(net9727),
    .B(_07823_),
    .Y(_07938_));
 sg13g2_a21oi_1 _30544_ (.A1(net9721),
    .A2(_07937_),
    .Y(_07939_),
    .B1(_07938_));
 sg13g2_nor2_1 _30545_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[17] ),
    .B(_07939_),
    .Y(_07940_));
 sg13g2_nand2_1 _30546_ (.Y(_07941_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[17] ),
    .B(_07939_));
 sg13g2_nor3_2 _30547_ (.A(net9733),
    .B(net9742),
    .C(_07870_),
    .Y(_07942_));
 sg13g2_nand2_1 _30548_ (.Y(_07943_),
    .A(net9722),
    .B(_07942_));
 sg13g2_o21ai_1 _30549_ (.B1(_07943_),
    .Y(_07944_),
    .A1(net9721),
    .A2(_07834_));
 sg13g2_nand2_1 _30550_ (.Y(_07945_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[16] ),
    .B(_07944_));
 sg13g2_a21o_1 _30551_ (.A2(_07845_),
    .A1(net9717),
    .B1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[15] ),
    .X(_07946_));
 sg13g2_nand3_1 _30552_ (.B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[15] ),
    .C(_07845_),
    .A(net9717),
    .Y(_07947_));
 sg13g2_inv_1 _30553_ (.Y(_07948_),
    .A(_07947_));
 sg13g2_and2_1 _30554_ (.A(net9717),
    .B(_07855_),
    .X(_07949_));
 sg13g2_nor2_1 _30555_ (.A(_10607_),
    .B(_07865_),
    .Y(_07950_));
 sg13g2_nor3_1 _30556_ (.A(net8983),
    .B(_00268_),
    .C(_07865_),
    .Y(_07951_));
 sg13g2_nor2b_1 _30557_ (.A(_07950_),
    .B_N(_00268_),
    .Y(_07952_));
 sg13g2_nand2_1 _30558_ (.Y(_07953_),
    .A(net9717),
    .B(_07874_));
 sg13g2_inv_1 _30559_ (.Y(_07954_),
    .A(_07953_));
 sg13g2_a21oi_1 _30560_ (.A1(net9717),
    .A2(_07885_),
    .Y(_07955_),
    .B1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[11] ));
 sg13g2_nor3_2 _30561_ (.A(net8983),
    .B(_10626_),
    .C(_07886_),
    .Y(_07956_));
 sg13g2_or3_1 _30562_ (.A(net8983),
    .B(_00265_),
    .C(_07906_),
    .X(_07957_));
 sg13g2_o21ai_1 _30563_ (.B1(_00265_),
    .Y(_07958_),
    .A1(net8983),
    .A2(_07906_));
 sg13g2_nand2_2 _30564_ (.Y(_07959_),
    .A(net9716),
    .B(_07914_));
 sg13g2_or2_1 _30565_ (.X(_07960_),
    .B(_07959_),
    .A(_00263_));
 sg13g2_inv_1 _30566_ (.Y(_07961_),
    .A(_07960_));
 sg13g2_nand2_1 _30567_ (.Y(_07962_),
    .A(net9716),
    .B(_07924_));
 sg13g2_nor2_1 _30568_ (.A(_00261_),
    .B(_07962_),
    .Y(_07963_));
 sg13g2_and2_1 _30569_ (.A(net9716),
    .B(_07928_),
    .X(_07964_));
 sg13g2_nor2b_1 _30570_ (.A(_00259_),
    .B_N(_07964_),
    .Y(_07965_));
 sg13g2_nor3_1 _30571_ (.A(net8983),
    .B(_00257_),
    .C(_07937_),
    .Y(_07966_));
 sg13g2_nand2_1 _30572_ (.Y(_07967_),
    .A(net9716),
    .B(_07942_));
 sg13g2_nor2_1 _30573_ (.A(_00253_),
    .B(_07967_),
    .Y(_07968_));
 sg13g2_o21ai_1 _30574_ (.B1(_00257_),
    .Y(_07969_),
    .A1(net8983),
    .A2(_07937_));
 sg13g2_nor2b_1 _30575_ (.A(_07966_),
    .B_N(_07969_),
    .Y(_07970_));
 sg13g2_a21oi_1 _30576_ (.A1(_07968_),
    .A2(_07969_),
    .Y(_07971_),
    .B1(_07966_));
 sg13g2_nor4_2 _30577_ (.A(net9734),
    .B(net9743),
    .C(net8983),
    .Y(_07972_),
    .D(_07852_));
 sg13g2_xor2_1 _30578_ (.B(_07972_),
    .A(_00258_),
    .X(_07973_));
 sg13g2_or2_1 _30579_ (.X(_07974_),
    .B(_07973_),
    .A(_07971_));
 sg13g2_nand2_1 _30580_ (.Y(_07975_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[2] ),
    .B(_07972_));
 sg13g2_o21ai_1 _30581_ (.B1(_07975_),
    .Y(_07976_),
    .A1(_07971_),
    .A2(_07973_));
 sg13g2_nand2b_1 _30582_ (.Y(_07977_),
    .B(_00259_),
    .A_N(_07964_));
 sg13g2_nand2b_1 _30583_ (.Y(_07978_),
    .B(_07977_),
    .A_N(_07965_));
 sg13g2_a21oi_1 _30584_ (.A1(_07976_),
    .A2(_07977_),
    .Y(_07979_),
    .B1(_07965_));
 sg13g2_nor3_2 _30585_ (.A(net9734),
    .B(net8983),
    .C(_07872_),
    .Y(_07980_));
 sg13g2_xor2_1 _30586_ (.B(_07980_),
    .A(_00260_),
    .X(_07981_));
 sg13g2_nor2_1 _30587_ (.A(_07979_),
    .B(_07981_),
    .Y(_07982_));
 sg13g2_nand2_1 _30588_ (.Y(_07983_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[4] ),
    .B(_07980_));
 sg13g2_o21ai_1 _30589_ (.B1(_07983_),
    .Y(_07984_),
    .A1(_07979_),
    .A2(_07981_));
 sg13g2_nand2_1 _30590_ (.Y(_07985_),
    .A(_00261_),
    .B(_07962_));
 sg13g2_nor2b_1 _30591_ (.A(_07963_),
    .B_N(_07985_),
    .Y(_07986_));
 sg13g2_a21oi_1 _30592_ (.A1(_07984_),
    .A2(_07985_),
    .Y(_07987_),
    .B1(_07963_));
 sg13g2_and2_1 _30593_ (.A(net9716),
    .B(_07919_),
    .X(_07988_));
 sg13g2_xor2_1 _30594_ (.B(_07988_),
    .A(_00262_),
    .X(_07989_));
 sg13g2_nor2_1 _30595_ (.A(_07987_),
    .B(_07989_),
    .Y(_07990_));
 sg13g2_nand2_1 _30596_ (.Y(_07991_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[6] ),
    .B(_07988_));
 sg13g2_o21ai_1 _30597_ (.B1(_07991_),
    .Y(_07992_),
    .A1(_07987_),
    .A2(_07989_));
 sg13g2_nand2_1 _30598_ (.Y(_07993_),
    .A(_00263_),
    .B(_07959_));
 sg13g2_and2_1 _30599_ (.A(_07960_),
    .B(_07993_),
    .X(_07994_));
 sg13g2_a21oi_2 _30600_ (.B1(_07961_),
    .Y(_07995_),
    .A2(_07993_),
    .A1(_07992_));
 sg13g2_and2_1 _30601_ (.A(net9716),
    .B(_07902_),
    .X(_07996_));
 sg13g2_xor2_1 _30602_ (.B(_07996_),
    .A(_00264_),
    .X(_07997_));
 sg13g2_nor2_1 _30603_ (.A(_07995_),
    .B(_07997_),
    .Y(_07998_));
 sg13g2_nand2_1 _30604_ (.Y(_07999_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[8] ),
    .B(_07996_));
 sg13g2_nor2b_1 _30605_ (.A(_07998_),
    .B_N(_07999_),
    .Y(_08000_));
 sg13g2_and2_1 _30606_ (.A(_07957_),
    .B(_07999_),
    .X(_08001_));
 sg13g2_o21ai_1 _30607_ (.B1(_08001_),
    .Y(_08002_),
    .A1(_07995_),
    .A2(_07997_));
 sg13g2_nand2_1 _30608_ (.Y(_08003_),
    .A(_07958_),
    .B(_08002_));
 sg13g2_nand2_1 _30609_ (.Y(_08004_),
    .A(net9716),
    .B(_07895_));
 sg13g2_xnor2_1 _30610_ (.Y(_08005_),
    .A(_00266_),
    .B(_08004_));
 sg13g2_nand3b_1 _30611_ (.B(_08002_),
    .C(_07958_),
    .Y(_08006_),
    .A_N(_08005_));
 sg13g2_nand3_1 _30612_ (.B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[10] ),
    .C(_07895_),
    .A(net9717),
    .Y(_08007_));
 sg13g2_nand2_1 _30613_ (.Y(_08008_),
    .A(_08006_),
    .B(_08007_));
 sg13g2_a21oi_2 _30614_ (.B1(_07955_),
    .Y(_08009_),
    .A2(_08007_),
    .A1(_08006_));
 sg13g2_xor2_1 _30615_ (.B(_07953_),
    .A(_00267_),
    .X(_08010_));
 sg13g2_o21ai_1 _30616_ (.B1(_08010_),
    .Y(_08011_),
    .A1(_07956_),
    .A2(_08009_));
 sg13g2_o21ai_1 _30617_ (.B1(_08011_),
    .Y(_08012_),
    .A1(_10627_),
    .A2(_07953_));
 sg13g2_nor2_1 _30618_ (.A(_07951_),
    .B(_07952_),
    .Y(_08013_));
 sg13g2_and2_1 _30619_ (.A(_08010_),
    .B(_08013_),
    .X(_08014_));
 sg13g2_o21ai_1 _30620_ (.B1(_08014_),
    .Y(_08015_),
    .A1(_07956_),
    .A2(_08009_));
 sg13g2_a21oi_1 _30621_ (.A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[12] ),
    .A2(_07954_),
    .Y(_08016_),
    .B1(_07951_));
 sg13g2_or2_1 _30622_ (.X(_08017_),
    .B(_08016_),
    .A(_07952_));
 sg13g2_and2_1 _30623_ (.A(_08015_),
    .B(_08017_),
    .X(_08018_));
 sg13g2_xnor2_1 _30624_ (.Y(_08019_),
    .A(_00269_),
    .B(_07949_));
 sg13g2_nor2b_1 _30625_ (.A(_08018_),
    .B_N(_08019_),
    .Y(_08020_));
 sg13g2_a21o_1 _30626_ (.A2(_07949_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[14] ),
    .B1(_08020_),
    .X(_08021_));
 sg13g2_and3_1 _30627_ (.X(_08022_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[14] ),
    .B(_07946_),
    .C(_07949_));
 sg13g2_and2_1 _30628_ (.A(_07946_),
    .B(_07947_),
    .X(_08023_));
 sg13g2_nand2_1 _30629_ (.Y(_08024_),
    .A(_08019_),
    .B(_08023_));
 sg13g2_a21oi_1 _30630_ (.A1(_08015_),
    .A2(_08017_),
    .Y(_08025_),
    .B1(_08024_));
 sg13g2_nor3_2 _30631_ (.A(_07948_),
    .B(_08022_),
    .C(_08025_),
    .Y(_08026_));
 sg13g2_nor2_1 _30632_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[16] ),
    .B(_07944_),
    .Y(_08027_));
 sg13g2_xor2_1 _30633_ (.B(_07944_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[16] ),
    .X(_08028_));
 sg13g2_o21ai_1 _30634_ (.B1(_07945_),
    .Y(_08029_),
    .A1(_08026_),
    .A2(_08027_));
 sg13g2_o21ai_1 _30635_ (.B1(_07941_),
    .Y(_08030_),
    .A1(_07940_),
    .A2(_07945_));
 sg13g2_inv_1 _30636_ (.Y(_08031_),
    .A(_08030_));
 sg13g2_nor2b_1 _30637_ (.A(_07940_),
    .B_N(_07941_),
    .Y(_08032_));
 sg13g2_nand2_1 _30638_ (.Y(_08033_),
    .A(_08028_),
    .B(_08032_));
 sg13g2_o21ai_1 _30639_ (.B1(_08031_),
    .Y(_08034_),
    .A1(_08026_),
    .A2(_08033_));
 sg13g2_xor2_1 _30640_ (.B(_07935_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[18] ),
    .X(_08035_));
 sg13g2_a21oi_2 _30641_ (.B1(_07936_),
    .Y(_08036_),
    .A2(_08035_),
    .A1(_08034_));
 sg13g2_and2_1 _30642_ (.A(_07931_),
    .B(_07933_),
    .X(_08037_));
 sg13g2_inv_1 _30643_ (.Y(_08038_),
    .A(_08037_));
 sg13g2_a21oi_2 _30644_ (.B1(_07932_),
    .Y(_08039_),
    .A2(_08036_),
    .A1(_07933_));
 sg13g2_nand3b_1 _30645_ (.B(net9719),
    .C(net9072),
    .Y(_08040_),
    .A_N(_07872_));
 sg13g2_o21ai_1 _30646_ (.B1(_08040_),
    .Y(_08041_),
    .A1(net9719),
    .A2(_07787_));
 sg13g2_nand2_1 _30647_ (.Y(_08042_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[20] ),
    .B(_08041_));
 sg13g2_xor2_1 _30648_ (.B(_08041_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[20] ),
    .X(_08043_));
 sg13g2_nand2_1 _30649_ (.Y(_08044_),
    .A(_08039_),
    .B(_08043_));
 sg13g2_nand2_1 _30650_ (.Y(_08045_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[21] ),
    .B(_07926_));
 sg13g2_and2_1 _30651_ (.A(_08042_),
    .B(_08045_),
    .X(_08046_));
 sg13g2_a21oi_1 _30652_ (.A1(_08044_),
    .A2(_08046_),
    .Y(_08047_),
    .B1(_07927_));
 sg13g2_nand2_1 _30653_ (.Y(_08048_),
    .A(_07923_),
    .B(_08047_));
 sg13g2_nand2_1 _30654_ (.Y(_08049_),
    .A(_07922_),
    .B(_08048_));
 sg13g2_nor2_2 _30655_ (.A(_07917_),
    .B(_07918_),
    .Y(_08050_));
 sg13g2_nand2_1 _30656_ (.Y(_08051_),
    .A(_07923_),
    .B(_08050_));
 sg13g2_nor3_1 _30657_ (.A(_07927_),
    .B(_08046_),
    .C(_08051_),
    .Y(_08052_));
 sg13g2_nor2b_1 _30658_ (.A(_07927_),
    .B_N(_08045_),
    .Y(_08053_));
 sg13g2_and4_1 _30659_ (.A(_07923_),
    .B(_08043_),
    .C(_08050_),
    .D(_08053_),
    .X(_08054_));
 sg13g2_o21ai_1 _30660_ (.B1(_07916_),
    .Y(_08055_),
    .A1(_07918_),
    .A2(_07922_));
 sg13g2_or2_1 _30661_ (.X(_08056_),
    .B(_08055_),
    .A(_08052_));
 sg13g2_a21oi_2 _30662_ (.B1(_08056_),
    .Y(_08057_),
    .A2(_08054_),
    .A1(_08039_));
 sg13g2_xor2_1 _30663_ (.B(_07903_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[24] ),
    .X(_08058_));
 sg13g2_nand2b_2 _30664_ (.Y(_08059_),
    .B(_08058_),
    .A_N(_08057_));
 sg13g2_o21ai_1 _30665_ (.B1(_07912_),
    .Y(_08060_),
    .A1(_07913_),
    .A2(_08059_));
 sg13g2_nand4_1 _30666_ (.B(_07900_),
    .C(_07910_),
    .A(_07899_),
    .Y(_08061_),
    .D(_07911_));
 sg13g2_nor2b_1 _30667_ (.A(_07898_),
    .B_N(_08061_),
    .Y(_08062_));
 sg13g2_nand4_1 _30668_ (.B(_07900_),
    .C(_07909_),
    .A(_07899_),
    .Y(_08063_),
    .D(_07911_));
 sg13g2_o21ai_1 _30669_ (.B1(_08062_),
    .Y(_08064_),
    .A1(_08059_),
    .A2(_08063_));
 sg13g2_and2_1 _30670_ (.A(_07881_),
    .B(_08064_),
    .X(_08065_));
 sg13g2_o21ai_1 _30671_ (.B1(_07869_),
    .Y(_08066_),
    .A1(_07878_),
    .A2(_08065_));
 sg13g2_o21ai_1 _30672_ (.B1(_07879_),
    .Y(_08067_),
    .A1(_07883_),
    .A2(_08062_));
 sg13g2_a21oi_1 _30673_ (.A1(_07861_),
    .A2(_08067_),
    .Y(_08068_),
    .B1(_07858_));
 sg13g2_nand3_1 _30674_ (.B(_07882_),
    .C(_08058_),
    .A(_07861_),
    .Y(_08069_));
 sg13g2_or2_1 _30675_ (.X(_08070_),
    .B(_08069_),
    .A(_08063_));
 sg13g2_o21ai_1 _30676_ (.B1(_08068_),
    .Y(_08071_),
    .A1(_08057_),
    .A2(_08070_));
 sg13g2_xnor2_1 _30677_ (.Y(_08072_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[32] ),
    .B(_07836_));
 sg13g2_a21o_1 _30678_ (.A2(_08072_),
    .A1(_08071_),
    .B1(_07837_),
    .X(_08073_));
 sg13g2_a221oi_1 _30679_ (.B2(_08072_),
    .C1(_07837_),
    .B1(_08071_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[33] ),
    .Y(_08074_),
    .A2(_07825_));
 sg13g2_a21oi_2 _30680_ (.B1(_08074_),
    .Y(_08075_),
    .A2(_07824_),
    .A1(_10636_));
 sg13g2_xnor2_1 _30681_ (.Y(_08076_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[34] ),
    .B(_07814_));
 sg13g2_nand2_1 _30682_ (.Y(_08077_),
    .A(_08075_),
    .B(_08076_));
 sg13g2_nand2_1 _30683_ (.Y(_08078_),
    .A(_07815_),
    .B(_08077_));
 sg13g2_o21ai_1 _30684_ (.B1(_07804_),
    .Y(_08079_),
    .A1(_07803_),
    .A2(_07815_));
 sg13g2_nor2b_1 _30685_ (.A(_07803_),
    .B_N(_07804_),
    .Y(_08080_));
 sg13g2_and2_1 _30686_ (.A(_08076_),
    .B(_08080_),
    .X(_08081_));
 sg13g2_a21o_1 _30687_ (.A2(_08081_),
    .A1(_08075_),
    .B1(_08079_),
    .X(_08082_));
 sg13g2_a21oi_1 _30688_ (.A1(_08075_),
    .A2(_08081_),
    .Y(_08083_),
    .B1(_08079_));
 sg13g2_xnor2_1 _30689_ (.Y(_08084_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[36] ),
    .B(_07788_));
 sg13g2_nor2_1 _30690_ (.A(_08083_),
    .B(_08084_),
    .Y(_08085_));
 sg13g2_or2_1 _30691_ (.X(_08086_),
    .B(_08084_),
    .A(_08083_));
 sg13g2_o21ai_1 _30692_ (.B1(_07778_),
    .Y(_08087_),
    .A1(_07791_),
    .A2(_08085_));
 sg13g2_nor3_1 _30693_ (.A(_07767_),
    .B(_07794_),
    .C(_08084_),
    .Y(_08088_));
 sg13g2_o21ai_1 _30694_ (.B1(_07764_),
    .Y(_08089_),
    .A1(_07767_),
    .A2(_07792_));
 sg13g2_a21o_1 _30695_ (.A2(_08088_),
    .A1(_08082_),
    .B1(_08089_),
    .X(_08090_));
 sg13g2_xor2_1 _30696_ (.B(_07735_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[40] ),
    .X(_08091_));
 sg13g2_and2_1 _30697_ (.A(_08090_),
    .B(_08091_),
    .X(_08092_));
 sg13g2_and2_1 _30698_ (.A(_07743_),
    .B(_08092_),
    .X(_08093_));
 sg13g2_and4_1 _30699_ (.A(_07712_),
    .B(_07742_),
    .C(_07743_),
    .D(_08091_),
    .X(_08094_));
 sg13g2_a221oi_1 _30700_ (.B2(_08094_),
    .C1(_07741_),
    .B1(_08090_),
    .A1(_07653_),
    .Y(_08095_),
    .A2(_07740_));
 sg13g2_nand2_1 _30701_ (.Y(_08096_),
    .A(net9729),
    .B(_07827_));
 sg13g2_xor2_1 _30702_ (.B(_08096_),
    .A(_00270_),
    .X(_08097_));
 sg13g2_inv_1 _30703_ (.Y(_08098_),
    .A(_08097_));
 sg13g2_nand3_1 _30704_ (.B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[48] ),
    .C(_07827_),
    .A(net9729),
    .Y(_08099_));
 sg13g2_o21ai_1 _30705_ (.B1(_08099_),
    .Y(_08100_),
    .A1(_08095_),
    .A2(_08098_));
 sg13g2_a21oi_1 _30706_ (.A1(_07625_),
    .A2(_08100_),
    .Y(_08101_),
    .B1(_07624_));
 sg13g2_xnor2_1 _30707_ (.Y(_08102_),
    .A(_00272_),
    .B(_07615_));
 sg13g2_or2_1 _30708_ (.X(_08103_),
    .B(_08102_),
    .A(_08101_));
 sg13g2_and2_1 _30709_ (.A(_07616_),
    .B(_08103_),
    .X(_08104_));
 sg13g2_nand2b_1 _30710_ (.Y(_08105_),
    .B(_07605_),
    .A_N(_07604_));
 sg13g2_a21oi_1 _30711_ (.A1(_07605_),
    .A2(_08104_),
    .Y(_08106_),
    .B1(_07604_));
 sg13g2_xnor2_1 _30712_ (.Y(_08107_),
    .A(_00273_),
    .B(_07596_));
 sg13g2_nand2_1 _30713_ (.Y(_08108_),
    .A(_08106_),
    .B(_08107_));
 sg13g2_nand2_1 _30714_ (.Y(_08109_),
    .A(_07597_),
    .B(_08108_));
 sg13g2_nand2b_1 _30715_ (.Y(_08110_),
    .B(_07587_),
    .A_N(_07586_));
 sg13g2_a21oi_1 _30716_ (.A1(_07587_),
    .A2(_08109_),
    .Y(_08111_),
    .B1(_07586_));
 sg13g2_o21ai_1 _30717_ (.B1(_07573_),
    .Y(_08112_),
    .A1(_07575_),
    .A2(_08111_));
 sg13g2_nand2_1 _30718_ (.Y(_08113_),
    .A(_07561_),
    .B(_08112_));
 sg13g2_a21oi_1 _30719_ (.A1(_07560_),
    .A2(_08113_),
    .Y(_08114_),
    .B1(_07551_));
 sg13g2_a21o_1 _30720_ (.A2(_07550_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[56] ),
    .B1(_08114_),
    .X(_08115_));
 sg13g2_a21oi_1 _30721_ (.A1(_07538_),
    .A2(_08115_),
    .Y(_08116_),
    .B1(_07539_));
 sg13g2_nand2_1 _30722_ (.Y(_08117_),
    .A(net9724),
    .B(_07695_));
 sg13g2_xnor2_1 _30723_ (.Y(_08118_),
    .A(_00279_),
    .B(_08117_));
 sg13g2_or2_1 _30724_ (.X(_08119_),
    .B(_08118_),
    .A(_08116_));
 sg13g2_nand3_1 _30725_ (.B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[58] ),
    .C(_07695_),
    .A(net9724),
    .Y(_08120_));
 sg13g2_and2_1 _30726_ (.A(_08119_),
    .B(_08120_),
    .X(_08121_));
 sg13g2_nor2_1 _30727_ (.A(_07528_),
    .B(_08121_),
    .Y(_08122_));
 sg13g2_nand2_1 _30728_ (.Y(_08123_),
    .A(net9725),
    .B(_07666_));
 sg13g2_xor2_1 _30729_ (.B(_08123_),
    .A(_00281_),
    .X(_08124_));
 sg13g2_o21ai_1 _30730_ (.B1(_08124_),
    .Y(_08125_),
    .A1(_07527_),
    .A2(_08122_));
 sg13g2_nand3_1 _30731_ (.B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[60] ),
    .C(_07666_),
    .A(net9725),
    .Y(_08126_));
 sg13g2_nor3_2 _30732_ (.A(net9074),
    .B(net9731),
    .C(_07576_),
    .Y(_08127_));
 sg13g2_xor2_1 _30733_ (.B(_08127_),
    .A(_00282_),
    .X(_08128_));
 sg13g2_a21oi_1 _30734_ (.A1(_08125_),
    .A2(_08126_),
    .Y(_08129_),
    .B1(_08128_));
 sg13g2_a21oi_1 _30735_ (.A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[61] ),
    .A2(_08127_),
    .Y(_08130_),
    .B1(_08129_));
 sg13g2_a21o_1 _30736_ (.A2(_07515_),
    .A1(net9724),
    .B1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[62] ),
    .X(_08131_));
 sg13g2_nand2_1 _30737_ (.Y(_08132_),
    .A(_07516_),
    .B(_08131_));
 sg13g2_o21ai_1 _30738_ (.B1(_07516_),
    .Y(_08133_),
    .A1(_08130_),
    .A2(_08132_));
 sg13g2_o21ai_1 _30739_ (.B1(net9210),
    .Y(_08134_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[63] ),
    .A2(_08133_));
 sg13g2_a21oi_1 _30740_ (.A1(net5132),
    .A2(_08133_),
    .Y(_08135_),
    .B1(_08134_));
 sg13g2_nor3_2 _30741_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[0] ),
    .B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[1] ),
    .C(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[2] ),
    .Y(_08136_));
 sg13g2_nand2_1 _30742_ (.Y(_08137_),
    .A(_10621_),
    .B(_08136_));
 sg13g2_nand3_1 _30743_ (.B(_10622_),
    .C(_08136_),
    .A(_10621_),
    .Y(_08138_));
 sg13g2_or2_1 _30744_ (.X(_08139_),
    .B(_08138_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[5] ));
 sg13g2_nor2_1 _30745_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[6] ),
    .B(_08139_),
    .Y(_08140_));
 sg13g2_nand2b_1 _30746_ (.Y(_08141_),
    .B(_08140_),
    .A_N(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[7] ));
 sg13g2_or2_2 _30747_ (.X(_08142_),
    .B(_08141_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[8] ));
 sg13g2_or3_2 _30748_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[9] ),
    .B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[10] ),
    .C(_08142_),
    .X(_08143_));
 sg13g2_nor3_1 _30749_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[11] ),
    .B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[12] ),
    .C(_08143_),
    .Y(_08144_));
 sg13g2_nand2b_1 _30750_ (.Y(_08145_),
    .B(_08144_),
    .A_N(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[13] ));
 sg13g2_or2_2 _30751_ (.X(_08146_),
    .B(_08145_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[14] ));
 sg13g2_or3_2 _30752_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[15] ),
    .B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[16] ),
    .C(_08146_),
    .X(_08147_));
 sg13g2_nor3_2 _30753_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[17] ),
    .B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[18] ),
    .C(_08147_),
    .Y(_08148_));
 sg13g2_nand2b_2 _30754_ (.Y(_08149_),
    .B(_08148_),
    .A_N(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[19] ));
 sg13g2_or2_1 _30755_ (.X(_08150_),
    .B(_08149_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[20] ));
 sg13g2_or3_2 _30756_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[21] ),
    .B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[22] ),
    .C(_08150_),
    .X(_08151_));
 sg13g2_nor3_1 _30757_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[23] ),
    .B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[24] ),
    .C(_08151_),
    .Y(_08152_));
 sg13g2_nor2b_2 _30758_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[25] ),
    .B_N(_08152_),
    .Y(_08153_));
 sg13g2_nand2b_1 _30759_ (.Y(_08154_),
    .B(_08153_),
    .A_N(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[26] ));
 sg13g2_or3_2 _30760_ (.A(net9205),
    .B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[28] ),
    .C(_08154_),
    .X(_08155_));
 sg13g2_or3_2 _30761_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[29] ),
    .B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[30] ),
    .C(_08155_),
    .X(_08156_));
 sg13g2_nand3b_1 _30762_ (.B(_10635_),
    .C(_10634_),
    .Y(_08157_),
    .A_N(_08156_));
 sg13g2_or3_2 _30763_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[33] ),
    .B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[34] ),
    .C(_08157_),
    .X(_08158_));
 sg13g2_or3_1 _30764_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[35] ),
    .B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[36] ),
    .C(_08158_),
    .X(_08159_));
 sg13g2_nor2_1 _30765_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[37] ),
    .B(_08159_),
    .Y(_08160_));
 sg13g2_nand2b_1 _30766_ (.Y(_08161_),
    .B(_08160_),
    .A_N(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[38] ));
 sg13g2_or3_2 _30767_ (.A(net9206),
    .B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[40] ),
    .C(_08161_),
    .X(_08162_));
 sg13g2_or3_2 _30768_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[41] ),
    .B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[42] ),
    .C(_08162_),
    .X(_08163_));
 sg13g2_or3_2 _30769_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[43] ),
    .B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[44] ),
    .C(_08163_),
    .X(_08164_));
 sg13g2_or3_2 _30770_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[45] ),
    .B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[46] ),
    .C(_08164_),
    .X(_08165_));
 sg13g2_nor3_2 _30771_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[47] ),
    .B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[48] ),
    .C(_08165_),
    .Y(_08166_));
 sg13g2_nand2b_2 _30772_ (.Y(_08167_),
    .B(_08166_),
    .A_N(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[49] ));
 sg13g2_or2_1 _30773_ (.X(_08168_),
    .B(_08167_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[50] ));
 sg13g2_or3_1 _30774_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[51] ),
    .B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[52] ),
    .C(_08168_),
    .X(_08169_));
 sg13g2_nor2_1 _30775_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[53] ),
    .B(_08169_),
    .Y(_08170_));
 sg13g2_nand2b_1 _30776_ (.Y(_08171_),
    .B(_08170_),
    .A_N(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[54] ));
 sg13g2_or2_1 _30777_ (.X(_08172_),
    .B(_08171_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[55] ));
 sg13g2_or2_2 _30778_ (.X(_08173_),
    .B(_08172_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[56] ));
 sg13g2_or3_2 _30779_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[57] ),
    .B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[58] ),
    .C(_08173_),
    .X(_08174_));
 sg13g2_nor3_2 _30780_ (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[59] ),
    .B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[60] ),
    .C(_08174_),
    .Y(_08175_));
 sg13g2_nand2b_1 _30781_ (.Y(_08176_),
    .B(_08175_),
    .A_N(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[61] ));
 sg13g2_or2_1 _30782_ (.X(_08177_),
    .B(_08176_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[62] ));
 sg13g2_o21ai_1 _30783_ (.B1(net9218),
    .Y(_08178_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[63] ),
    .A2(_08177_));
 sg13g2_a21oi_1 _30784_ (.A1(net5132),
    .A2(_08177_),
    .Y(_08179_),
    .B1(_08178_));
 sg13g2_nand2_1 _30785_ (.Y(_08180_),
    .A(net9209),
    .B(net7712));
 sg13g2_a21oi_2 _30786_ (.B1(net7755),
    .Y(_08181_),
    .A2(net8987),
    .A1(net9077));
 sg13g2_o21ai_1 _30787_ (.B1(net7710),
    .Y(_08182_),
    .A1(net9221),
    .A2(net9212));
 sg13g2_o21ai_1 _30788_ (.B1(net7708),
    .Y(_08183_),
    .A1(_08135_),
    .A2(_08179_));
 sg13g2_o21ai_1 _30789_ (.B1(_08183_),
    .Y(_02145_),
    .A1(_10643_),
    .A2(net7710));
 sg13g2_nand2_1 _30790_ (.Y(_08184_),
    .A(net4615),
    .B(net7753));
 sg13g2_xor2_1 _30791_ (.B(_08132_),
    .A(_08130_),
    .X(_08185_));
 sg13g2_a21oi_1 _30792_ (.A1(net4615),
    .A2(_08176_),
    .Y(_08186_),
    .B1(net9077));
 sg13g2_a22oi_1 _30793_ (.Y(_08187_),
    .B1(_08186_),
    .B2(_08177_),
    .A2(_08185_),
    .A1(net9211));
 sg13g2_o21ai_1 _30794_ (.B1(_08184_),
    .Y(_02146_),
    .A1(net7693),
    .A2(_08187_));
 sg13g2_nand2_1 _30795_ (.Y(_08188_),
    .A(net4807),
    .B(net7753));
 sg13g2_nand3_1 _30796_ (.B(_08126_),
    .C(_08128_),
    .A(_08125_),
    .Y(_08189_));
 sg13g2_nor2_1 _30797_ (.A(net8987),
    .B(_08129_),
    .Y(_08190_));
 sg13g2_xnor2_1 _30798_ (.Y(_08191_),
    .A(net4807),
    .B(_08175_));
 sg13g2_a22oi_1 _30799_ (.Y(_08192_),
    .B1(_08191_),
    .B2(net9219),
    .A2(_08190_),
    .A1(_08189_));
 sg13g2_o21ai_1 _30800_ (.B1(_08188_),
    .Y(_02147_),
    .A1(net7693),
    .A2(_08192_));
 sg13g2_nand2_1 _30801_ (.Y(_08193_),
    .A(net4949),
    .B(net7752));
 sg13g2_or3_1 _30802_ (.A(_07527_),
    .B(_08122_),
    .C(_08124_),
    .X(_08194_));
 sg13g2_and2_1 _30803_ (.A(net9210),
    .B(_08125_),
    .X(_08195_));
 sg13g2_o21ai_1 _30804_ (.B1(net4949),
    .Y(_08196_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[59] ),
    .A2(_08174_));
 sg13g2_nor2_1 _30805_ (.A(net9077),
    .B(_08175_),
    .Y(_08197_));
 sg13g2_a22oi_1 _30806_ (.Y(_08198_),
    .B1(_08196_),
    .B2(_08197_),
    .A2(_08195_),
    .A1(_08194_));
 sg13g2_o21ai_1 _30807_ (.B1(_08193_),
    .Y(_02148_),
    .A1(net7692),
    .A2(_08198_));
 sg13g2_nand2_1 _30808_ (.Y(_08199_),
    .A(net5102),
    .B(net7753));
 sg13g2_nand2_1 _30809_ (.Y(_08200_),
    .A(_07528_),
    .B(_08121_));
 sg13g2_nor2_1 _30810_ (.A(net8987),
    .B(_08122_),
    .Y(_08201_));
 sg13g2_xor2_1 _30811_ (.B(_08174_),
    .A(net5102),
    .X(_08202_));
 sg13g2_a22oi_1 _30812_ (.Y(_08203_),
    .B1(_08202_),
    .B2(net9218),
    .A2(_08201_),
    .A1(_08200_));
 sg13g2_o21ai_1 _30813_ (.B1(_08199_),
    .Y(_02149_),
    .A1(net7692),
    .A2(_08203_));
 sg13g2_nand2_1 _30814_ (.Y(_08204_),
    .A(_08116_),
    .B(_08118_));
 sg13g2_nand3_1 _30815_ (.B(_08119_),
    .C(_08204_),
    .A(net9210),
    .Y(_08205_));
 sg13g2_o21ai_1 _30816_ (.B1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[58] ),
    .Y(_08206_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[57] ),
    .A2(_08173_));
 sg13g2_nand3_1 _30817_ (.B(_08174_),
    .C(_08206_),
    .A(net9218),
    .Y(_08207_));
 sg13g2_a21oi_1 _30818_ (.A1(_08205_),
    .A2(_08207_),
    .Y(_08208_),
    .B1(net7692));
 sg13g2_a21o_1 _30819_ (.A2(net7752),
    .A1(net4887),
    .B1(_08208_),
    .X(_02150_));
 sg13g2_xor2_1 _30820_ (.B(_07537_),
    .A(_00278_),
    .X(_08209_));
 sg13g2_o21ai_1 _30821_ (.B1(net9210),
    .Y(_08210_),
    .A1(_08115_),
    .A2(_08209_));
 sg13g2_a21oi_1 _30822_ (.A1(_08115_),
    .A2(_08209_),
    .Y(_08211_),
    .B1(_08210_));
 sg13g2_o21ai_1 _30823_ (.B1(net9218),
    .Y(_08212_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[57] ),
    .A2(_08173_));
 sg13g2_a21oi_1 _30824_ (.A1(net5111),
    .A2(_08173_),
    .Y(_08213_),
    .B1(_08212_));
 sg13g2_o21ai_1 _30825_ (.B1(net7708),
    .Y(_08214_),
    .A1(_08211_),
    .A2(_08213_));
 sg13g2_o21ai_1 _30826_ (.B1(_08214_),
    .Y(_02151_),
    .A1(_10642_),
    .A2(net7710));
 sg13g2_nand2_1 _30827_ (.Y(_08215_),
    .A(net4531),
    .B(net7752));
 sg13g2_nand3_1 _30828_ (.B(_07560_),
    .C(_08113_),
    .A(_07551_),
    .Y(_08216_));
 sg13g2_nor2_1 _30829_ (.A(net8987),
    .B(_08114_),
    .Y(_08217_));
 sg13g2_a21oi_1 _30830_ (.A1(net4531),
    .A2(_08172_),
    .Y(_08218_),
    .B1(net9077));
 sg13g2_a22oi_1 _30831_ (.Y(_08219_),
    .B1(_08218_),
    .B2(_08173_),
    .A2(_08217_),
    .A1(_08216_));
 sg13g2_o21ai_1 _30832_ (.B1(_08215_),
    .Y(_02152_),
    .A1(net7692),
    .A2(_08219_));
 sg13g2_a21oi_1 _30833_ (.A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[55] ),
    .A2(_08171_),
    .Y(_08220_),
    .B1(net9077));
 sg13g2_nand2_1 _30834_ (.Y(_08221_),
    .A(_08172_),
    .B(_08220_));
 sg13g2_nand3_1 _30835_ (.B(_07561_),
    .C(_08112_),
    .A(_07560_),
    .Y(_08222_));
 sg13g2_a21oi_1 _30836_ (.A1(_07560_),
    .A2(_07561_),
    .Y(_08223_),
    .B1(_08112_));
 sg13g2_nand2_1 _30837_ (.Y(_08224_),
    .A(net9210),
    .B(_08222_));
 sg13g2_o21ai_1 _30838_ (.B1(_08221_),
    .Y(_08225_),
    .A1(_08223_),
    .A2(_08224_));
 sg13g2_a22oi_1 _30839_ (.Y(_08226_),
    .B1(net7708),
    .B2(_08225_),
    .A2(net7752),
    .A1(net4658));
 sg13g2_inv_1 _30840_ (.Y(_02153_),
    .A(net4659));
 sg13g2_nand2_1 _30841_ (.Y(_08227_),
    .A(net4772),
    .B(net7752));
 sg13g2_xnor2_1 _30842_ (.Y(_08228_),
    .A(net4772),
    .B(_08170_));
 sg13g2_xnor2_1 _30843_ (.Y(_08229_),
    .A(_07574_),
    .B(_08111_));
 sg13g2_a22oi_1 _30844_ (.Y(_08230_),
    .B1(_08229_),
    .B2(net9210),
    .A2(_08228_),
    .A1(net9218));
 sg13g2_o21ai_1 _30845_ (.B1(_08227_),
    .Y(_02154_),
    .A1(net7692),
    .A2(_08230_));
 sg13g2_nand2_1 _30846_ (.Y(_08231_),
    .A(net3860),
    .B(net7752));
 sg13g2_xnor2_1 _30847_ (.Y(_08232_),
    .A(_08109_),
    .B(_08110_));
 sg13g2_nand2_1 _30848_ (.Y(_08233_),
    .A(net3860),
    .B(_08169_));
 sg13g2_nor2_1 _30849_ (.A(net9077),
    .B(_08170_),
    .Y(_08234_));
 sg13g2_a22oi_1 _30850_ (.Y(_08235_),
    .B1(_08233_),
    .B2(_08234_),
    .A2(_08232_),
    .A1(net9210));
 sg13g2_o21ai_1 _30851_ (.B1(_08231_),
    .Y(_02155_),
    .A1(net7692),
    .A2(_08235_));
 sg13g2_o21ai_1 _30852_ (.B1(net9211),
    .Y(_08236_),
    .A1(_08106_),
    .A2(_08107_));
 sg13g2_nand2b_1 _30853_ (.Y(_08237_),
    .B(_08108_),
    .A_N(_08236_));
 sg13g2_o21ai_1 _30854_ (.B1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[52] ),
    .Y(_08238_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[51] ),
    .A2(_08168_));
 sg13g2_nand3_1 _30855_ (.B(_08169_),
    .C(_08238_),
    .A(net9218),
    .Y(_08239_));
 sg13g2_a21oi_1 _30856_ (.A1(_08237_),
    .A2(_08239_),
    .Y(_08240_),
    .B1(net7693));
 sg13g2_a21o_1 _30857_ (.A2(net7752),
    .A1(net4928),
    .B1(_08240_),
    .X(_02156_));
 sg13g2_o21ai_1 _30858_ (.B1(net9211),
    .Y(_08241_),
    .A1(_08104_),
    .A2(_08105_));
 sg13g2_a21oi_1 _30859_ (.A1(_08104_),
    .A2(_08105_),
    .Y(_08242_),
    .B1(_08241_));
 sg13g2_o21ai_1 _30860_ (.B1(net9219),
    .Y(_08243_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[51] ),
    .A2(_08168_));
 sg13g2_a21oi_1 _30861_ (.A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[51] ),
    .A2(_08168_),
    .Y(_08244_),
    .B1(_08243_));
 sg13g2_o21ai_1 _30862_ (.B1(net7708),
    .Y(_08245_),
    .A1(_08242_),
    .A2(_08244_));
 sg13g2_o21ai_1 _30863_ (.B1(_08245_),
    .Y(_02157_),
    .A1(_10641_),
    .A2(net7710));
 sg13g2_nand2_1 _30864_ (.Y(_08246_),
    .A(net4834),
    .B(net7754));
 sg13g2_xor2_1 _30865_ (.B(_08167_),
    .A(net4834),
    .X(_08247_));
 sg13g2_a21oi_1 _30866_ (.A1(_08101_),
    .A2(_08102_),
    .Y(_08248_),
    .B1(net8986));
 sg13g2_a22oi_1 _30867_ (.Y(_08249_),
    .B1(_08248_),
    .B2(_08103_),
    .A2(_08247_),
    .A1(net9220));
 sg13g2_o21ai_1 _30868_ (.B1(_08246_),
    .Y(_02158_),
    .A1(net7693),
    .A2(_08249_));
 sg13g2_nand2_1 _30869_ (.Y(_08250_),
    .A(net4367),
    .B(net7754));
 sg13g2_nor2b_1 _30870_ (.A(_07624_),
    .B_N(_07625_),
    .Y(_08251_));
 sg13g2_xor2_1 _30871_ (.B(_08251_),
    .A(_08100_),
    .X(_08252_));
 sg13g2_nor2b_1 _30872_ (.A(_08166_),
    .B_N(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[49] ),
    .Y(_08253_));
 sg13g2_nor2_1 _30873_ (.A(net9078),
    .B(_08253_),
    .Y(_08254_));
 sg13g2_a22oi_1 _30874_ (.Y(_08255_),
    .B1(_08254_),
    .B2(_08167_),
    .A2(_08252_),
    .A1(net9213));
 sg13g2_o21ai_1 _30875_ (.B1(_08250_),
    .Y(_02159_),
    .A1(net7694),
    .A2(_08255_));
 sg13g2_nand2_1 _30876_ (.Y(_08256_),
    .A(net4666),
    .B(net7754));
 sg13g2_o21ai_1 _30877_ (.B1(net4666),
    .Y(_08257_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[47] ),
    .A2(_08165_));
 sg13g2_nor2_1 _30878_ (.A(_10508_),
    .B(_08166_),
    .Y(_08258_));
 sg13g2_xnor2_1 _30879_ (.Y(_08259_),
    .A(_08095_),
    .B(_08097_));
 sg13g2_a22oi_1 _30880_ (.Y(_08260_),
    .B1(_08259_),
    .B2(net9213),
    .A2(_08258_),
    .A1(_08257_));
 sg13g2_o21ai_1 _30881_ (.B1(_08256_),
    .Y(_02160_),
    .A1(net7694),
    .A2(_08260_));
 sg13g2_o21ai_1 _30882_ (.B1(_07710_),
    .Y(_08261_),
    .A1(_07738_),
    .A2(_08093_));
 sg13g2_a21oi_1 _30883_ (.A1(_07708_),
    .A2(_08261_),
    .Y(_08262_),
    .B1(_07694_));
 sg13g2_and2_1 _30884_ (.A(_07682_),
    .B(_08262_),
    .X(_08263_));
 sg13g2_o21ai_1 _30885_ (.B1(_07664_),
    .Y(_08264_),
    .A1(_07679_),
    .A2(_08263_));
 sg13g2_or2_1 _30886_ (.X(_08265_),
    .B(_08264_),
    .A(_07652_));
 sg13g2_and2_1 _30887_ (.A(_07650_),
    .B(_08265_),
    .X(_08266_));
 sg13g2_o21ai_1 _30888_ (.B1(net9213),
    .Y(_08267_),
    .A1(_07637_),
    .A2(_08266_));
 sg13g2_a21oi_1 _30889_ (.A1(_07637_),
    .A2(_08266_),
    .Y(_08268_),
    .B1(_08267_));
 sg13g2_o21ai_1 _30890_ (.B1(net9222),
    .Y(_08269_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[47] ),
    .A2(_08165_));
 sg13g2_a21oi_1 _30891_ (.A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[47] ),
    .A2(_08165_),
    .Y(_08270_),
    .B1(_08269_));
 sg13g2_o21ai_1 _30892_ (.B1(net7707),
    .Y(_08271_),
    .A1(_08268_),
    .A2(_08270_));
 sg13g2_o21ai_1 _30893_ (.B1(_08271_),
    .Y(_02161_),
    .A1(_10640_),
    .A2(net7711));
 sg13g2_a21oi_1 _30894_ (.A1(_07652_),
    .A2(_08264_),
    .Y(_08272_),
    .B1(net8986));
 sg13g2_nand2_1 _30895_ (.Y(_08273_),
    .A(_08265_),
    .B(_08272_));
 sg13g2_o21ai_1 _30896_ (.B1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[46] ),
    .Y(_08274_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[45] ),
    .A2(_08164_));
 sg13g2_nand3_1 _30897_ (.B(_08165_),
    .C(_08274_),
    .A(net9220),
    .Y(_08275_));
 sg13g2_a21oi_1 _30898_ (.A1(_08273_),
    .A2(_08275_),
    .Y(_08276_),
    .B1(net7694));
 sg13g2_a21o_1 _30899_ (.A2(net7754),
    .A1(net5288),
    .B1(_08276_),
    .X(_02162_));
 sg13g2_a21o_1 _30900_ (.A2(_07677_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[44] ),
    .B1(_08263_),
    .X(_08277_));
 sg13g2_o21ai_1 _30901_ (.B1(net9213),
    .Y(_08278_),
    .A1(_07681_),
    .A2(_08277_));
 sg13g2_a21oi_1 _30902_ (.A1(_07681_),
    .A2(_08277_),
    .Y(_08279_),
    .B1(_08278_));
 sg13g2_o21ai_1 _30903_ (.B1(net9220),
    .Y(_08280_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[45] ),
    .A2(_08164_));
 sg13g2_a21oi_1 _30904_ (.A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[45] ),
    .A2(_08164_),
    .Y(_08281_),
    .B1(_08280_));
 sg13g2_o21ai_1 _30905_ (.B1(net7707),
    .Y(_08282_),
    .A1(_08279_),
    .A2(_08281_));
 sg13g2_o21ai_1 _30906_ (.B1(_08282_),
    .Y(_02163_),
    .A1(_10639_),
    .A2(net7712));
 sg13g2_nor2_1 _30907_ (.A(net8986),
    .B(_08263_),
    .Y(_08283_));
 sg13g2_o21ai_1 _30908_ (.B1(_08283_),
    .Y(_08284_),
    .A1(_07682_),
    .A2(_08262_));
 sg13g2_o21ai_1 _30909_ (.B1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[44] ),
    .Y(_08285_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[43] ),
    .A2(_08163_));
 sg13g2_nand3_1 _30910_ (.B(_08164_),
    .C(_08285_),
    .A(net9214),
    .Y(_08286_));
 sg13g2_a21oi_1 _30911_ (.A1(_08284_),
    .A2(_08286_),
    .Y(_08287_),
    .B1(net7691));
 sg13g2_a21o_1 _30912_ (.A2(net7750),
    .A1(net5461),
    .B1(_08287_),
    .X(_02164_));
 sg13g2_and2_1 _30913_ (.A(_07706_),
    .B(_08261_),
    .X(_08288_));
 sg13g2_nand2b_1 _30914_ (.Y(_08289_),
    .B(_08288_),
    .A_N(_07711_));
 sg13g2_nand2b_1 _30915_ (.Y(_08290_),
    .B(_07711_),
    .A_N(_08288_));
 sg13g2_nand3_1 _30916_ (.B(_08289_),
    .C(_08290_),
    .A(net9208),
    .Y(_08291_));
 sg13g2_o21ai_1 _30917_ (.B1(net9216),
    .Y(_08292_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[43] ),
    .A2(_08163_));
 sg13g2_a21o_1 _30918_ (.A2(_08163_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[43] ),
    .B1(_08292_),
    .X(_08293_));
 sg13g2_a21oi_1 _30919_ (.A1(_08291_),
    .A2(_08293_),
    .Y(_08294_),
    .B1(net7691));
 sg13g2_a21o_1 _30920_ (.A2(net7750),
    .A1(net5484),
    .B1(_08294_),
    .X(_02165_));
 sg13g2_o21ai_1 _30921_ (.B1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[42] ),
    .Y(_08295_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[41] ),
    .A2(_08162_));
 sg13g2_nand3_1 _30922_ (.B(_08163_),
    .C(_08295_),
    .A(net9214),
    .Y(_08296_));
 sg13g2_or3_1 _30923_ (.A(_07710_),
    .B(_07738_),
    .C(_08093_),
    .X(_08297_));
 sg13g2_nand3_1 _30924_ (.B(_08261_),
    .C(_08297_),
    .A(net9208),
    .Y(_08298_));
 sg13g2_a21oi_1 _30925_ (.A1(_08296_),
    .A2(_08298_),
    .Y(_08299_),
    .B1(net7691));
 sg13g2_a21o_1 _30926_ (.A2(net7750),
    .A1(net5379),
    .B1(_08299_),
    .X(_02166_));
 sg13g2_nand2_1 _30927_ (.Y(_08300_),
    .A(net5353),
    .B(net7750));
 sg13g2_nor3_1 _30928_ (.A(_07736_),
    .B(_07743_),
    .C(_08092_),
    .Y(_08301_));
 sg13g2_o21ai_1 _30929_ (.B1(_07743_),
    .Y(_08302_),
    .A1(_07736_),
    .A2(_08092_));
 sg13g2_nor2_1 _30930_ (.A(net8985),
    .B(_08301_),
    .Y(_08303_));
 sg13g2_o21ai_1 _30931_ (.B1(net9216),
    .Y(_08304_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[41] ),
    .A2(_08162_));
 sg13g2_a21oi_1 _30932_ (.A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[41] ),
    .A2(_08162_),
    .Y(_08305_),
    .B1(_08304_));
 sg13g2_a21oi_1 _30933_ (.A1(_08302_),
    .A2(_08303_),
    .Y(_08306_),
    .B1(_08305_));
 sg13g2_o21ai_1 _30934_ (.B1(_08300_),
    .Y(_02167_),
    .A1(net7691),
    .A2(_08306_));
 sg13g2_o21ai_1 _30935_ (.B1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[40] ),
    .Y(_08307_),
    .A1(net9206),
    .A2(_08161_));
 sg13g2_nand3_1 _30936_ (.B(_08162_),
    .C(_08307_),
    .A(net9216),
    .Y(_08308_));
 sg13g2_nor2_1 _30937_ (.A(net8985),
    .B(_08092_),
    .Y(_08309_));
 sg13g2_o21ai_1 _30938_ (.B1(_08309_),
    .Y(_08310_),
    .A1(_08090_),
    .A2(_08091_));
 sg13g2_a21oi_1 _30939_ (.A1(_08308_),
    .A2(_08310_),
    .Y(_08311_),
    .B1(net7690));
 sg13g2_a21o_1 _30940_ (.A2(net7750),
    .A1(net5372),
    .B1(_08311_),
    .X(_02168_));
 sg13g2_nand2b_1 _30941_ (.Y(_08312_),
    .B(_07766_),
    .A_N(_08087_));
 sg13g2_and2_1 _30942_ (.A(_07762_),
    .B(_08312_),
    .X(_08313_));
 sg13g2_nand2b_1 _30943_ (.Y(_08314_),
    .B(_08313_),
    .A_N(_07765_));
 sg13g2_nand2b_1 _30944_ (.Y(_08315_),
    .B(_07765_),
    .A_N(_08313_));
 sg13g2_nand3_1 _30945_ (.B(_08314_),
    .C(_08315_),
    .A(net9207),
    .Y(_08316_));
 sg13g2_o21ai_1 _30946_ (.B1(net9215),
    .Y(_08317_),
    .A1(net9206),
    .A2(_08161_));
 sg13g2_a21o_1 _30947_ (.A2(_08161_),
    .A1(net9206),
    .B1(_08317_),
    .X(_08318_));
 sg13g2_a21oi_1 _30948_ (.A1(_08316_),
    .A2(_08318_),
    .Y(_08319_),
    .B1(net7690));
 sg13g2_a21o_1 _30949_ (.A2(net7749),
    .A1(net9206),
    .B1(_08319_),
    .X(_02169_));
 sg13g2_nand2_1 _30950_ (.Y(_08320_),
    .A(net5114),
    .B(net7749));
 sg13g2_xnor2_1 _30951_ (.Y(_08321_),
    .A(_07766_),
    .B(_08087_));
 sg13g2_xnor2_1 _30952_ (.Y(_08322_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[38] ),
    .B(_08160_));
 sg13g2_a22oi_1 _30953_ (.Y(_08323_),
    .B1(_08322_),
    .B2(net9215),
    .A2(_08321_),
    .A1(net9207));
 sg13g2_o21ai_1 _30954_ (.B1(_08320_),
    .Y(_02170_),
    .A1(net7690),
    .A2(_08323_));
 sg13g2_nand2_1 _30955_ (.Y(_08324_),
    .A(_07789_),
    .B(_08086_));
 sg13g2_o21ai_1 _30956_ (.B1(net9207),
    .Y(_08325_),
    .A1(_07793_),
    .A2(_08324_));
 sg13g2_a21oi_1 _30957_ (.A1(_07793_),
    .A2(_08324_),
    .Y(_08326_),
    .B1(_08325_));
 sg13g2_o21ai_1 _30958_ (.B1(net9215),
    .Y(_08327_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[37] ),
    .A2(_08159_));
 sg13g2_a21oi_1 _30959_ (.A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[37] ),
    .A2(_08159_),
    .Y(_08328_),
    .B1(_08327_));
 sg13g2_o21ai_1 _30960_ (.B1(net7709),
    .Y(_08329_),
    .A1(_08326_),
    .A2(_08328_));
 sg13g2_o21ai_1 _30961_ (.B1(_08329_),
    .Y(_02171_),
    .A1(_10638_),
    .A2(net7712));
 sg13g2_o21ai_1 _30962_ (.B1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[36] ),
    .Y(_08330_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[35] ),
    .A2(_08158_));
 sg13g2_nand3_1 _30963_ (.B(_08159_),
    .C(_08330_),
    .A(net9215),
    .Y(_08331_));
 sg13g2_nand2_1 _30964_ (.Y(_08332_),
    .A(_08083_),
    .B(_08084_));
 sg13g2_nand3_1 _30965_ (.B(_08086_),
    .C(_08332_),
    .A(net9207),
    .Y(_08333_));
 sg13g2_a21oi_1 _30966_ (.A1(_08331_),
    .A2(_08333_),
    .Y(_08334_),
    .B1(net7690));
 sg13g2_a21o_1 _30967_ (.A2(net7749),
    .A1(net5472),
    .B1(_08334_),
    .X(_02172_));
 sg13g2_o21ai_1 _30968_ (.B1(net9208),
    .Y(_08335_),
    .A1(_08078_),
    .A2(_08080_));
 sg13g2_a21oi_1 _30969_ (.A1(_08078_),
    .A2(_08080_),
    .Y(_08336_),
    .B1(_08335_));
 sg13g2_o21ai_1 _30970_ (.B1(net9214),
    .Y(_08337_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[35] ),
    .A2(_08158_));
 sg13g2_a21oi_1 _30971_ (.A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[35] ),
    .A2(_08158_),
    .Y(_08338_),
    .B1(_08337_));
 sg13g2_o21ai_1 _30972_ (.B1(net7709),
    .Y(_08339_),
    .A1(_08336_),
    .A2(_08338_));
 sg13g2_o21ai_1 _30973_ (.B1(_08339_),
    .Y(_02173_),
    .A1(_10637_),
    .A2(net7712));
 sg13g2_xnor2_1 _30974_ (.Y(_08340_),
    .A(_08075_),
    .B(_08076_));
 sg13g2_o21ai_1 _30975_ (.B1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[34] ),
    .Y(_08341_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[33] ),
    .A2(_08157_));
 sg13g2_nand3_1 _30976_ (.B(_08158_),
    .C(_08341_),
    .A(net9214),
    .Y(_08342_));
 sg13g2_o21ai_1 _30977_ (.B1(_08342_),
    .Y(_08343_),
    .A1(net8984),
    .A2(_08340_));
 sg13g2_a22oi_1 _30978_ (.Y(_08344_),
    .B1(net7709),
    .B2(_08343_),
    .A2(net7750),
    .A1(net5405));
 sg13g2_inv_1 _30979_ (.Y(_02174_),
    .A(_08344_));
 sg13g2_xnor2_1 _30980_ (.Y(_08345_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[33] ),
    .B(_07824_));
 sg13g2_o21ai_1 _30981_ (.B1(net9213),
    .Y(_08346_),
    .A1(_08073_),
    .A2(_08345_));
 sg13g2_a21oi_1 _30982_ (.A1(_08073_),
    .A2(_08345_),
    .Y(_08347_),
    .B1(_08346_));
 sg13g2_o21ai_1 _30983_ (.B1(net9220),
    .Y(_08348_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[33] ),
    .A2(_08157_));
 sg13g2_a21oi_1 _30984_ (.A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[33] ),
    .A2(_08157_),
    .Y(_08349_),
    .B1(_08348_));
 sg13g2_o21ai_1 _30985_ (.B1(net7707),
    .Y(_08350_),
    .A1(_08347_),
    .A2(_08349_));
 sg13g2_o21ai_1 _30986_ (.B1(_08350_),
    .Y(_02175_),
    .A1(_10636_),
    .A2(net7710));
 sg13g2_xnor2_1 _30987_ (.Y(_08351_),
    .A(_08071_),
    .B(_08072_));
 sg13g2_o21ai_1 _30988_ (.B1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[32] ),
    .Y(_08352_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[31] ),
    .A2(_08156_));
 sg13g2_nand3_1 _30989_ (.B(_08157_),
    .C(_08352_),
    .A(net9220),
    .Y(_08353_));
 sg13g2_o21ai_1 _30990_ (.B1(_08353_),
    .Y(_08354_),
    .A1(net8986),
    .A2(_08351_));
 sg13g2_nand2_1 _30991_ (.Y(_08355_),
    .A(net7707),
    .B(_08354_));
 sg13g2_o21ai_1 _30992_ (.B1(_08355_),
    .Y(_02176_),
    .A1(_10635_),
    .A2(net7711));
 sg13g2_nand2b_1 _30993_ (.Y(_08356_),
    .B(_07860_),
    .A_N(_08066_));
 sg13g2_nand2_1 _30994_ (.Y(_08357_),
    .A(_07857_),
    .B(_08356_));
 sg13g2_o21ai_1 _30995_ (.B1(net9212),
    .Y(_08358_),
    .A1(_07859_),
    .A2(_08357_));
 sg13g2_a21oi_1 _30996_ (.A1(_07859_),
    .A2(_08357_),
    .Y(_08359_),
    .B1(_08358_));
 sg13g2_o21ai_1 _30997_ (.B1(net9221),
    .Y(_08360_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[31] ),
    .A2(_08156_));
 sg13g2_a21oi_1 _30998_ (.A1(net5335),
    .A2(_08156_),
    .Y(_08361_),
    .B1(_08360_));
 sg13g2_o21ai_1 _30999_ (.B1(net7707),
    .Y(_08362_),
    .A1(_08359_),
    .A2(_08361_));
 sg13g2_o21ai_1 _31000_ (.B1(_08362_),
    .Y(_02177_),
    .A1(_10634_),
    .A2(net7711));
 sg13g2_nand2_1 _31001_ (.Y(_08363_),
    .A(net5122),
    .B(net7755));
 sg13g2_xnor2_1 _31002_ (.Y(_08364_),
    .A(_07860_),
    .B(_08066_));
 sg13g2_o21ai_1 _31003_ (.B1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[30] ),
    .Y(_08365_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[29] ),
    .A2(_08155_));
 sg13g2_and2_1 _31004_ (.A(net9221),
    .B(_08365_),
    .X(_08366_));
 sg13g2_a22oi_1 _31005_ (.Y(_08367_),
    .B1(_08366_),
    .B2(_08156_),
    .A2(_08364_),
    .A1(net9213));
 sg13g2_o21ai_1 _31006_ (.B1(_08363_),
    .Y(_02178_),
    .A1(net7694),
    .A2(_08367_));
 sg13g2_a21o_1 _31007_ (.A2(_07876_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[28] ),
    .B1(_08065_),
    .X(_08368_));
 sg13g2_o21ai_1 _31008_ (.B1(net9212),
    .Y(_08369_),
    .A1(_07880_),
    .A2(_08368_));
 sg13g2_a21oi_1 _31009_ (.A1(_07880_),
    .A2(_08368_),
    .Y(_08370_),
    .B1(_08369_));
 sg13g2_o21ai_1 _31010_ (.B1(net9221),
    .Y(_08371_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[29] ),
    .A2(_08155_));
 sg13g2_a21oi_1 _31011_ (.A1(net5427),
    .A2(_08155_),
    .Y(_08372_),
    .B1(_08371_));
 sg13g2_o21ai_1 _31012_ (.B1(_08181_),
    .Y(_08373_),
    .A1(_08370_),
    .A2(_08372_));
 sg13g2_o21ai_1 _31013_ (.B1(_08373_),
    .Y(_02179_),
    .A1(_10632_),
    .A2(net7711));
 sg13g2_o21ai_1 _31014_ (.B1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[28] ),
    .Y(_08374_),
    .A1(net9205),
    .A2(_08154_));
 sg13g2_nand3_1 _31015_ (.B(_08155_),
    .C(_08374_),
    .A(net9221),
    .Y(_08375_));
 sg13g2_o21ai_1 _31016_ (.B1(net9212),
    .Y(_08376_),
    .A1(_07881_),
    .A2(_08064_));
 sg13g2_o21ai_1 _31017_ (.B1(_08375_),
    .Y(_08377_),
    .A1(_08065_),
    .A2(_08376_));
 sg13g2_a22oi_1 _31018_ (.Y(_08378_),
    .B1(_08181_),
    .B2(_08377_),
    .A2(net7755),
    .A1(net5334));
 sg13g2_inv_1 _31019_ (.Y(_02180_),
    .A(_08378_));
 sg13g2_nand2_1 _31020_ (.Y(_08379_),
    .A(_07899_),
    .B(_08060_));
 sg13g2_nand2_1 _31021_ (.Y(_08380_),
    .A(_07897_),
    .B(_08379_));
 sg13g2_o21ai_1 _31022_ (.B1(net9212),
    .Y(_08381_),
    .A1(_07900_),
    .A2(_08380_));
 sg13g2_a21o_1 _31023_ (.A2(_08380_),
    .A1(_07900_),
    .B1(_08381_),
    .X(_08382_));
 sg13g2_o21ai_1 _31024_ (.B1(net9221),
    .Y(_08383_),
    .A1(net9205),
    .A2(_08154_));
 sg13g2_a21o_1 _31025_ (.A2(_08154_),
    .A1(net9205),
    .B1(_08383_),
    .X(_08384_));
 sg13g2_a21oi_1 _31026_ (.A1(_08382_),
    .A2(_08384_),
    .Y(_08385_),
    .B1(net7694));
 sg13g2_a21o_1 _31027_ (.A2(net7755),
    .A1(net9205),
    .B1(_08385_),
    .X(_02181_));
 sg13g2_nand2_1 _31028_ (.Y(_08386_),
    .A(net5254),
    .B(net7755));
 sg13g2_xor2_1 _31029_ (.B(_08060_),
    .A(_07899_),
    .X(_08387_));
 sg13g2_xnor2_1 _31030_ (.Y(_08388_),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[26] ),
    .B(_08153_));
 sg13g2_a22oi_1 _31031_ (.Y(_08389_),
    .B1(_08388_),
    .B2(net9221),
    .A2(_08387_),
    .A1(net9212));
 sg13g2_o21ai_1 _31032_ (.B1(_08386_),
    .Y(_02182_),
    .A1(net7694),
    .A2(_08389_));
 sg13g2_nand2_1 _31033_ (.Y(_08390_),
    .A(net5192),
    .B(net7755));
 sg13g2_nand3_1 _31034_ (.B(_07913_),
    .C(_08059_),
    .A(_07904_),
    .Y(_08391_));
 sg13g2_a21oi_1 _31035_ (.A1(_07904_),
    .A2(_08059_),
    .Y(_08392_),
    .B1(_07913_));
 sg13g2_nor2_1 _31036_ (.A(net8986),
    .B(_08392_),
    .Y(_08393_));
 sg13g2_nand2b_1 _31037_ (.Y(_08394_),
    .B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[25] ),
    .A_N(_08152_));
 sg13g2_nor2_1 _31038_ (.A(net9077),
    .B(_08153_),
    .Y(_08395_));
 sg13g2_a22oi_1 _31039_ (.Y(_08396_),
    .B1(_08394_),
    .B2(_08395_),
    .A2(_08393_),
    .A1(_08391_));
 sg13g2_o21ai_1 _31040_ (.B1(_08390_),
    .Y(_02183_),
    .A1(net7694),
    .A2(_08396_));
 sg13g2_o21ai_1 _31041_ (.B1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[24] ),
    .Y(_08397_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[23] ),
    .A2(_08151_));
 sg13g2_nand2_1 _31042_ (.Y(_08398_),
    .A(net9219),
    .B(_08397_));
 sg13g2_nand2b_1 _31043_ (.Y(_08399_),
    .B(_08057_),
    .A_N(_08058_));
 sg13g2_nand3_1 _31044_ (.B(_08059_),
    .C(_08399_),
    .A(net9212),
    .Y(_08400_));
 sg13g2_o21ai_1 _31045_ (.B1(_08400_),
    .Y(_08401_),
    .A1(_08152_),
    .A2(_08398_));
 sg13g2_a22oi_1 _31046_ (.Y(_08402_),
    .B1(net7708),
    .B2(_08401_),
    .A2(net7754),
    .A1(net5356));
 sg13g2_inv_1 _31047_ (.Y(_02184_),
    .A(_08402_));
 sg13g2_o21ai_1 _31048_ (.B1(net9211),
    .Y(_08403_),
    .A1(_08049_),
    .A2(_08050_));
 sg13g2_a21oi_1 _31049_ (.A1(_08049_),
    .A2(_08050_),
    .Y(_08404_),
    .B1(_08403_));
 sg13g2_o21ai_1 _31050_ (.B1(net9218),
    .Y(_08405_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[23] ),
    .A2(_08151_));
 sg13g2_a21oi_1 _31051_ (.A1(net5378),
    .A2(_08151_),
    .Y(_08406_),
    .B1(_08405_));
 sg13g2_o21ai_1 _31052_ (.B1(net7708),
    .Y(_08407_),
    .A1(_08404_),
    .A2(_08406_));
 sg13g2_o21ai_1 _31053_ (.B1(_08407_),
    .Y(_02185_),
    .A1(_10631_),
    .A2(net7710));
 sg13g2_nand2_1 _31054_ (.Y(_08408_),
    .A(net4969),
    .B(net7752));
 sg13g2_xor2_1 _31055_ (.B(_08047_),
    .A(_07923_),
    .X(_08409_));
 sg13g2_o21ai_1 _31056_ (.B1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[22] ),
    .Y(_08410_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[21] ),
    .A2(_08150_));
 sg13g2_and2_1 _31057_ (.A(_08151_),
    .B(_08410_),
    .X(_08411_));
 sg13g2_a22oi_1 _31058_ (.Y(_08412_),
    .B1(_08411_),
    .B2(net9219),
    .A2(_08409_),
    .A1(net9211));
 sg13g2_o21ai_1 _31059_ (.B1(_08408_),
    .Y(_02186_),
    .A1(net7692),
    .A2(_08412_));
 sg13g2_o21ai_1 _31060_ (.B1(net9218),
    .Y(_08413_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[21] ),
    .A2(_08150_));
 sg13g2_a21oi_1 _31061_ (.A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[21] ),
    .A2(_08150_),
    .Y(_08414_),
    .B1(_08413_));
 sg13g2_nand2_1 _31062_ (.Y(_08415_),
    .A(_08042_),
    .B(_08044_));
 sg13g2_o21ai_1 _31063_ (.B1(net9210),
    .Y(_08416_),
    .A1(_08053_),
    .A2(_08415_));
 sg13g2_a21oi_1 _31064_ (.A1(_08053_),
    .A2(_08415_),
    .Y(_08417_),
    .B1(_08416_));
 sg13g2_o21ai_1 _31065_ (.B1(net7708),
    .Y(_08418_),
    .A1(_08414_),
    .A2(_08417_));
 sg13g2_o21ai_1 _31066_ (.B1(_08418_),
    .Y(_02187_),
    .A1(_10630_),
    .A2(net7710));
 sg13g2_a21oi_1 _31067_ (.A1(_08039_),
    .A2(_08043_),
    .Y(_08419_),
    .B1(net8987));
 sg13g2_o21ai_1 _31068_ (.B1(_08419_),
    .Y(_08420_),
    .A1(_08039_),
    .A2(_08043_));
 sg13g2_a21oi_1 _31069_ (.A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[20] ),
    .A2(_08149_),
    .Y(_08421_),
    .B1(net9077));
 sg13g2_nand2_1 _31070_ (.Y(_08422_),
    .A(_08150_),
    .B(_08421_));
 sg13g2_a21oi_1 _31071_ (.A1(_08420_),
    .A2(_08422_),
    .Y(_08423_),
    .B1(net7692));
 sg13g2_a21o_1 _31072_ (.A2(net7753),
    .A1(net5161),
    .B1(_08423_),
    .X(_02188_));
 sg13g2_a21oi_1 _31073_ (.A1(_08036_),
    .A2(_08038_),
    .Y(_08424_),
    .B1(net8986));
 sg13g2_o21ai_1 _31074_ (.B1(_08424_),
    .Y(_08425_),
    .A1(_08036_),
    .A2(_08038_));
 sg13g2_nand2b_1 _31075_ (.Y(_08426_),
    .B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[19] ),
    .A_N(_08148_));
 sg13g2_nand3_1 _31076_ (.B(_08149_),
    .C(_08426_),
    .A(net9221),
    .Y(_08427_));
 sg13g2_a21oi_1 _31077_ (.A1(_08425_),
    .A2(_08427_),
    .Y(_08428_),
    .B1(net7695));
 sg13g2_a21o_1 _31078_ (.A2(net7754),
    .A1(net5092),
    .B1(_08428_),
    .X(_02189_));
 sg13g2_xnor2_1 _31079_ (.Y(_08429_),
    .A(_08034_),
    .B(_08035_));
 sg13g2_o21ai_1 _31080_ (.B1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[18] ),
    .Y(_08430_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[17] ),
    .A2(_08147_));
 sg13g2_nand3b_1 _31081_ (.B(_08430_),
    .C(net9220),
    .Y(_08431_),
    .A_N(_08148_));
 sg13g2_o21ai_1 _31082_ (.B1(_08431_),
    .Y(_08432_),
    .A1(net8986),
    .A2(_08429_));
 sg13g2_a22oi_1 _31083_ (.Y(_08433_),
    .B1(net7707),
    .B2(_08432_),
    .A2(net7754),
    .A1(net5121));
 sg13g2_inv_1 _31084_ (.Y(_02190_),
    .A(_08433_));
 sg13g2_o21ai_1 _31085_ (.B1(net9213),
    .Y(_08434_),
    .A1(_08029_),
    .A2(_08032_));
 sg13g2_a21oi_1 _31086_ (.A1(_08029_),
    .A2(_08032_),
    .Y(_08435_),
    .B1(_08434_));
 sg13g2_o21ai_1 _31087_ (.B1(net9220),
    .Y(_08436_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[17] ),
    .A2(_08147_));
 sg13g2_a21oi_1 _31088_ (.A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[17] ),
    .A2(_08147_),
    .Y(_08437_),
    .B1(_08436_));
 sg13g2_o21ai_1 _31089_ (.B1(net7707),
    .Y(_08438_),
    .A1(_08435_),
    .A2(_08437_));
 sg13g2_o21ai_1 _31090_ (.B1(_08438_),
    .Y(_02191_),
    .A1(_10629_),
    .A2(net7710));
 sg13g2_xor2_1 _31091_ (.B(_08028_),
    .A(_08026_),
    .X(_08439_));
 sg13g2_o21ai_1 _31092_ (.B1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[16] ),
    .Y(_08440_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[15] ),
    .A2(_08146_));
 sg13g2_nand3_1 _31093_ (.B(_08147_),
    .C(_08440_),
    .A(net9220),
    .Y(_08441_));
 sg13g2_o21ai_1 _31094_ (.B1(_08441_),
    .Y(_08442_),
    .A1(net8986),
    .A2(_08439_));
 sg13g2_a22oi_1 _31095_ (.Y(_08443_),
    .B1(net7707),
    .B2(_08442_),
    .A2(net7754),
    .A1(net5112));
 sg13g2_inv_1 _31096_ (.Y(_02192_),
    .A(_08443_));
 sg13g2_o21ai_1 _31097_ (.B1(net9208),
    .Y(_08444_),
    .A1(_08021_),
    .A2(_08023_));
 sg13g2_a21oi_1 _31098_ (.A1(_08021_),
    .A2(_08023_),
    .Y(_08445_),
    .B1(_08444_));
 sg13g2_o21ai_1 _31099_ (.B1(net9214),
    .Y(_08446_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[15] ),
    .A2(_08146_));
 sg13g2_a21oi_1 _31100_ (.A1(net5264),
    .A2(_08146_),
    .Y(_08447_),
    .B1(_08446_));
 sg13g2_o21ai_1 _31101_ (.B1(net7709),
    .Y(_08448_),
    .A1(_08445_),
    .A2(_08447_));
 sg13g2_o21ai_1 _31102_ (.B1(_08448_),
    .Y(_02193_),
    .A1(_10628_),
    .A2(net7712));
 sg13g2_nand2_1 _31103_ (.Y(_08449_),
    .A(net4729),
    .B(net7750));
 sg13g2_xnor2_1 _31104_ (.Y(_08450_),
    .A(_08018_),
    .B(_08019_));
 sg13g2_a21oi_1 _31105_ (.A1(net4729),
    .A2(_08145_),
    .Y(_08451_),
    .B1(net9078));
 sg13g2_a22oi_1 _31106_ (.Y(_08452_),
    .B1(_08451_),
    .B2(_08146_),
    .A2(_08450_),
    .A1(net9208));
 sg13g2_o21ai_1 _31107_ (.B1(_08449_),
    .Y(_02194_),
    .A1(net7691),
    .A2(_08452_));
 sg13g2_a21oi_1 _31108_ (.A1(_08012_),
    .A2(_08013_),
    .Y(_08453_),
    .B1(net8985));
 sg13g2_o21ai_1 _31109_ (.B1(_08453_),
    .Y(_08454_),
    .A1(_08012_),
    .A2(_08013_));
 sg13g2_nand2b_1 _31110_ (.Y(_08455_),
    .B(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[13] ),
    .A_N(_08144_));
 sg13g2_nand3_1 _31111_ (.B(_08145_),
    .C(_08455_),
    .A(net9214),
    .Y(_08456_));
 sg13g2_a21oi_1 _31112_ (.A1(_08454_),
    .A2(_08456_),
    .Y(_08457_),
    .B1(net7691));
 sg13g2_a21o_1 _31113_ (.A2(net7750),
    .A1(net4297),
    .B1(_08457_),
    .X(_02195_));
 sg13g2_or3_1 _31114_ (.A(_07956_),
    .B(_08009_),
    .C(_08010_),
    .X(_08458_));
 sg13g2_nand3_1 _31115_ (.B(_08011_),
    .C(_08458_),
    .A(net9208),
    .Y(_08459_));
 sg13g2_o21ai_1 _31116_ (.B1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[12] ),
    .Y(_08460_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[11] ),
    .A2(_08143_));
 sg13g2_nand3b_1 _31117_ (.B(_08460_),
    .C(net9214),
    .Y(_08461_),
    .A_N(_08144_));
 sg13g2_a21o_1 _31118_ (.A2(_08461_),
    .A1(_08459_),
    .B1(net7691),
    .X(_08462_));
 sg13g2_o21ai_1 _31119_ (.B1(_08462_),
    .Y(_02196_),
    .A1(_10627_),
    .A2(net7712));
 sg13g2_nor2_1 _31120_ (.A(_07955_),
    .B(_07956_),
    .Y(_08463_));
 sg13g2_o21ai_1 _31121_ (.B1(net9207),
    .Y(_08464_),
    .A1(_08008_),
    .A2(_08463_));
 sg13g2_a21oi_1 _31122_ (.A1(_08008_),
    .A2(_08463_),
    .Y(_08465_),
    .B1(_08464_));
 sg13g2_o21ai_1 _31123_ (.B1(net9214),
    .Y(_08466_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[11] ),
    .A2(_08143_));
 sg13g2_a21oi_1 _31124_ (.A1(net5425),
    .A2(_08143_),
    .Y(_08467_),
    .B1(_08466_));
 sg13g2_o21ai_1 _31125_ (.B1(net7709),
    .Y(_08468_),
    .A1(_08465_),
    .A2(_08467_));
 sg13g2_o21ai_1 _31126_ (.B1(_08468_),
    .Y(_02197_),
    .A1(_10626_),
    .A2(net7712));
 sg13g2_nand2_1 _31127_ (.Y(_08469_),
    .A(net4160),
    .B(net7749));
 sg13g2_xor2_1 _31128_ (.B(_08005_),
    .A(_08003_),
    .X(_08470_));
 sg13g2_o21ai_1 _31129_ (.B1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[10] ),
    .Y(_08471_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[9] ),
    .A2(_08142_));
 sg13g2_and2_1 _31130_ (.A(_08143_),
    .B(_08471_),
    .X(_08472_));
 sg13g2_a22oi_1 _31131_ (.Y(_08473_),
    .B1(_08472_),
    .B2(net9215),
    .A2(_08470_),
    .A1(net9207));
 sg13g2_o21ai_1 _31132_ (.B1(_08469_),
    .Y(_02198_),
    .A1(net7690),
    .A2(_08473_));
 sg13g2_nand2_1 _31133_ (.Y(_08474_),
    .A(_07957_),
    .B(_07958_));
 sg13g2_o21ai_1 _31134_ (.B1(net9207),
    .Y(_08475_),
    .A1(_08000_),
    .A2(_08474_));
 sg13g2_a21oi_1 _31135_ (.A1(_08000_),
    .A2(_08474_),
    .Y(_08476_),
    .B1(_08475_));
 sg13g2_o21ai_1 _31136_ (.B1(net9215),
    .Y(_08477_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[9] ),
    .A2(_08142_));
 sg13g2_a21oi_1 _31137_ (.A1(net5083),
    .A2(_08142_),
    .Y(_08478_),
    .B1(_08477_));
 sg13g2_o21ai_1 _31138_ (.B1(net7709),
    .Y(_08479_),
    .A1(_08476_),
    .A2(_08478_));
 sg13g2_o21ai_1 _31139_ (.B1(_08479_),
    .Y(_02199_),
    .A1(_10625_),
    .A2(net7712));
 sg13g2_nand2_1 _31140_ (.Y(_08480_),
    .A(_07995_),
    .B(_07997_));
 sg13g2_nand3b_1 _31141_ (.B(_08480_),
    .C(net9207),
    .Y(_08481_),
    .A_N(_07998_));
 sg13g2_a21oi_1 _31142_ (.A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[8] ),
    .A2(_08141_),
    .Y(_08482_),
    .B1(net9078));
 sg13g2_nand2_1 _31143_ (.Y(_08483_),
    .A(_08142_),
    .B(_08482_));
 sg13g2_nand2_1 _31144_ (.Y(_08484_),
    .A(_08481_),
    .B(_08483_));
 sg13g2_a22oi_1 _31145_ (.Y(_08485_),
    .B1(net7709),
    .B2(_08484_),
    .A2(net7749),
    .A1(net4324));
 sg13g2_inv_1 _31146_ (.Y(_02200_),
    .A(net4325));
 sg13g2_nand2_1 _31147_ (.Y(_08486_),
    .A(net3971),
    .B(net7749));
 sg13g2_nor2_1 _31148_ (.A(_07992_),
    .B(_07994_),
    .Y(_08487_));
 sg13g2_a21o_1 _31149_ (.A2(_07994_),
    .A1(_07992_),
    .B1(net8984),
    .X(_08488_));
 sg13g2_nor2_1 _31150_ (.A(_08487_),
    .B(_08488_),
    .Y(_08489_));
 sg13g2_xnor2_1 _31151_ (.Y(_08490_),
    .A(net3971),
    .B(_08140_));
 sg13g2_a21oi_1 _31152_ (.A1(net9215),
    .A2(_08490_),
    .Y(_08491_),
    .B1(_08489_));
 sg13g2_o21ai_1 _31153_ (.B1(_08486_),
    .Y(_02201_),
    .A1(net7690),
    .A2(_08491_));
 sg13g2_nand2_1 _31154_ (.Y(_08492_),
    .A(net4530),
    .B(net7749));
 sg13g2_nand2_1 _31155_ (.Y(_08493_),
    .A(_07987_),
    .B(_07989_));
 sg13g2_nor2_1 _31156_ (.A(net8985),
    .B(_07990_),
    .Y(_08494_));
 sg13g2_xor2_1 _31157_ (.B(_08139_),
    .A(net4530),
    .X(_08495_));
 sg13g2_a22oi_1 _31158_ (.Y(_08496_),
    .B1(_08495_),
    .B2(net9215),
    .A2(_08494_),
    .A1(_08493_));
 sg13g2_o21ai_1 _31159_ (.B1(_08492_),
    .Y(_02202_),
    .A1(net7690),
    .A2(_08496_));
 sg13g2_nand2_1 _31160_ (.Y(_08497_),
    .A(net3229),
    .B(net7751));
 sg13g2_a21oi_1 _31161_ (.A1(net3229),
    .A2(_08138_),
    .Y(_08498_),
    .B1(net9078));
 sg13g2_xnor2_1 _31162_ (.Y(_08499_),
    .A(_07984_),
    .B(_07986_));
 sg13g2_nor2_1 _31163_ (.A(net8985),
    .B(_08499_),
    .Y(_08500_));
 sg13g2_a21oi_1 _31164_ (.A1(_08139_),
    .A2(_08498_),
    .Y(_08501_),
    .B1(_08500_));
 sg13g2_o21ai_1 _31165_ (.B1(_08497_),
    .Y(_02203_),
    .A1(net7690),
    .A2(_08501_));
 sg13g2_nand2_1 _31166_ (.Y(_08502_),
    .A(_07979_),
    .B(_07981_));
 sg13g2_nor2_1 _31167_ (.A(net8984),
    .B(_07982_),
    .Y(_08503_));
 sg13g2_xnor2_1 _31168_ (.Y(_08504_),
    .A(_10622_),
    .B(_08137_));
 sg13g2_a221oi_1 _31169_ (.B2(net9217),
    .C1(net7751),
    .B1(_08504_),
    .A1(_08502_),
    .Y(_08505_),
    .A2(_08503_));
 sg13g2_a21oi_1 _31170_ (.A1(_10622_),
    .A2(net7751),
    .Y(_02204_),
    .B1(_08505_));
 sg13g2_xnor2_1 _31171_ (.Y(_08506_),
    .A(_07976_),
    .B(_07978_));
 sg13g2_xnor2_1 _31172_ (.Y(_08507_),
    .A(net5214),
    .B(_08136_));
 sg13g2_a221oi_1 _31173_ (.B2(net9217),
    .C1(net7751),
    .B1(_08507_),
    .A1(net9209),
    .Y(_08508_),
    .A2(_08506_));
 sg13g2_a21oi_1 _31174_ (.A1(_10621_),
    .A2(net7751),
    .Y(_02205_),
    .B1(_08508_));
 sg13g2_nand2_1 _31175_ (.Y(_08509_),
    .A(_07971_),
    .B(_07973_));
 sg13g2_nand3_1 _31176_ (.B(_07974_),
    .C(_08509_),
    .A(net9209),
    .Y(_08510_));
 sg13g2_o21ai_1 _31177_ (.B1(net5201),
    .Y(_08511_),
    .A1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[0] ),
    .A2(net5066));
 sg13g2_nor2_1 _31178_ (.A(net9078),
    .B(_08136_),
    .Y(_08512_));
 sg13g2_a21oi_1 _31179_ (.A1(_08511_),
    .A2(_08512_),
    .Y(_08513_),
    .B1(net7751));
 sg13g2_a22oi_1 _31180_ (.Y(_02206_),
    .B1(_08510_),
    .B2(_08513_),
    .A2(net7751),
    .A1(_10620_));
 sg13g2_xor2_1 _31181_ (.B(_07970_),
    .A(_07968_),
    .X(_08514_));
 sg13g2_xor2_1 _31182_ (.B(net5066),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[0] ),
    .X(_08515_));
 sg13g2_a221oi_1 _31183_ (.B2(net9217),
    .C1(net7751),
    .B1(_08515_),
    .A1(net9209),
    .Y(_08516_),
    .A2(_08514_));
 sg13g2_a21oi_1 _31184_ (.A1(_10619_),
    .A2(net7749),
    .Y(_02207_),
    .B1(_08516_));
 sg13g2_o21ai_1 _31185_ (.B1(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[0] ),
    .Y(_08517_),
    .A1(net9217),
    .A2(_07479_));
 sg13g2_xnor2_1 _31186_ (.Y(_08518_),
    .A(net4491),
    .B(_07967_));
 sg13g2_o21ai_1 _31187_ (.B1(_08517_),
    .Y(_02208_),
    .A1(_08180_),
    .A2(_08518_));
 sg13g2_o21ai_1 _31188_ (.B1(net8494),
    .Y(_08519_),
    .A1(_10646_),
    .A2(net8373));
 sg13g2_nand2b_2 _31189_ (.Y(_08520_),
    .B(_08519_),
    .A_N(_13303_));
 sg13g2_nand4_1 _31190_ (.B(net9425),
    .C(net9427),
    .A(net9423),
    .Y(_08521_),
    .D(_10891_));
 sg13g2_and4_1 _31191_ (.A(_10894_),
    .B(_10896_),
    .C(_10934_),
    .D(_08521_),
    .X(_08522_));
 sg13g2_nand2_1 _31192_ (.Y(_08523_),
    .A(net9406),
    .B(net8846));
 sg13g2_a21oi_2 _31193_ (.B1(_08523_),
    .Y(_08524_),
    .A2(_08522_),
    .A1(_10936_));
 sg13g2_nor3_2 _31194_ (.A(net9294),
    .B(_10903_),
    .C(net8842),
    .Y(_08525_));
 sg13g2_nor3_1 _31195_ (.A(net9294),
    .B(_10971_),
    .C(_11012_),
    .Y(_08526_));
 sg13g2_nor3_1 _31196_ (.A(_08524_),
    .B(_08525_),
    .C(_08526_),
    .Y(_08527_));
 sg13g2_a22oi_1 _31197_ (.Y(_08528_),
    .B1(_13835_),
    .B2(\soc_I.clint_I.addr[0] ),
    .A2(\soc_I.clint_I.addr[1] ),
    .A1(net9705));
 sg13g2_or3_1 _31198_ (.A(net9051),
    .B(_10975_),
    .C(_08528_),
    .X(_08529_));
 sg13g2_o21ai_1 _31199_ (.B1(_08529_),
    .Y(_08530_),
    .A1(_08520_),
    .A2(_08527_));
 sg13g2_nand3b_1 _31200_ (.B(net8846),
    .C(net9001),
    .Y(_08531_),
    .A_N(_10905_));
 sg13g2_nand2_1 _31201_ (.Y(_08532_),
    .A(net9398),
    .B(_11055_));
 sg13g2_or2_1 _31202_ (.X(_08533_),
    .B(_08532_),
    .A(_10971_));
 sg13g2_a21oi_1 _31203_ (.A1(_08531_),
    .A2(_08533_),
    .Y(_08534_),
    .B1(_08528_));
 sg13g2_and3_1 _31204_ (.X(_08535_),
    .A(net9398),
    .B(_10969_),
    .C(_03849_));
 sg13g2_nor2_1 _31205_ (.A(net9444),
    .B(net9462),
    .Y(_08536_));
 sg13g2_or2_2 _31206_ (.X(_08537_),
    .B(net9471),
    .A(net9446));
 sg13g2_nor3_1 _31207_ (.A(net9423),
    .B(net9434),
    .C(net9708),
    .Y(_08538_));
 sg13g2_nand4_1 _31208_ (.B(_10924_),
    .C(_12584_),
    .A(\soc_I.kianv_I.Instr[6] ),
    .Y(_08539_),
    .D(_08538_));
 sg13g2_nor4_2 _31209_ (.A(_11000_),
    .B(_12609_),
    .C(net8594),
    .Y(_08540_),
    .D(_08539_));
 sg13g2_nand4_1 _31210_ (.B(_10906_),
    .C(net8923),
    .A(net9160),
    .Y(_08541_),
    .D(_08540_));
 sg13g2_nor2b_2 _31211_ (.A(net9446),
    .B_N(net9470),
    .Y(_08542_));
 sg13g2_nand2b_1 _31212_ (.Y(_08543_),
    .B(net9470),
    .A_N(net9446));
 sg13g2_nor2_2 _31213_ (.A(net9496),
    .B(net9141),
    .Y(_08544_));
 sg13g2_nand4_1 _31214_ (.B(_10458_),
    .C(_10895_),
    .A(\soc_I.kianv_I.Instr[28] ),
    .Y(_08545_),
    .D(net8766));
 sg13g2_nor2_1 _31215_ (.A(net8909),
    .B(_08545_),
    .Y(_08546_));
 sg13g2_nand3_1 _31216_ (.B(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[3] ),
    .C(\soc_I.kianv_I.control_unit_I.main_fsm_I.mip[3] ),
    .A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[3] ),
    .Y(_08547_));
 sg13g2_nand2_2 _31217_ (.Y(_08548_),
    .A(_04085_),
    .B(_08547_));
 sg13g2_nor3_2 _31218_ (.A(net9294),
    .B(_10981_),
    .C(_08548_),
    .Y(_08549_));
 sg13g2_and2_1 _31219_ (.A(_11011_),
    .B(_08549_),
    .X(_08550_));
 sg13g2_nor2_2 _31220_ (.A(net9712),
    .B(_11000_),
    .Y(_08551_));
 sg13g2_nand2_1 _31221_ (.Y(_08552_),
    .A(\soc_I.kianv_I.Instr[25] ),
    .B(_08551_));
 sg13g2_o21ai_1 _31222_ (.B1(_08551_),
    .Y(_08553_),
    .A1(\soc_I.kianv_I.Instr[25] ),
    .A2(_00285_));
 sg13g2_and2_1 _31223_ (.A(_08549_),
    .B(_08552_),
    .X(_08554_));
 sg13g2_and2_2 _31224_ (.A(_08550_),
    .B(_08553_),
    .X(_08555_));
 sg13g2_inv_1 _31225_ (.Y(_08556_),
    .A(_08555_));
 sg13g2_a21oi_1 _31226_ (.A1(_08540_),
    .A2(_08546_),
    .Y(_08557_),
    .B1(_08556_));
 sg13g2_nand3_1 _31227_ (.B(net9487),
    .C(_10893_),
    .A(net9430),
    .Y(_08558_));
 sg13g2_nor3_2 _31228_ (.A(net9522),
    .B(net8918),
    .C(_08558_),
    .Y(_08559_));
 sg13g2_nand2_1 _31229_ (.Y(_08560_),
    .A(_08540_),
    .B(_08559_));
 sg13g2_nor3_1 _31230_ (.A(_00214_),
    .B(_11005_),
    .C(_13291_),
    .Y(_08561_));
 sg13g2_nand2b_1 _31231_ (.Y(_08562_),
    .B(_11008_),
    .A_N(_08561_));
 sg13g2_nor4_1 _31232_ (.A(net9712),
    .B(net9713),
    .C(net9715),
    .D(_13291_),
    .Y(_08563_));
 sg13g2_nor4_1 _31233_ (.A(_11065_),
    .B(_13292_),
    .C(_08562_),
    .D(_08563_),
    .Y(_08564_));
 sg13g2_and3_1 _31234_ (.X(_08565_),
    .A(_10906_),
    .B(net8923),
    .C(_08540_));
 sg13g2_nand4_1 _31235_ (.B(_08557_),
    .C(_08560_),
    .A(_08541_),
    .Y(_08566_),
    .D(_08564_));
 sg13g2_nand2_1 _31236_ (.Y(_08567_),
    .A(net9398),
    .B(_03810_));
 sg13g2_nand3_1 _31237_ (.B(_08557_),
    .C(_08565_),
    .A(net8764),
    .Y(_08568_));
 sg13g2_o21ai_1 _31238_ (.B1(_08568_),
    .Y(_08569_),
    .A1(_11753_),
    .A2(_08567_));
 sg13g2_nor3_2 _31239_ (.A(net9295),
    .B(_10843_),
    .C(_03811_),
    .Y(_08570_));
 sg13g2_nor2_1 _31240_ (.A(net9296),
    .B(_03809_),
    .Y(_08571_));
 sg13g2_a21oi_1 _31241_ (.A1(net9398),
    .A2(net8673),
    .Y(_08572_),
    .B1(_08571_));
 sg13g2_inv_1 _31242_ (.Y(_08573_),
    .A(_08572_));
 sg13g2_nand3_1 _31243_ (.B(_10980_),
    .C(_08548_),
    .A(net9403),
    .Y(_08574_));
 sg13g2_nor2_1 _31244_ (.A(net9295),
    .B(_03821_),
    .Y(_08575_));
 sg13g2_nor2_1 _31245_ (.A(net9295),
    .B(_03816_),
    .Y(_08576_));
 sg13g2_a21oi_1 _31246_ (.A1(_03812_),
    .A2(_03816_),
    .Y(_08577_),
    .B1(net9294));
 sg13g2_nor2b_1 _31247_ (.A(_08577_),
    .B_N(_08574_),
    .Y(_08578_));
 sg13g2_nor4_2 _31248_ (.A(net9200),
    .B(net9296),
    .C(_10861_),
    .Y(_08579_),
    .D(_03811_));
 sg13g2_nor4_1 _31249_ (.A(_08570_),
    .B(_08573_),
    .C(_08575_),
    .D(_08579_),
    .Y(_08580_));
 sg13g2_nor2_1 _31250_ (.A(net9499),
    .B(net9536),
    .Y(_08581_));
 sg13g2_nand3_1 _31251_ (.B(_08565_),
    .C(net8875),
    .A(_08555_),
    .Y(_08582_));
 sg13g2_nand4_1 _31252_ (.B(_08578_),
    .C(_08580_),
    .A(_08566_),
    .Y(_08583_),
    .D(_08582_));
 sg13g2_nor4_1 _31253_ (.A(_08534_),
    .B(_08535_),
    .C(_08569_),
    .D(_08583_),
    .Y(_08584_));
 sg13g2_nand2b_1 _31254_ (.Y(_02209_),
    .B(_08584_),
    .A_N(_08530_));
 sg13g2_o21ai_1 _31255_ (.B1(_10602_),
    .Y(_08585_),
    .A1(_10596_),
    .A2(_13283_));
 sg13g2_nor3_1 _31256_ (.A(_10851_),
    .B(net8859),
    .C(_05887_),
    .Y(_08586_));
 sg13g2_and2_1 _31257_ (.A(net7472),
    .B(_08528_),
    .X(_08587_));
 sg13g2_inv_2 _31258_ (.Y(_08588_),
    .A(_08587_));
 sg13g2_nor3_2 _31259_ (.A(_10905_),
    .B(_08523_),
    .C(_08588_),
    .Y(_08589_));
 sg13g2_nor2b_1 _31260_ (.A(net4795),
    .B_N(_08589_),
    .Y(_08590_));
 sg13g2_nor3_1 _31261_ (.A(net9294),
    .B(_10970_),
    .C(_03849_),
    .Y(_08591_));
 sg13g2_nand4_1 _31262_ (.B(_10985_),
    .C(_03809_),
    .A(_10865_),
    .Y(_08592_),
    .D(_04252_));
 sg13g2_nor2_1 _31263_ (.A(net9294),
    .B(_10985_),
    .Y(_08593_));
 sg13g2_nor2_1 _31264_ (.A(net9295),
    .B(_10865_),
    .Y(_08594_));
 sg13g2_a22oi_1 _31265_ (.Y(_08595_),
    .B1(_08592_),
    .B2(_10602_),
    .A2(_08555_),
    .A1(_11004_));
 sg13g2_nand3_1 _31266_ (.B(_08557_),
    .C(_08559_),
    .A(_08540_),
    .Y(_08596_));
 sg13g2_or3_1 _31267_ (.A(_13293_),
    .B(_08556_),
    .C(_08562_),
    .X(_08597_));
 sg13g2_nand3_1 _31268_ (.B(_08596_),
    .C(_08597_),
    .A(_08595_),
    .Y(_08598_));
 sg13g2_nor3_2 _31269_ (.A(net9045),
    .B(_10596_),
    .C(_13283_),
    .Y(_08599_));
 sg13g2_nor2_1 _31270_ (.A(net9295),
    .B(_10975_),
    .Y(_08600_));
 sg13g2_a22oi_1 _31271_ (.Y(_08601_),
    .B1(_08600_),
    .B2(_08528_),
    .A2(_08599_),
    .A1(net8743));
 sg13g2_o21ai_1 _31272_ (.B1(_08601_),
    .Y(_08602_),
    .A1(_08585_),
    .A2(_08586_));
 sg13g2_nor4_1 _31273_ (.A(_08590_),
    .B(_08591_),
    .C(_08598_),
    .D(_08602_),
    .Y(_08603_));
 sg13g2_a22oi_1 _31274_ (.Y(_08604_),
    .B1(_08599_),
    .B2(_10851_),
    .A2(_08589_),
    .A1(net4795));
 sg13g2_nor2b_1 _31275_ (.A(net7483),
    .B_N(_08520_),
    .Y(_08605_));
 sg13g2_and2_1 _31276_ (.A(_08524_),
    .B(_08605_),
    .X(_08606_));
 sg13g2_a21o_1 _31277_ (.A2(_08599_),
    .A1(net8859),
    .B1(_08606_),
    .X(_08607_));
 sg13g2_a221oi_1 _31278_ (.B2(_08525_),
    .C1(_08607_),
    .B1(_08605_),
    .A1(_05887_),
    .Y(_08608_),
    .A2(_08599_));
 sg13g2_nand3_1 _31279_ (.B(_08604_),
    .C(_08608_),
    .A(_08603_),
    .Y(_02210_));
 sg13g2_nand2_1 _31280_ (.Y(_08609_),
    .A(_11062_),
    .B(_08554_));
 sg13g2_nand2_1 _31281_ (.Y(_08610_),
    .A(_08601_),
    .B(_08609_));
 sg13g2_nor2_1 _31282_ (.A(_08534_),
    .B(_08610_),
    .Y(_08611_));
 sg13g2_nor2_1 _31283_ (.A(_10855_),
    .B(_08585_),
    .Y(_08612_));
 sg13g2_or2_1 _31284_ (.X(_08613_),
    .B(_08612_),
    .A(_08576_));
 sg13g2_nand3b_1 _31285_ (.B(_08550_),
    .C(_08551_),
    .Y(_08614_),
    .A_N(_00285_));
 sg13g2_nor2_2 _31286_ (.A(\soc_I.kianv_I.control_unit_I.mul_ready ),
    .B(\soc_I.kianv_I.control_unit_I.div_ready ),
    .Y(_08615_));
 sg13g2_nand3_1 _31287_ (.B(_13831_),
    .C(_08615_),
    .A(net9398),
    .Y(_08616_));
 sg13g2_nand3_1 _31288_ (.B(_08614_),
    .C(_08616_),
    .A(_08596_),
    .Y(_08617_));
 sg13g2_nor3_1 _31289_ (.A(_08530_),
    .B(_08593_),
    .C(_08617_),
    .Y(_08618_));
 sg13g2_nand2b_1 _31290_ (.Y(_08619_),
    .B(_13831_),
    .A_N(_08615_));
 sg13g2_a21oi_1 _31291_ (.A1(_13830_),
    .A2(_03810_),
    .Y(_08620_),
    .B1(net8807));
 sg13g2_a21oi_1 _31292_ (.A1(_08619_),
    .A2(_08620_),
    .Y(_08621_),
    .B1(net9294));
 sg13g2_nand2_1 _31293_ (.Y(_08622_),
    .A(_10957_),
    .B(_08550_));
 sg13g2_inv_1 _31294_ (.Y(_08623_),
    .A(_08622_));
 sg13g2_nand2_1 _31295_ (.Y(_08624_),
    .A(_08550_),
    .B(_08561_));
 sg13g2_o21ai_1 _31296_ (.B1(_08624_),
    .Y(_08625_),
    .A1(net9294),
    .A2(_10968_));
 sg13g2_nand3_1 _31297_ (.B(_11006_),
    .C(_08555_),
    .A(_10955_),
    .Y(_08626_));
 sg13g2_nand3b_1 _31298_ (.B(_11006_),
    .C(_08555_),
    .Y(_08627_),
    .A_N(_10954_));
 sg13g2_nor4_1 _31299_ (.A(_08594_),
    .B(_08621_),
    .C(_08623_),
    .D(_08625_),
    .Y(_08628_));
 sg13g2_o21ai_1 _31300_ (.B1(_08628_),
    .Y(_08629_),
    .A1(net9295),
    .A2(_03814_));
 sg13g2_a21oi_1 _31301_ (.A1(_11007_),
    .A2(_08554_),
    .Y(_08630_),
    .B1(_08629_));
 sg13g2_nand4_1 _31302_ (.B(_08618_),
    .C(_08627_),
    .A(_08566_),
    .Y(_08631_),
    .D(_08630_));
 sg13g2_nor3_1 _31303_ (.A(_08607_),
    .B(_08613_),
    .C(_08631_),
    .Y(_08632_));
 sg13g2_nand2_1 _31304_ (.Y(_02211_),
    .A(_08611_),
    .B(_08632_));
 sg13g2_nor4_1 _31305_ (.A(net9051),
    .B(_10981_),
    .C(_11010_),
    .D(_08548_),
    .Y(_08633_));
 sg13g2_nand3_1 _31306_ (.B(_08551_),
    .C(_08633_),
    .A(_00285_),
    .Y(_08634_));
 sg13g2_o21ai_1 _31307_ (.B1(_08634_),
    .Y(_08635_),
    .A1(_10852_),
    .A2(_08585_));
 sg13g2_a21oi_1 _31308_ (.A1(_10837_),
    .A2(_08599_),
    .Y(_08636_),
    .B1(_08575_));
 sg13g2_o21ai_1 _31309_ (.B1(_08636_),
    .Y(_08637_),
    .A1(_08533_),
    .A2(_08588_));
 sg13g2_nor4_1 _31310_ (.A(net9204),
    .B(_10847_),
    .C(_10849_),
    .D(_08585_),
    .Y(_08638_));
 sg13g2_nor2_1 _31311_ (.A(_08569_),
    .B(_08590_),
    .Y(_08639_));
 sg13g2_a21oi_1 _31312_ (.A1(_10884_),
    .A2(_10887_),
    .Y(_08640_),
    .B1(net9051));
 sg13g2_nor4_1 _31313_ (.A(_08570_),
    .B(_08617_),
    .C(_08621_),
    .D(_08640_),
    .Y(_08641_));
 sg13g2_nand3_1 _31314_ (.B(_08639_),
    .C(_08641_),
    .A(_08574_),
    .Y(_08642_));
 sg13g2_nor4_1 _31315_ (.A(_08635_),
    .B(_08637_),
    .C(_08638_),
    .D(_08642_),
    .Y(_08643_));
 sg13g2_and2_1 _31316_ (.A(_08604_),
    .B(_08622_),
    .X(_08644_));
 sg13g2_nand3_1 _31317_ (.B(_08643_),
    .C(_08644_),
    .A(_08611_),
    .Y(_02212_));
 sg13g2_nor4_1 _31318_ (.A(_08579_),
    .B(_08594_),
    .C(_08621_),
    .D(_08640_),
    .Y(_08645_));
 sg13g2_nand2_1 _31319_ (.Y(_08646_),
    .A(_08526_),
    .B(_08605_));
 sg13g2_nand4_1 _31320_ (.B(_08639_),
    .C(_08645_),
    .A(_08626_),
    .Y(_08647_),
    .D(_08646_));
 sg13g2_a221oi_1 _31321_ (.B2(_08525_),
    .C1(_08647_),
    .B1(_08605_),
    .A1(_10850_),
    .Y(_08648_),
    .A2(_08599_));
 sg13g2_a22oi_1 _31322_ (.Y(_08649_),
    .B1(_08555_),
    .B2(_11056_),
    .A2(_08549_),
    .A1(_11010_));
 sg13g2_nand4_1 _31323_ (.B(_08597_),
    .C(_08618_),
    .A(_08582_),
    .Y(_08650_),
    .D(_08649_));
 sg13g2_nor2_1 _31324_ (.A(_08635_),
    .B(_08650_),
    .Y(_08651_));
 sg13g2_nand2_1 _31325_ (.Y(_02213_),
    .A(_08648_),
    .B(_08651_));
 sg13g2_nor4_1 _31326_ (.A(_08570_),
    .B(_08573_),
    .C(_08591_),
    .D(_08625_),
    .Y(_08652_));
 sg13g2_o21ai_1 _31327_ (.B1(_08652_),
    .Y(_08653_),
    .A1(net9295),
    .A2(net7374));
 sg13g2_nor3_1 _31328_ (.A(_08613_),
    .B(_08637_),
    .C(_08653_),
    .Y(_08654_));
 sg13g2_nand3_1 _31329_ (.B(_08648_),
    .C(_08654_),
    .A(_08644_),
    .Y(_02214_));
 sg13g2_nand2_1 _31330_ (.Y(_08655_),
    .A(_14199_),
    .B(_14370_));
 sg13g2_nand2_1 _31331_ (.Y(_08656_),
    .A(net3708),
    .B(net7864));
 sg13g2_o21ai_1 _31332_ (.B1(_08656_),
    .Y(_02215_),
    .A1(net7486),
    .A2(net7864));
 sg13g2_nand2_1 _31333_ (.Y(_08657_),
    .A(net2882),
    .B(net7861));
 sg13g2_o21ai_1 _31334_ (.B1(_08657_),
    .Y(_02216_),
    .A1(net7666),
    .A2(net7861));
 sg13g2_nand2_1 _31335_ (.Y(_08658_),
    .A(net3614),
    .B(net7861));
 sg13g2_o21ai_1 _31336_ (.B1(_08658_),
    .Y(_02217_),
    .A1(net7614),
    .A2(net7861));
 sg13g2_nand2_1 _31337_ (.Y(_08659_),
    .A(net3101),
    .B(net7862));
 sg13g2_o21ai_1 _31338_ (.B1(_08659_),
    .Y(_02218_),
    .A1(net7607),
    .A2(net7862));
 sg13g2_nand2_1 _31339_ (.Y(_08660_),
    .A(net4072),
    .B(net7864));
 sg13g2_o21ai_1 _31340_ (.B1(_08660_),
    .Y(_02219_),
    .A1(net7589),
    .A2(net7864));
 sg13g2_nand2_1 _31341_ (.Y(_08661_),
    .A(net2982),
    .B(net7865));
 sg13g2_o21ai_1 _31342_ (.B1(_08661_),
    .Y(_02220_),
    .A1(net7599),
    .A2(net7865));
 sg13g2_nand2_1 _31343_ (.Y(_08662_),
    .A(net3573),
    .B(net7863));
 sg13g2_o21ai_1 _31344_ (.B1(_08662_),
    .Y(_02221_),
    .A1(net7592),
    .A2(net7863));
 sg13g2_nand2_1 _31345_ (.Y(_08663_),
    .A(net4191),
    .B(net7857));
 sg13g2_o21ai_1 _31346_ (.B1(_08663_),
    .Y(_02222_),
    .A1(net7606),
    .A2(net7857));
 sg13g2_nand2_1 _31347_ (.Y(_08664_),
    .A(net3641),
    .B(net7865));
 sg13g2_o21ai_1 _31348_ (.B1(_08664_),
    .Y(_02223_),
    .A1(net7560),
    .A2(net7865));
 sg13g2_nand2_1 _31349_ (.Y(_08665_),
    .A(net3501),
    .B(net7863));
 sg13g2_o21ai_1 _31350_ (.B1(_08665_),
    .Y(_02224_),
    .A1(net7574),
    .A2(net7863));
 sg13g2_nand2_1 _31351_ (.Y(_08666_),
    .A(net3204),
    .B(net7862));
 sg13g2_o21ai_1 _31352_ (.B1(_08666_),
    .Y(_02225_),
    .A1(net7547),
    .A2(net7862));
 sg13g2_nand2_1 _31353_ (.Y(_08667_),
    .A(net3873),
    .B(net7857));
 sg13g2_o21ai_1 _31354_ (.B1(_08667_),
    .Y(_02226_),
    .A1(net7573),
    .A2(net7857));
 sg13g2_nand2_1 _31355_ (.Y(_08668_),
    .A(net3841),
    .B(net7863));
 sg13g2_o21ai_1 _31356_ (.B1(_08668_),
    .Y(_02227_),
    .A1(net7540),
    .A2(net7863));
 sg13g2_nand2_1 _31357_ (.Y(_08669_),
    .A(net3771),
    .B(net7863));
 sg13g2_o21ai_1 _31358_ (.B1(_08669_),
    .Y(_02228_),
    .A1(net7551),
    .A2(net7863));
 sg13g2_nand2_1 _31359_ (.Y(_08670_),
    .A(net3714),
    .B(net7859));
 sg13g2_o21ai_1 _31360_ (.B1(_08670_),
    .Y(_02229_),
    .A1(net7583),
    .A2(net7859));
 sg13g2_nand2_1 _31361_ (.Y(_08671_),
    .A(net3144),
    .B(net7858));
 sg13g2_o21ai_1 _31362_ (.B1(_08671_),
    .Y(_02230_),
    .A1(net7565),
    .A2(net7859));
 sg13g2_nand2_1 _31363_ (.Y(_08672_),
    .A(net3958),
    .B(net7857));
 sg13g2_o21ai_1 _31364_ (.B1(_08672_),
    .Y(_02231_),
    .A1(net7526),
    .A2(net7857));
 sg13g2_nand2_1 _31365_ (.Y(_08673_),
    .A(net3648),
    .B(net7857));
 sg13g2_o21ai_1 _31366_ (.B1(_08673_),
    .Y(_02232_),
    .A1(net7539),
    .A2(net7857));
 sg13g2_nand2_1 _31367_ (.Y(_08674_),
    .A(net3100),
    .B(net7858));
 sg13g2_o21ai_1 _31368_ (.B1(_08674_),
    .Y(_02233_),
    .A1(net7530),
    .A2(net7858));
 sg13g2_nand2_1 _31369_ (.Y(_08675_),
    .A(net3036),
    .B(net7859));
 sg13g2_o21ai_1 _31370_ (.B1(_08675_),
    .Y(_02234_),
    .A1(net7516),
    .A2(net7859));
 sg13g2_nand2_1 _31371_ (.Y(_08676_),
    .A(net3851),
    .B(net7864));
 sg13g2_o21ai_1 _31372_ (.B1(_08676_),
    .Y(_02235_),
    .A1(net7506),
    .A2(net7864));
 sg13g2_nand2_1 _31373_ (.Y(_08677_),
    .A(net3078),
    .B(net7860));
 sg13g2_o21ai_1 _31374_ (.B1(_08677_),
    .Y(_02236_),
    .A1(net7511),
    .A2(net7860));
 sg13g2_nand2_1 _31375_ (.Y(_08678_),
    .A(net3003),
    .B(net7861));
 sg13g2_o21ai_1 _31376_ (.B1(_08678_),
    .Y(_02237_),
    .A1(net7497),
    .A2(net7861));
 sg13g2_nand2_1 _31377_ (.Y(_08679_),
    .A(net3202),
    .B(net7858));
 sg13g2_o21ai_1 _31378_ (.B1(_08679_),
    .Y(_02238_),
    .A1(net7501),
    .A2(net7858));
 sg13g2_nand2_1 _31379_ (.Y(_08680_),
    .A(net3275),
    .B(net7865));
 sg13g2_o21ai_1 _31380_ (.B1(_08680_),
    .Y(_02239_),
    .A1(net7645),
    .A2(net7865));
 sg13g2_nand2_1 _31381_ (.Y(_08681_),
    .A(net3541),
    .B(net7864));
 sg13g2_o21ai_1 _31382_ (.B1(_08681_),
    .Y(_02240_),
    .A1(net7651),
    .A2(net7864));
 sg13g2_nand2_1 _31383_ (.Y(_08682_),
    .A(net3027),
    .B(net7861));
 sg13g2_o21ai_1 _31384_ (.B1(_08682_),
    .Y(_02241_),
    .A1(net7653),
    .A2(net7861));
 sg13g2_nand2_1 _31385_ (.Y(_08683_),
    .A(net3482),
    .B(net7860));
 sg13g2_o21ai_1 _31386_ (.B1(_08683_),
    .Y(_02242_),
    .A1(net7660),
    .A2(net7860));
 sg13g2_nand2_1 _31387_ (.Y(_08684_),
    .A(net3129),
    .B(net7860));
 sg13g2_o21ai_1 _31388_ (.B1(_08684_),
    .Y(_02243_),
    .A1(net7636),
    .A2(net7860));
 sg13g2_nand2_1 _31389_ (.Y(_08685_),
    .A(net3220),
    .B(net7865));
 sg13g2_o21ai_1 _31390_ (.B1(_08685_),
    .Y(_02244_),
    .A1(net7626),
    .A2(net7865));
 sg13g2_nand2_1 _31391_ (.Y(_08686_),
    .A(net3936),
    .B(net7867));
 sg13g2_o21ai_1 _31392_ (.B1(_08686_),
    .Y(_02245_),
    .A1(net7620),
    .A2(net7860));
 sg13g2_nand2_1 _31393_ (.Y(_08687_),
    .A(net3050),
    .B(net7858));
 sg13g2_o21ai_1 _31394_ (.B1(_08687_),
    .Y(_02246_),
    .A1(net7632),
    .A2(net7858));
 sg13g2_nand2_1 _31395_ (.Y(_08688_),
    .A(_14301_),
    .B(_14370_));
 sg13g2_nand2_1 _31396_ (.Y(_08689_),
    .A(net3329),
    .B(net7854));
 sg13g2_o21ai_1 _31397_ (.B1(_08689_),
    .Y(_02247_),
    .A1(net7486),
    .A2(net7854));
 sg13g2_nand2_1 _31398_ (.Y(_08690_),
    .A(net3874),
    .B(net7851));
 sg13g2_o21ai_1 _31399_ (.B1(_08690_),
    .Y(_02248_),
    .A1(net7664),
    .A2(net7851));
 sg13g2_nand2_1 _31400_ (.Y(_08691_),
    .A(net3434),
    .B(net7853));
 sg13g2_o21ai_1 _31401_ (.B1(_08691_),
    .Y(_02249_),
    .A1(net7614),
    .A2(net7853));
 sg13g2_nand2_1 _31402_ (.Y(_08692_),
    .A(net3813),
    .B(net7852));
 sg13g2_o21ai_1 _31403_ (.B1(_08692_),
    .Y(_02250_),
    .A1(net7608),
    .A2(net7852));
 sg13g2_nand2_1 _31404_ (.Y(_08693_),
    .A(net3790),
    .B(net7854));
 sg13g2_o21ai_1 _31405_ (.B1(_08693_),
    .Y(_02251_),
    .A1(net7589),
    .A2(net7854));
 sg13g2_nand2_1 _31406_ (.Y(_08694_),
    .A(net3314),
    .B(net7855));
 sg13g2_o21ai_1 _31407_ (.B1(_08694_),
    .Y(_02252_),
    .A1(net7599),
    .A2(net7855));
 sg13g2_nand2_1 _31408_ (.Y(_08695_),
    .A(net3183),
    .B(net7852));
 sg13g2_o21ai_1 _31409_ (.B1(_08695_),
    .Y(_02253_),
    .A1(net7592),
    .A2(net7852));
 sg13g2_nand2_1 _31410_ (.Y(_08696_),
    .A(net3094),
    .B(net7848));
 sg13g2_o21ai_1 _31411_ (.B1(_08696_),
    .Y(_02254_),
    .A1(net7604),
    .A2(net7848));
 sg13g2_nand2_1 _31412_ (.Y(_08697_),
    .A(net3491),
    .B(net7855));
 sg13g2_o21ai_1 _31413_ (.B1(_08697_),
    .Y(_02255_),
    .A1(net7558),
    .A2(net7855));
 sg13g2_nand2_1 _31414_ (.Y(_08698_),
    .A(net2861),
    .B(net7851));
 sg13g2_o21ai_1 _31415_ (.B1(_08698_),
    .Y(_02256_),
    .A1(net7574),
    .A2(net7851));
 sg13g2_nand2_1 _31416_ (.Y(_08699_),
    .A(net3850),
    .B(net7853));
 sg13g2_o21ai_1 _31417_ (.B1(_08699_),
    .Y(_02257_),
    .A1(net7547),
    .A2(net7853));
 sg13g2_nand2_1 _31418_ (.Y(_08700_),
    .A(net3564),
    .B(net7846));
 sg13g2_o21ai_1 _31419_ (.B1(_08700_),
    .Y(_02258_),
    .A1(net7573),
    .A2(net7846));
 sg13g2_nand2_1 _31420_ (.Y(_08701_),
    .A(net3235),
    .B(net7851));
 sg13g2_o21ai_1 _31421_ (.B1(_08701_),
    .Y(_02259_),
    .A1(net7542),
    .A2(net7851));
 sg13g2_nand2_1 _31422_ (.Y(_08702_),
    .A(net3397),
    .B(net7851));
 sg13g2_o21ai_1 _31423_ (.B1(_08702_),
    .Y(_02260_),
    .A1(net7551),
    .A2(net7851));
 sg13g2_nand2_1 _31424_ (.Y(_08703_),
    .A(net3741),
    .B(net7849));
 sg13g2_o21ai_1 _31425_ (.B1(_08703_),
    .Y(_02261_),
    .A1(net7583),
    .A2(net7849));
 sg13g2_nand2_1 _31426_ (.Y(_08704_),
    .A(net2895),
    .B(net7846));
 sg13g2_o21ai_1 _31427_ (.B1(_08704_),
    .Y(_02262_),
    .A1(net7565),
    .A2(net7846));
 sg13g2_nand2_1 _31428_ (.Y(_08705_),
    .A(net3021),
    .B(net7846));
 sg13g2_o21ai_1 _31429_ (.B1(_08705_),
    .Y(_02263_),
    .A1(net7526),
    .A2(net7846));
 sg13g2_nand2_1 _31430_ (.Y(_08706_),
    .A(net3666),
    .B(net7846));
 sg13g2_o21ai_1 _31431_ (.B1(_08706_),
    .Y(_02264_),
    .A1(net7538),
    .A2(net7846));
 sg13g2_nand2_1 _31432_ (.Y(_08707_),
    .A(net3549),
    .B(net7848));
 sg13g2_o21ai_1 _31433_ (.B1(_08707_),
    .Y(_02265_),
    .A1(net7530),
    .A2(net7848));
 sg13g2_nand2_1 _31434_ (.Y(_08708_),
    .A(net3132),
    .B(net7850));
 sg13g2_o21ai_1 _31435_ (.B1(_08708_),
    .Y(_02266_),
    .A1(net7516),
    .A2(net7848));
 sg13g2_nand2_1 _31436_ (.Y(_08709_),
    .A(net3699),
    .B(net7854));
 sg13g2_o21ai_1 _31437_ (.B1(_08709_),
    .Y(_02267_),
    .A1(net7506),
    .A2(net7854));
 sg13g2_nand2_1 _31438_ (.Y(_08710_),
    .A(net3428),
    .B(net7850));
 sg13g2_o21ai_1 _31439_ (.B1(_08710_),
    .Y(_02268_),
    .A1(net7511),
    .A2(net7850));
 sg13g2_nand2_1 _31440_ (.Y(_08711_),
    .A(net3017),
    .B(net7852));
 sg13g2_o21ai_1 _31441_ (.B1(_08711_),
    .Y(_02269_),
    .A1(net7494),
    .A2(net7852));
 sg13g2_nand2_1 _31442_ (.Y(_08712_),
    .A(net3739),
    .B(net7847));
 sg13g2_o21ai_1 _31443_ (.B1(_08712_),
    .Y(_02270_),
    .A1(net7501),
    .A2(net7847));
 sg13g2_nand2_1 _31444_ (.Y(_08713_),
    .A(net3242),
    .B(net7855));
 sg13g2_o21ai_1 _31445_ (.B1(_08713_),
    .Y(_02271_),
    .A1(net7642),
    .A2(net7855));
 sg13g2_nand2_1 _31446_ (.Y(_08714_),
    .A(net3031),
    .B(net7854));
 sg13g2_o21ai_1 _31447_ (.B1(_08714_),
    .Y(_02272_),
    .A1(net7651),
    .A2(net7854));
 sg13g2_nand2_1 _31448_ (.Y(_08715_),
    .A(net3876),
    .B(net7852));
 sg13g2_o21ai_1 _31449_ (.B1(_08715_),
    .Y(_02273_),
    .A1(net7657),
    .A2(net7852));
 sg13g2_nand2_1 _31450_ (.Y(_08716_),
    .A(net3815),
    .B(net7849));
 sg13g2_o21ai_1 _31451_ (.B1(_08716_),
    .Y(_02274_),
    .A1(net7659),
    .A2(net7849));
 sg13g2_nand2_1 _31452_ (.Y(_08717_),
    .A(net3452),
    .B(net7849));
 sg13g2_o21ai_1 _31453_ (.B1(_08717_),
    .Y(_02275_),
    .A1(net7636),
    .A2(net7849));
 sg13g2_nand2_1 _31454_ (.Y(_08718_),
    .A(net3480),
    .B(net7855));
 sg13g2_o21ai_1 _31455_ (.B1(_08718_),
    .Y(_02276_),
    .A1(net7626),
    .A2(net7855));
 sg13g2_nand2_1 _31456_ (.Y(_08719_),
    .A(net3861),
    .B(net7849));
 sg13g2_o21ai_1 _31457_ (.B1(_08719_),
    .Y(_02277_),
    .A1(net7619),
    .A2(net7849));
 sg13g2_nand2_1 _31458_ (.Y(_08720_),
    .A(net3338),
    .B(net7847));
 sg13g2_o21ai_1 _31459_ (.B1(_08720_),
    .Y(_02278_),
    .A1(net7632),
    .A2(net7847));
 sg13g2_nand2_1 _31460_ (.Y(_08721_),
    .A(net2642),
    .B(net8584));
 sg13g2_o21ai_1 _31461_ (.B1(_08721_),
    .Y(_02279_),
    .A1(net9170),
    .A2(net8584));
 sg13g2_mux2_1 _31462_ (.A0(net9288),
    .A1(net4211),
    .S(net8584),
    .X(_02280_));
 sg13g2_mux2_1 _31463_ (.A0(net9287),
    .A1(net4107),
    .S(net8584),
    .X(_02281_));
 sg13g2_mux2_1 _31464_ (.A0(net9284),
    .A1(net4254),
    .S(net8584),
    .X(_02282_));
 sg13g2_mux2_1 _31465_ (.A0(net9283),
    .A1(net4016),
    .S(_06952_),
    .X(_02283_));
 sg13g2_mux2_1 _31466_ (.A0(net9281),
    .A1(net4037),
    .S(net8584),
    .X(_02284_));
 sg13g2_mux2_1 _31467_ (.A0(net9277),
    .A1(net4106),
    .S(net8584),
    .X(_02285_));
 sg13g2_mux2_1 _31468_ (.A0(\soc_I.rx_uart_i.fifo_i.din[7] ),
    .A1(net4112),
    .S(net8584),
    .X(_02286_));
 sg13g2_nand2_1 _31469_ (.Y(_08722_),
    .A(_14123_),
    .B(_02801_));
 sg13g2_nand2_1 _31470_ (.Y(_08723_),
    .A(net2841),
    .B(net8530));
 sg13g2_o21ai_1 _31471_ (.B1(_08723_),
    .Y(_02287_),
    .A1(net9170),
    .A2(net8530));
 sg13g2_mux2_1 _31472_ (.A0(net9288),
    .A1(net4091),
    .S(net8530),
    .X(_02288_));
 sg13g2_mux2_1 _31473_ (.A0(net9287),
    .A1(net3956),
    .S(net8530),
    .X(_02289_));
 sg13g2_mux2_1 _31474_ (.A0(net9284),
    .A1(net4053),
    .S(net8530),
    .X(_02290_));
 sg13g2_mux2_1 _31475_ (.A0(net9283),
    .A1(net4010),
    .S(_08722_),
    .X(_02291_));
 sg13g2_mux2_1 _31476_ (.A0(net9281),
    .A1(net4014),
    .S(net8530),
    .X(_02292_));
 sg13g2_mux2_1 _31477_ (.A0(net9277),
    .A1(net4218),
    .S(net8530),
    .X(_02293_));
 sg13g2_mux2_1 _31478_ (.A0(net9276),
    .A1(net4318),
    .S(net8530),
    .X(_02294_));
 sg13g2_nand2_1 _31479_ (.Y(_08724_),
    .A(_14123_),
    .B(_02810_));
 sg13g2_nand2_1 _31480_ (.Y(_08725_),
    .A(net2708),
    .B(net8579));
 sg13g2_o21ai_1 _31481_ (.B1(_08725_),
    .Y(_02295_),
    .A1(net9170),
    .A2(net8579));
 sg13g2_mux2_1 _31482_ (.A0(net9288),
    .A1(net4198),
    .S(net8579),
    .X(_02296_));
 sg13g2_mux2_1 _31483_ (.A0(net9287),
    .A1(net4260),
    .S(net8579),
    .X(_02297_));
 sg13g2_mux2_1 _31484_ (.A0(net9284),
    .A1(net4547),
    .S(net8579),
    .X(_02298_));
 sg13g2_mux2_1 _31485_ (.A0(net9283),
    .A1(net4040),
    .S(_08724_),
    .X(_02299_));
 sg13g2_mux2_1 _31486_ (.A0(net9281),
    .A1(net3949),
    .S(net8579),
    .X(_02300_));
 sg13g2_mux2_1 _31487_ (.A0(net9277),
    .A1(net4101),
    .S(net8579),
    .X(_02301_));
 sg13g2_mux2_1 _31488_ (.A0(net9275),
    .A1(net4036),
    .S(net8579),
    .X(_02302_));
 sg13g2_nand4_1 _31489_ (.B(_14127_),
    .C(net8371),
    .A(net9710),
    .Y(_08726_),
    .D(_14199_));
 sg13g2_nand2_1 _31490_ (.Y(_08727_),
    .A(net3114),
    .B(net8070));
 sg13g2_o21ai_1 _31491_ (.B1(_08727_),
    .Y(_02303_),
    .A1(net7488),
    .A2(net8070));
 sg13g2_nand2_1 _31492_ (.Y(_08728_),
    .A(net3500),
    .B(net8074));
 sg13g2_o21ai_1 _31493_ (.B1(_08728_),
    .Y(_02304_),
    .A1(net7664),
    .A2(net8074));
 sg13g2_nand2_1 _31494_ (.Y(_08729_),
    .A(net3008),
    .B(net8070));
 sg13g2_o21ai_1 _31495_ (.B1(_08729_),
    .Y(_02305_),
    .A1(net7612),
    .A2(net8070));
 sg13g2_nand2_1 _31496_ (.Y(_08730_),
    .A(net3612),
    .B(net8072));
 sg13g2_o21ai_1 _31497_ (.B1(_08730_),
    .Y(_02306_),
    .A1(net7610),
    .A2(net8072));
 sg13g2_nand2_1 _31498_ (.Y(_08731_),
    .A(net3801),
    .B(net8070));
 sg13g2_o21ai_1 _31499_ (.B1(_08731_),
    .Y(_02307_),
    .A1(net7589),
    .A2(net8070));
 sg13g2_nand2_1 _31500_ (.Y(_08732_),
    .A(net3756),
    .B(net8068));
 sg13g2_o21ai_1 _31501_ (.B1(_08732_),
    .Y(_02308_),
    .A1(net7599),
    .A2(net8068));
 sg13g2_nand2_1 _31502_ (.Y(_08733_),
    .A(net3070),
    .B(net8071));
 sg13g2_o21ai_1 _31503_ (.B1(_08733_),
    .Y(_02309_),
    .A1(net7595),
    .A2(net8071));
 sg13g2_nand2_1 _31504_ (.Y(_08734_),
    .A(net3899),
    .B(net8064));
 sg13g2_o21ai_1 _31505_ (.B1(_08734_),
    .Y(_02310_),
    .A1(net7603),
    .A2(net8064));
 sg13g2_nand2_1 _31506_ (.Y(_08735_),
    .A(net2730),
    .B(net8069));
 sg13g2_o21ai_1 _31507_ (.B1(_08735_),
    .Y(_02311_),
    .A1(net7560),
    .A2(net8069));
 sg13g2_nand2_1 _31508_ (.Y(_08736_),
    .A(net3025),
    .B(net8073));
 sg13g2_o21ai_1 _31509_ (.B1(_08736_),
    .Y(_02312_),
    .A1(net7574),
    .A2(net8073));
 sg13g2_nand2_1 _31510_ (.Y(_08737_),
    .A(net3018),
    .B(net8072));
 sg13g2_o21ai_1 _31511_ (.B1(_08737_),
    .Y(_02313_),
    .A1(net7549),
    .A2(net8072));
 sg13g2_nand2_1 _31512_ (.Y(_08738_),
    .A(net3959),
    .B(net8064));
 sg13g2_o21ai_1 _31513_ (.B1(_08738_),
    .Y(_02314_),
    .A1(net7569),
    .A2(net8064));
 sg13g2_nand2_1 _31514_ (.Y(_08739_),
    .A(net3429),
    .B(net8071));
 sg13g2_o21ai_1 _31515_ (.B1(_08739_),
    .Y(_02315_),
    .A1(net7544),
    .A2(net8071));
 sg13g2_nand2_1 _31516_ (.Y(_08740_),
    .A(net3327),
    .B(net8073));
 sg13g2_o21ai_1 _31517_ (.B1(_08740_),
    .Y(_02316_),
    .A1(net7555),
    .A2(net8073));
 sg13g2_nand2_1 _31518_ (.Y(_08741_),
    .A(net3721),
    .B(net8066));
 sg13g2_o21ai_1 _31519_ (.B1(_08741_),
    .Y(_02317_),
    .A1(net7583),
    .A2(net8066));
 sg13g2_nand2_1 _31520_ (.Y(_08742_),
    .A(net3442),
    .B(net8065));
 sg13g2_o21ai_1 _31521_ (.B1(_08742_),
    .Y(_02318_),
    .A1(net7563),
    .A2(net8065));
 sg13g2_nand2_1 _31522_ (.Y(_08743_),
    .A(net3787),
    .B(net8064));
 sg13g2_o21ai_1 _31523_ (.B1(_08743_),
    .Y(_02319_),
    .A1(net7523),
    .A2(net8064));
 sg13g2_nand2_1 _31524_ (.Y(_08744_),
    .A(net3724),
    .B(net8064));
 sg13g2_o21ai_1 _31525_ (.B1(_08744_),
    .Y(_02320_),
    .A1(net7534),
    .A2(net8064));
 sg13g2_nand2_1 _31526_ (.Y(_08745_),
    .A(net3766),
    .B(net8065));
 sg13g2_o21ai_1 _31527_ (.B1(_08745_),
    .Y(_02321_),
    .A1(net7528),
    .A2(net8065));
 sg13g2_nand2_1 _31528_ (.Y(_08746_),
    .A(net3814),
    .B(net8066));
 sg13g2_o21ai_1 _31529_ (.B1(_08746_),
    .Y(_02322_),
    .A1(net7520),
    .A2(net8066));
 sg13g2_nand2_1 _31530_ (.Y(_08747_),
    .A(net3402),
    .B(net8070));
 sg13g2_o21ai_1 _31531_ (.B1(_08747_),
    .Y(_02323_),
    .A1(net7506),
    .A2(net8070));
 sg13g2_nand2_1 _31532_ (.Y(_08748_),
    .A(net3773),
    .B(net8068));
 sg13g2_o21ai_1 _31533_ (.B1(_08748_),
    .Y(_02324_),
    .A1(net7514),
    .A2(net8068));
 sg13g2_nand2_1 _31534_ (.Y(_08749_),
    .A(net3396),
    .B(net8071));
 sg13g2_o21ai_1 _31535_ (.B1(_08749_),
    .Y(_02325_),
    .A1(net7495),
    .A2(net8071));
 sg13g2_nand2_1 _31536_ (.Y(_08750_),
    .A(net3759),
    .B(net8065));
 sg13g2_o21ai_1 _31537_ (.B1(_08750_),
    .Y(_02326_),
    .A1(net7499),
    .A2(net8065));
 sg13g2_nand2_1 _31538_ (.Y(_08751_),
    .A(net3506),
    .B(net8068));
 sg13g2_o21ai_1 _31539_ (.B1(_08751_),
    .Y(_02327_),
    .A1(net7643),
    .A2(net8068));
 sg13g2_nand2_1 _31540_ (.Y(_08752_),
    .A(net3356),
    .B(net8068));
 sg13g2_o21ai_1 _31541_ (.B1(_08752_),
    .Y(_02328_),
    .A1(net7648),
    .A2(net8068));
 sg13g2_nand2_1 _31542_ (.Y(_08753_),
    .A(net3269),
    .B(net8071));
 sg13g2_o21ai_1 _31543_ (.B1(_08753_),
    .Y(_02329_),
    .A1(net7654),
    .A2(net8071));
 sg13g2_nand2_1 _31544_ (.Y(_08754_),
    .A(net4236),
    .B(net8066));
 sg13g2_o21ai_1 _31545_ (.B1(_08754_),
    .Y(_02330_),
    .A1(net7658),
    .A2(net8066));
 sg13g2_nand2_1 _31546_ (.Y(_08755_),
    .A(net3693),
    .B(net8066));
 sg13g2_o21ai_1 _31547_ (.B1(_08755_),
    .Y(_02331_),
    .A1(net7640),
    .A2(net8066));
 sg13g2_nand2_1 _31548_ (.Y(_08756_),
    .A(net3715),
    .B(net8069));
 sg13g2_o21ai_1 _31549_ (.B1(_08756_),
    .Y(_02332_),
    .A1(net7628),
    .A2(net8069));
 sg13g2_nand2_1 _31550_ (.Y(_08757_),
    .A(net4031),
    .B(net8067));
 sg13g2_o21ai_1 _31551_ (.B1(_08757_),
    .Y(_02333_),
    .A1(net7622),
    .A2(net8067));
 sg13g2_nand2_1 _31552_ (.Y(_08758_),
    .A(net3870),
    .B(net8067));
 sg13g2_o21ai_1 _31553_ (.B1(_08758_),
    .Y(_02334_),
    .A1(net7630),
    .A2(net8067));
 sg13g2_nand2_2 _31554_ (.Y(_08759_),
    .A(net8961),
    .B(_03742_));
 sg13g2_nand2_1 _31555_ (.Y(_08760_),
    .A(net3847),
    .B(net7844));
 sg13g2_o21ai_1 _31556_ (.B1(_08760_),
    .Y(_02335_),
    .A1(net7485),
    .A2(net7844));
 sg13g2_nand2_1 _31557_ (.Y(_08761_),
    .A(net3211),
    .B(net7843));
 sg13g2_o21ai_1 _31558_ (.B1(_08761_),
    .Y(_02336_),
    .A1(net7665),
    .A2(net7843));
 sg13g2_nand2_1 _31559_ (.Y(_08762_),
    .A(net2957),
    .B(net7844));
 sg13g2_o21ai_1 _31560_ (.B1(_08762_),
    .Y(_02337_),
    .A1(net7612),
    .A2(net7844));
 sg13g2_nand2_1 _31561_ (.Y(_08763_),
    .A(net3833),
    .B(net7844));
 sg13g2_o21ai_1 _31562_ (.B1(_08763_),
    .Y(_02338_),
    .A1(net7607),
    .A2(net7845));
 sg13g2_nand2_1 _31563_ (.Y(_08764_),
    .A(net3829),
    .B(net7841));
 sg13g2_o21ai_1 _31564_ (.B1(_08764_),
    .Y(_02339_),
    .A1(net7587),
    .A2(net7841));
 sg13g2_nand2_1 _31565_ (.Y(_08765_),
    .A(net3767),
    .B(net7840));
 sg13g2_o21ai_1 _31566_ (.B1(_08765_),
    .Y(_02340_),
    .A1(net7601),
    .A2(net7840));
 sg13g2_nand2_1 _31567_ (.Y(_08766_),
    .A(net3305),
    .B(net7843));
 sg13g2_o21ai_1 _31568_ (.B1(_08766_),
    .Y(_02341_),
    .A1(net7593),
    .A2(net7843));
 sg13g2_nand2_1 _31569_ (.Y(_08767_),
    .A(net3069),
    .B(net7836));
 sg13g2_o21ai_1 _31570_ (.B1(_08767_),
    .Y(_02342_),
    .A1(net7606),
    .A2(net7836));
 sg13g2_nand2_1 _31571_ (.Y(_08768_),
    .A(net3631),
    .B(net7840));
 sg13g2_o21ai_1 _31572_ (.B1(_08768_),
    .Y(_02343_),
    .A1(net7559),
    .A2(net7840));
 sg13g2_nand2_1 _31573_ (.Y(_08769_),
    .A(net3067),
    .B(net7842));
 sg13g2_o21ai_1 _31574_ (.B1(_08769_),
    .Y(_02344_),
    .A1(net7578),
    .A2(net7842));
 sg13g2_nand2_1 _31575_ (.Y(_08770_),
    .A(net2819),
    .B(net7842));
 sg13g2_o21ai_1 _31576_ (.B1(_08770_),
    .Y(_02345_),
    .A1(net7546),
    .A2(net7842));
 sg13g2_nand2_1 _31577_ (.Y(_08771_),
    .A(net3044),
    .B(net7835));
 sg13g2_o21ai_1 _31578_ (.B1(_08771_),
    .Y(_02346_),
    .A1(net7571),
    .A2(net7835));
 sg13g2_nand2_1 _31579_ (.Y(_08772_),
    .A(net3411),
    .B(net7842));
 sg13g2_o21ai_1 _31580_ (.B1(_08772_),
    .Y(_02347_),
    .A1(net7541),
    .A2(net7842));
 sg13g2_nand2_1 _31581_ (.Y(_08773_),
    .A(net2899),
    .B(net7842));
 sg13g2_o21ai_1 _31582_ (.B1(_08773_),
    .Y(_02348_),
    .A1(net7554),
    .A2(net7842));
 sg13g2_nand2_1 _31583_ (.Y(_08774_),
    .A(net3497),
    .B(net7838));
 sg13g2_o21ai_1 _31584_ (.B1(_08774_),
    .Y(_02349_),
    .A1(net7580),
    .A2(net7838));
 sg13g2_nand2_1 _31585_ (.Y(_08775_),
    .A(net2855),
    .B(net7835));
 sg13g2_o21ai_1 _31586_ (.B1(_08775_),
    .Y(_02350_),
    .A1(net7566),
    .A2(net7835));
 sg13g2_nand2_1 _31587_ (.Y(_08776_),
    .A(net3370),
    .B(net7835));
 sg13g2_o21ai_1 _31588_ (.B1(_08776_),
    .Y(_02351_),
    .A1(net7526),
    .A2(net7835));
 sg13g2_nand2_1 _31589_ (.Y(_08777_),
    .A(net3777),
    .B(net7835));
 sg13g2_o21ai_1 _31590_ (.B1(_08777_),
    .Y(_02352_),
    .A1(net7539),
    .A2(net7835));
 sg13g2_nand2_1 _31591_ (.Y(_08778_),
    .A(net3566),
    .B(net7836));
 sg13g2_o21ai_1 _31592_ (.B1(_08778_),
    .Y(_02353_),
    .A1(net7531),
    .A2(net7836));
 sg13g2_nand2_1 _31593_ (.Y(_08779_),
    .A(net3302),
    .B(net7838));
 sg13g2_o21ai_1 _31594_ (.B1(_08779_),
    .Y(_02354_),
    .A1(net7517),
    .A2(net7838));
 sg13g2_nand2_1 _31595_ (.Y(_08780_),
    .A(net3040),
    .B(net7841));
 sg13g2_o21ai_1 _31596_ (.B1(_08780_),
    .Y(_02355_),
    .A1(net7504),
    .A2(net7841));
 sg13g2_nand2_1 _31597_ (.Y(_08781_),
    .A(net3108),
    .B(_08759_));
 sg13g2_o21ai_1 _31598_ (.B1(_08781_),
    .Y(_02356_),
    .A1(net7512),
    .A2(net7839));
 sg13g2_nand2_1 _31599_ (.Y(_08782_),
    .A(net3770),
    .B(net7845));
 sg13g2_o21ai_1 _31600_ (.B1(_08782_),
    .Y(_02357_),
    .A1(net7494),
    .A2(net7843));
 sg13g2_nand2_1 _31601_ (.Y(_08783_),
    .A(net3754),
    .B(net7837));
 sg13g2_o21ai_1 _31602_ (.B1(_08783_),
    .Y(_02358_),
    .A1(net7503),
    .A2(net7837));
 sg13g2_nand2_1 _31603_ (.Y(_08784_),
    .A(net3125),
    .B(net7840));
 sg13g2_o21ai_1 _31604_ (.B1(_08784_),
    .Y(_02359_),
    .A1(net7646),
    .A2(net7840));
 sg13g2_nand2_1 _31605_ (.Y(_08785_),
    .A(net3779),
    .B(net7844));
 sg13g2_o21ai_1 _31606_ (.B1(_08785_),
    .Y(_02360_),
    .A1(net7649),
    .A2(net7844));
 sg13g2_nand2_1 _31607_ (.Y(_08786_),
    .A(net3789),
    .B(net7843));
 sg13g2_o21ai_1 _31608_ (.B1(_08786_),
    .Y(_02361_),
    .A1(net7656),
    .A2(net7843));
 sg13g2_nand2_1 _31609_ (.Y(_08787_),
    .A(net3894),
    .B(net7839));
 sg13g2_o21ai_1 _31610_ (.B1(_08787_),
    .Y(_02362_),
    .A1(net7661),
    .A2(net7839));
 sg13g2_nand2_1 _31611_ (.Y(_08788_),
    .A(net3360),
    .B(net7839));
 sg13g2_o21ai_1 _31612_ (.B1(_08788_),
    .Y(_02363_),
    .A1(net7640),
    .A2(net7839));
 sg13g2_nand2_1 _31613_ (.Y(_08789_),
    .A(net3653),
    .B(net7840));
 sg13g2_o21ai_1 _31614_ (.B1(_08789_),
    .Y(_02364_),
    .A1(net7628),
    .A2(net7840));
 sg13g2_nand2_1 _31615_ (.Y(_08790_),
    .A(net3116),
    .B(net7839));
 sg13g2_o21ai_1 _31616_ (.B1(_08790_),
    .Y(_02365_),
    .A1(net7619),
    .A2(net7839));
 sg13g2_nand2_1 _31617_ (.Y(_08791_),
    .A(net3409),
    .B(net7836));
 sg13g2_o21ai_1 _31618_ (.B1(_08791_),
    .Y(_02366_),
    .A1(net7630),
    .A2(net7836));
 sg13g2_nand2_1 _31619_ (.Y(_08792_),
    .A(_14301_),
    .B(_03742_));
 sg13g2_nand2_1 _31620_ (.Y(_08793_),
    .A(net3683),
    .B(net7833));
 sg13g2_o21ai_1 _31621_ (.B1(_08793_),
    .Y(_02367_),
    .A1(net7487),
    .A2(net7833));
 sg13g2_nand2_1 _31622_ (.Y(_08794_),
    .A(net3509),
    .B(net7831));
 sg13g2_o21ai_1 _31623_ (.B1(_08794_),
    .Y(_02368_),
    .A1(net7665),
    .A2(net7831));
 sg13g2_nand2_1 _31624_ (.Y(_08795_),
    .A(net3158),
    .B(net7831));
 sg13g2_o21ai_1 _31625_ (.B1(_08795_),
    .Y(_02369_),
    .A1(net7615),
    .A2(net7831));
 sg13g2_nand2_1 _31626_ (.Y(_08796_),
    .A(net2970),
    .B(net7832));
 sg13g2_o21ai_1 _31627_ (.B1(_08796_),
    .Y(_02370_),
    .A1(net7607),
    .A2(net7832));
 sg13g2_nand2_1 _31628_ (.Y(_08797_),
    .A(net2785),
    .B(net7829));
 sg13g2_o21ai_1 _31629_ (.B1(_08797_),
    .Y(_02371_),
    .A1(net7586),
    .A2(net7829));
 sg13g2_nand2_1 _31630_ (.Y(_08798_),
    .A(net2845),
    .B(net7828));
 sg13g2_o21ai_1 _31631_ (.B1(_08798_),
    .Y(_02372_),
    .A1(net7597),
    .A2(net7828));
 sg13g2_nand2_1 _31632_ (.Y(_08799_),
    .A(net2823),
    .B(net7832));
 sg13g2_o21ai_1 _31633_ (.B1(_08799_),
    .Y(_02373_),
    .A1(net7593),
    .A2(net7832));
 sg13g2_nand2_1 _31634_ (.Y(_08800_),
    .A(net2858),
    .B(net7825));
 sg13g2_o21ai_1 _31635_ (.B1(_08800_),
    .Y(_02374_),
    .A1(net7606),
    .A2(net7825));
 sg13g2_nand2_1 _31636_ (.Y(_08801_),
    .A(net2907),
    .B(net7828));
 sg13g2_o21ai_1 _31637_ (.B1(_08801_),
    .Y(_02375_),
    .A1(net7557),
    .A2(net7828));
 sg13g2_nand2_1 _31638_ (.Y(_08802_),
    .A(net2797),
    .B(net7830));
 sg13g2_o21ai_1 _31639_ (.B1(_08802_),
    .Y(_02376_),
    .A1(net7578),
    .A2(net7830));
 sg13g2_nand2_1 _31640_ (.Y(_08803_),
    .A(net3000),
    .B(net7830));
 sg13g2_o21ai_1 _31641_ (.B1(_08803_),
    .Y(_02377_),
    .A1(net7546),
    .A2(net7830));
 sg13g2_nand2_1 _31642_ (.Y(_08804_),
    .A(net3226),
    .B(net7824));
 sg13g2_o21ai_1 _31643_ (.B1(_08804_),
    .Y(_02378_),
    .A1(net7571),
    .A2(net7824));
 sg13g2_nand2_1 _31644_ (.Y(_08805_),
    .A(net2865),
    .B(net7830));
 sg13g2_o21ai_1 _31645_ (.B1(_08805_),
    .Y(_02379_),
    .A1(net7541),
    .A2(net7830));
 sg13g2_nand2_1 _31646_ (.Y(_08806_),
    .A(net3247),
    .B(net7830));
 sg13g2_o21ai_1 _31647_ (.B1(_08806_),
    .Y(_02380_),
    .A1(net7554),
    .A2(net7830));
 sg13g2_nand2_1 _31648_ (.Y(_08807_),
    .A(net2863),
    .B(net7826));
 sg13g2_o21ai_1 _31649_ (.B1(_08807_),
    .Y(_02381_),
    .A1(net7580),
    .A2(net7826));
 sg13g2_nand2_1 _31650_ (.Y(_08808_),
    .A(net2831),
    .B(net7824));
 sg13g2_o21ai_1 _31651_ (.B1(_08808_),
    .Y(_02382_),
    .A1(net7566),
    .A2(net7825));
 sg13g2_nand2_1 _31652_ (.Y(_08809_),
    .A(net2943),
    .B(net7824));
 sg13g2_o21ai_1 _31653_ (.B1(_08809_),
    .Y(_02383_),
    .A1(net7526),
    .A2(net7824));
 sg13g2_nand2_1 _31654_ (.Y(_08810_),
    .A(net2753),
    .B(net7824));
 sg13g2_o21ai_1 _31655_ (.B1(_08810_),
    .Y(_02384_),
    .A1(net7537),
    .A2(net7824));
 sg13g2_nand2_1 _31656_ (.Y(_08811_),
    .A(net2893),
    .B(net7826));
 sg13g2_o21ai_1 _31657_ (.B1(_08811_),
    .Y(_02385_),
    .A1(net7532),
    .A2(net7826));
 sg13g2_nand2_1 _31658_ (.Y(_08812_),
    .A(net2874),
    .B(net7826));
 sg13g2_o21ai_1 _31659_ (.B1(_08812_),
    .Y(_02386_),
    .A1(net7517),
    .A2(net7826));
 sg13g2_nand2_1 _31660_ (.Y(_08813_),
    .A(net2937),
    .B(net7829));
 sg13g2_o21ai_1 _31661_ (.B1(_08813_),
    .Y(_02387_),
    .A1(net7504),
    .A2(net7829));
 sg13g2_nand2_1 _31662_ (.Y(_08814_),
    .A(net2921),
    .B(net7834));
 sg13g2_o21ai_1 _31663_ (.B1(_08814_),
    .Y(_02388_),
    .A1(net7512),
    .A2(net7827));
 sg13g2_nand2_1 _31664_ (.Y(_08815_),
    .A(net3197),
    .B(net7831));
 sg13g2_o21ai_1 _31665_ (.B1(_08815_),
    .Y(_02389_),
    .A1(net7494),
    .A2(net7831));
 sg13g2_nand2_1 _31666_ (.Y(_08816_),
    .A(net3570),
    .B(net7825));
 sg13g2_o21ai_1 _31667_ (.B1(_08816_),
    .Y(_02390_),
    .A1(net7503),
    .A2(net7825));
 sg13g2_nand2_1 _31668_ (.Y(_08817_),
    .A(net3423),
    .B(net7828));
 sg13g2_o21ai_1 _31669_ (.B1(_08817_),
    .Y(_02391_),
    .A1(net7646),
    .A2(net7828));
 sg13g2_nand2_1 _31670_ (.Y(_08818_),
    .A(net2883),
    .B(net7833));
 sg13g2_o21ai_1 _31671_ (.B1(_08818_),
    .Y(_02392_),
    .A1(net7649),
    .A2(net7833));
 sg13g2_nand2_1 _31672_ (.Y(_08819_),
    .A(net3895),
    .B(net7831));
 sg13g2_o21ai_1 _31673_ (.B1(_08819_),
    .Y(_02393_),
    .A1(net7656),
    .A2(net7831));
 sg13g2_nand2_1 _31674_ (.Y(_08820_),
    .A(net3110),
    .B(net7827));
 sg13g2_o21ai_1 _31675_ (.B1(_08820_),
    .Y(_02394_),
    .A1(net7661),
    .A2(net7827));
 sg13g2_nand2_1 _31676_ (.Y(_08821_),
    .A(net2821),
    .B(net7827));
 sg13g2_o21ai_1 _31677_ (.B1(_08821_),
    .Y(_02395_),
    .A1(net7638),
    .A2(net7827));
 sg13g2_nand2_1 _31678_ (.Y(_08822_),
    .A(net3030),
    .B(net7828));
 sg13g2_o21ai_1 _31679_ (.B1(_08822_),
    .Y(_02396_),
    .A1(net7628),
    .A2(net7828));
 sg13g2_nand2_1 _31680_ (.Y(_08823_),
    .A(net3446),
    .B(net7827));
 sg13g2_o21ai_1 _31681_ (.B1(_08823_),
    .Y(_02397_),
    .A1(net7620),
    .A2(net7827));
 sg13g2_nand2_1 _31682_ (.Y(_08824_),
    .A(net3091),
    .B(net7824));
 sg13g2_o21ai_1 _31683_ (.B1(_08824_),
    .Y(_02398_),
    .A1(net7630),
    .A2(net7825));
 sg13g2_nand2_2 _31684_ (.Y(_08825_),
    .A(_14130_),
    .B(_14302_));
 sg13g2_nand2_1 _31685_ (.Y(_08826_),
    .A(net2910),
    .B(net8062));
 sg13g2_o21ai_1 _31686_ (.B1(_08826_),
    .Y(_02399_),
    .A1(net7488),
    .A2(net8062));
 sg13g2_nand2_1 _31687_ (.Y(_08827_),
    .A(net2975),
    .B(net8062));
 sg13g2_o21ai_1 _31688_ (.B1(_08827_),
    .Y(_02400_),
    .A1(net7667),
    .A2(net8062));
 sg13g2_nand2_1 _31689_ (.Y(_08828_),
    .A(net2787),
    .B(net8062));
 sg13g2_o21ai_1 _31690_ (.B1(_08828_),
    .Y(_02401_),
    .A1(net7612),
    .A2(net8062));
 sg13g2_nand2_1 _31691_ (.Y(_08829_),
    .A(net2948),
    .B(net8060));
 sg13g2_o21ai_1 _31692_ (.B1(_08829_),
    .Y(_02402_),
    .A1(net7609),
    .A2(net8060));
 sg13g2_nand2_1 _31693_ (.Y(_08830_),
    .A(net3664),
    .B(net8057));
 sg13g2_o21ai_1 _31694_ (.B1(_08830_),
    .Y(_02403_),
    .A1(net7586),
    .A2(net8057));
 sg13g2_nand2_1 _31695_ (.Y(_08831_),
    .A(net2816),
    .B(net8057));
 sg13g2_o21ai_1 _31696_ (.B1(_08831_),
    .Y(_02404_),
    .A1(net7598),
    .A2(net8057));
 sg13g2_nand2_1 _31697_ (.Y(_08832_),
    .A(net3026),
    .B(net8059));
 sg13g2_o21ai_1 _31698_ (.B1(_08832_),
    .Y(_02405_),
    .A1(net7594),
    .A2(net8059));
 sg13g2_nand2_1 _31699_ (.Y(_08833_),
    .A(net3361),
    .B(net8053));
 sg13g2_o21ai_1 _31700_ (.B1(_08833_),
    .Y(_02406_),
    .A1(net7602),
    .A2(net8053));
 sg13g2_nand2_1 _31701_ (.Y(_08834_),
    .A(net2961),
    .B(net8058));
 sg13g2_o21ai_1 _31702_ (.B1(_08834_),
    .Y(_02407_),
    .A1(net7559),
    .A2(net8058));
 sg13g2_nand2_1 _31703_ (.Y(_08835_),
    .A(net3074),
    .B(net8061));
 sg13g2_o21ai_1 _31704_ (.B1(_08835_),
    .Y(_02408_),
    .A1(net7576),
    .A2(net8061));
 sg13g2_nand2_1 _31705_ (.Y(_08836_),
    .A(net2864),
    .B(net8059));
 sg13g2_o21ai_1 _31706_ (.B1(_08836_),
    .Y(_02409_),
    .A1(net7548),
    .A2(net8059));
 sg13g2_nand2_1 _31707_ (.Y(_08837_),
    .A(net3250),
    .B(net8053));
 sg13g2_o21ai_1 _31708_ (.B1(_08837_),
    .Y(_02410_),
    .A1(net7568),
    .A2(net8053));
 sg13g2_nand2_1 _31709_ (.Y(_08838_),
    .A(net3807),
    .B(net8059));
 sg13g2_o21ai_1 _31710_ (.B1(_08838_),
    .Y(_02411_),
    .A1(net7544),
    .A2(net8059));
 sg13g2_nand2_1 _31711_ (.Y(_08839_),
    .A(net3177),
    .B(net8061));
 sg13g2_o21ai_1 _31712_ (.B1(_08839_),
    .Y(_02412_),
    .A1(net7552),
    .A2(net8061));
 sg13g2_nand2_1 _31713_ (.Y(_08840_),
    .A(net4267),
    .B(net8056));
 sg13g2_o21ai_1 _31714_ (.B1(_08840_),
    .Y(_02413_),
    .A1(_12964_),
    .A2(net8056));
 sg13g2_nand2_1 _31715_ (.Y(_08841_),
    .A(net2966),
    .B(net8054));
 sg13g2_o21ai_1 _31716_ (.B1(_08841_),
    .Y(_02414_),
    .A1(net7564),
    .A2(net8054));
 sg13g2_nand2_1 _31717_ (.Y(_08842_),
    .A(net2927),
    .B(net8053));
 sg13g2_o21ai_1 _31718_ (.B1(_08842_),
    .Y(_02415_),
    .A1(net7522),
    .A2(net8053));
 sg13g2_nand2_1 _31719_ (.Y(_08843_),
    .A(net3209),
    .B(net8053));
 sg13g2_o21ai_1 _31720_ (.B1(_08843_),
    .Y(_02416_),
    .A1(net7534),
    .A2(net8053));
 sg13g2_nand2_1 _31721_ (.Y(_08844_),
    .A(net2806),
    .B(net8054));
 sg13g2_o21ai_1 _31722_ (.B1(_08844_),
    .Y(_02417_),
    .A1(net7528),
    .A2(net8054));
 sg13g2_nand2_1 _31723_ (.Y(_08845_),
    .A(net2891),
    .B(net8055));
 sg13g2_o21ai_1 _31724_ (.B1(_08845_),
    .Y(_02418_),
    .A1(net7518),
    .A2(net8055));
 sg13g2_nand2_1 _31725_ (.Y(_08846_),
    .A(net3278),
    .B(net8058));
 sg13g2_o21ai_1 _31726_ (.B1(_08846_),
    .Y(_02419_),
    .A1(net7505),
    .A2(net8058));
 sg13g2_nand2_1 _31727_ (.Y(_08847_),
    .A(net3537),
    .B(net8057));
 sg13g2_o21ai_1 _31728_ (.B1(_08847_),
    .Y(_02420_),
    .A1(net7513),
    .A2(net8057));
 sg13g2_nand2_1 _31729_ (.Y(_08848_),
    .A(net3702),
    .B(net8060));
 sg13g2_o21ai_1 _31730_ (.B1(_08848_),
    .Y(_02421_),
    .A1(net7496),
    .A2(net8060));
 sg13g2_nand2_1 _31731_ (.Y(_08849_),
    .A(net2880),
    .B(net8054));
 sg13g2_o21ai_1 _31732_ (.B1(_08849_),
    .Y(_02422_),
    .A1(net7502),
    .A2(net8054));
 sg13g2_nand2_1 _31733_ (.Y(_08850_),
    .A(net3536),
    .B(net8057));
 sg13g2_o21ai_1 _31734_ (.B1(_08850_),
    .Y(_02423_),
    .A1(net7643),
    .A2(net8057));
 sg13g2_nand2_1 _31735_ (.Y(_08851_),
    .A(net2834),
    .B(net8062));
 sg13g2_o21ai_1 _31736_ (.B1(_08851_),
    .Y(_02424_),
    .A1(net7650),
    .A2(net8062));
 sg13g2_nand2_1 _31737_ (.Y(_08852_),
    .A(net3389),
    .B(net8059));
 sg13g2_o21ai_1 _31738_ (.B1(_08852_),
    .Y(_02425_),
    .A1(net7655),
    .A2(net8059));
 sg13g2_nand2_1 _31739_ (.Y(_08853_),
    .A(net3511),
    .B(net8055));
 sg13g2_o21ai_1 _31740_ (.B1(_08853_),
    .Y(_02426_),
    .A1(net7659),
    .A2(net8055));
 sg13g2_nand2_1 _31741_ (.Y(_08854_),
    .A(net2960),
    .B(net8055));
 sg13g2_o21ai_1 _31742_ (.B1(_08854_),
    .Y(_02427_),
    .A1(net7638),
    .A2(net8055));
 sg13g2_nand2_1 _31743_ (.Y(_08855_),
    .A(net2932),
    .B(net8058));
 sg13g2_o21ai_1 _31744_ (.B1(_08855_),
    .Y(_02428_),
    .A1(net7625),
    .A2(net8058));
 sg13g2_nand2_1 _31745_ (.Y(_08856_),
    .A(net3267),
    .B(net8055));
 sg13g2_o21ai_1 _31746_ (.B1(_08856_),
    .Y(_02429_),
    .A1(net7622),
    .A2(net8055));
 sg13g2_nand2_1 _31747_ (.Y(_08857_),
    .A(net2852),
    .B(net8056));
 sg13g2_o21ai_1 _31748_ (.B1(_08857_),
    .Y(_02430_),
    .A1(net7631),
    .A2(net8056));
 sg13g2_nand3_1 _31749_ (.B(net8371),
    .C(_14130_),
    .A(net8961),
    .Y(_08858_));
 sg13g2_nand2_1 _31750_ (.Y(_08859_),
    .A(net2645),
    .B(net8051));
 sg13g2_o21ai_1 _31751_ (.B1(_08859_),
    .Y(_02431_),
    .A1(net7488),
    .A2(net8051));
 sg13g2_nand2_1 _31752_ (.Y(_08860_),
    .A(net4042),
    .B(net8051));
 sg13g2_o21ai_1 _31753_ (.B1(_08860_),
    .Y(_02432_),
    .A1(net7667),
    .A2(net8051));
 sg13g2_nand2_1 _31754_ (.Y(_08861_),
    .A(net3613),
    .B(net8051));
 sg13g2_o21ai_1 _31755_ (.B1(_08861_),
    .Y(_02433_),
    .A1(net7613),
    .A2(net8051));
 sg13g2_nand2_1 _31756_ (.Y(_08862_),
    .A(net3595),
    .B(net8049));
 sg13g2_o21ai_1 _31757_ (.B1(_08862_),
    .Y(_02434_),
    .A1(net7609),
    .A2(net8049));
 sg13g2_nand2_1 _31758_ (.Y(_08863_),
    .A(net3744),
    .B(net8046));
 sg13g2_o21ai_1 _31759_ (.B1(_08863_),
    .Y(_02435_),
    .A1(net7588),
    .A2(net8046));
 sg13g2_nand2_1 _31760_ (.Y(_08864_),
    .A(net3535),
    .B(net8046));
 sg13g2_o21ai_1 _31761_ (.B1(_08864_),
    .Y(_02436_),
    .A1(net7598),
    .A2(net8046));
 sg13g2_nand2_1 _31762_ (.Y(_08865_),
    .A(net3301),
    .B(net8048));
 sg13g2_o21ai_1 _31763_ (.B1(_08865_),
    .Y(_02437_),
    .A1(net7594),
    .A2(net8048));
 sg13g2_nand2_1 _31764_ (.Y(_08866_),
    .A(net3675),
    .B(net8042));
 sg13g2_o21ai_1 _31765_ (.B1(_08866_),
    .Y(_02438_),
    .A1(net7602),
    .A2(net8042));
 sg13g2_nand2_1 _31766_ (.Y(_08867_),
    .A(net3263),
    .B(net8047));
 sg13g2_o21ai_1 _31767_ (.B1(_08867_),
    .Y(_02439_),
    .A1(net7557),
    .A2(net8047));
 sg13g2_nand2_1 _31768_ (.Y(_08868_),
    .A(net3172),
    .B(net8050));
 sg13g2_o21ai_1 _31769_ (.B1(_08868_),
    .Y(_02440_),
    .A1(net7574),
    .A2(net8050));
 sg13g2_nand2_1 _31770_ (.Y(_08869_),
    .A(net3033),
    .B(net8048));
 sg13g2_o21ai_1 _31771_ (.B1(_08869_),
    .Y(_02441_),
    .A1(net7550),
    .A2(net8048));
 sg13g2_nand2_1 _31772_ (.Y(_08870_),
    .A(net4013),
    .B(net8042));
 sg13g2_o21ai_1 _31773_ (.B1(_08870_),
    .Y(_02442_),
    .A1(net7568),
    .A2(net8042));
 sg13g2_nand2_1 _31774_ (.Y(_08871_),
    .A(net3608),
    .B(net8048));
 sg13g2_o21ai_1 _31775_ (.B1(_08871_),
    .Y(_02443_),
    .A1(net7544),
    .A2(net8048));
 sg13g2_nand2_1 _31776_ (.Y(_08872_),
    .A(net3159),
    .B(net8050));
 sg13g2_o21ai_1 _31777_ (.B1(_08872_),
    .Y(_02444_),
    .A1(net7552),
    .A2(net8050));
 sg13g2_nand2_1 _31778_ (.Y(_08873_),
    .A(net3192),
    .B(net8045));
 sg13g2_o21ai_1 _31779_ (.B1(_08873_),
    .Y(_02445_),
    .A1(net7585),
    .A2(net8045));
 sg13g2_nand2_1 _31780_ (.Y(_08874_),
    .A(net3898),
    .B(net8043));
 sg13g2_o21ai_1 _31781_ (.B1(_08874_),
    .Y(_02446_),
    .A1(net7565),
    .A2(net8043));
 sg13g2_nand2_1 _31782_ (.Y(_08875_),
    .A(net3520),
    .B(net8042));
 sg13g2_o21ai_1 _31783_ (.B1(_08875_),
    .Y(_02447_),
    .A1(net7522),
    .A2(net8042));
 sg13g2_nand2_1 _31784_ (.Y(_08876_),
    .A(net3636),
    .B(net8043));
 sg13g2_o21ai_1 _31785_ (.B1(_08876_),
    .Y(_02448_),
    .A1(net7535),
    .A2(net8043));
 sg13g2_nand2_1 _31786_ (.Y(_08877_),
    .A(net3578),
    .B(net8042));
 sg13g2_o21ai_1 _31787_ (.B1(_08877_),
    .Y(_02449_),
    .A1(net7528),
    .A2(net8042));
 sg13g2_nand2_1 _31788_ (.Y(_08878_),
    .A(net3788),
    .B(net8044));
 sg13g2_o21ai_1 _31789_ (.B1(_08878_),
    .Y(_02450_),
    .A1(net7516),
    .A2(net8044));
 sg13g2_nand2_1 _31790_ (.Y(_08879_),
    .A(net2904),
    .B(net8047));
 sg13g2_o21ai_1 _31791_ (.B1(_08879_),
    .Y(_02451_),
    .A1(net7505),
    .A2(net8047));
 sg13g2_nand2_1 _31792_ (.Y(_08880_),
    .A(net2987),
    .B(net8046));
 sg13g2_o21ai_1 _31793_ (.B1(_08880_),
    .Y(_02452_),
    .A1(net7512),
    .A2(net8046));
 sg13g2_nand2_1 _31794_ (.Y(_08881_),
    .A(net3697),
    .B(net8049));
 sg13g2_o21ai_1 _31795_ (.B1(_08881_),
    .Y(_02453_),
    .A1(net7496),
    .A2(net8049));
 sg13g2_nand2_1 _31796_ (.Y(_08882_),
    .A(net3709),
    .B(net8043));
 sg13g2_o21ai_1 _31797_ (.B1(_08882_),
    .Y(_02454_),
    .A1(net7500),
    .A2(net8043));
 sg13g2_nand2_1 _31798_ (.Y(_08883_),
    .A(net4157),
    .B(net8046));
 sg13g2_o21ai_1 _31799_ (.B1(_08883_),
    .Y(_02455_),
    .A1(net7643),
    .A2(net8046));
 sg13g2_nand2_1 _31800_ (.Y(_08884_),
    .A(net3483),
    .B(net8051));
 sg13g2_o21ai_1 _31801_ (.B1(_08884_),
    .Y(_02456_),
    .A1(net7650),
    .A2(net8051));
 sg13g2_nand2_1 _31802_ (.Y(_08885_),
    .A(net3525),
    .B(net8048));
 sg13g2_o21ai_1 _31803_ (.B1(_08885_),
    .Y(_02457_),
    .A1(net7655),
    .A2(net8048));
 sg13g2_nand2_1 _31804_ (.Y(_08886_),
    .A(net3505),
    .B(net8044));
 sg13g2_o21ai_1 _31805_ (.B1(_08886_),
    .Y(_02458_),
    .A1(net7659),
    .A2(net8044));
 sg13g2_nand2_1 _31806_ (.Y(_08887_),
    .A(net3580),
    .B(net8044));
 sg13g2_o21ai_1 _31807_ (.B1(_08887_),
    .Y(_02459_),
    .A1(net7638),
    .A2(net8044));
 sg13g2_nand2_1 _31808_ (.Y(_08888_),
    .A(net3474),
    .B(net8047));
 sg13g2_o21ai_1 _31809_ (.B1(_08888_),
    .Y(_02460_),
    .A1(net7625),
    .A2(net8047));
 sg13g2_nand2_1 _31810_ (.Y(_08889_),
    .A(net3173),
    .B(net8044));
 sg13g2_o21ai_1 _31811_ (.B1(_08889_),
    .Y(_02461_),
    .A1(net7621),
    .A2(net8044));
 sg13g2_nand2_1 _31812_ (.Y(_08890_),
    .A(net3077),
    .B(net8045));
 sg13g2_o21ai_1 _31813_ (.B1(_08890_),
    .Y(_02462_),
    .A1(net7630),
    .A2(net8045));
 sg13g2_nand3_1 _31814_ (.B(net8372),
    .C(_14199_),
    .A(_12607_),
    .Y(_08891_));
 sg13g2_nand2_1 _31815_ (.Y(_08892_),
    .A(net3324),
    .B(net8040));
 sg13g2_o21ai_1 _31816_ (.B1(_08892_),
    .Y(_02463_),
    .A1(net7486),
    .A2(net8040));
 sg13g2_nand2_1 _31817_ (.Y(_08893_),
    .A(net3222),
    .B(net8040));
 sg13g2_o21ai_1 _31818_ (.B1(_08893_),
    .Y(_02464_),
    .A1(net7663),
    .A2(net8040));
 sg13g2_nand2_1 _31819_ (.Y(_08894_),
    .A(net3335),
    .B(net8040));
 sg13g2_o21ai_1 _31820_ (.B1(_08894_),
    .Y(_02465_),
    .A1(net7612),
    .A2(net8040));
 sg13g2_nand2_1 _31821_ (.Y(_08895_),
    .A(net4025),
    .B(net8038));
 sg13g2_o21ai_1 _31822_ (.B1(_08895_),
    .Y(_02466_),
    .A1(net7609),
    .A2(net8038));
 sg13g2_nand2_1 _31823_ (.Y(_08896_),
    .A(net3682),
    .B(net8036));
 sg13g2_o21ai_1 _31824_ (.B1(_08896_),
    .Y(_02467_),
    .A1(net7588),
    .A2(net8036));
 sg13g2_nand2_1 _31825_ (.Y(_08897_),
    .A(net3412),
    .B(net8035));
 sg13g2_o21ai_1 _31826_ (.B1(_08897_),
    .Y(_02468_),
    .A1(net7600),
    .A2(net8035));
 sg13g2_nand2_1 _31827_ (.Y(_08898_),
    .A(net3291),
    .B(net8037));
 sg13g2_o21ai_1 _31828_ (.B1(_08898_),
    .Y(_02469_),
    .A1(net7594),
    .A2(net8037));
 sg13g2_nand2_1 _31829_ (.Y(_08899_),
    .A(net3552),
    .B(net8030));
 sg13g2_o21ai_1 _31830_ (.B1(_08899_),
    .Y(_02470_),
    .A1(net7602),
    .A2(net8030));
 sg13g2_nand2_1 _31831_ (.Y(_08900_),
    .A(net4174),
    .B(net8036));
 sg13g2_o21ai_1 _31832_ (.B1(_08900_),
    .Y(_02471_),
    .A1(net7562),
    .A2(net8036));
 sg13g2_nand2_1 _31833_ (.Y(_08901_),
    .A(net3983),
    .B(net8039));
 sg13g2_o21ai_1 _31834_ (.B1(_08901_),
    .Y(_02472_),
    .A1(net7577),
    .A2(net8039));
 sg13g2_nand2_1 _31835_ (.Y(_08902_),
    .A(net3479),
    .B(net8037));
 sg13g2_o21ai_1 _31836_ (.B1(_08902_),
    .Y(_02473_),
    .A1(net7548),
    .A2(net8037));
 sg13g2_nand2_1 _31837_ (.Y(_08903_),
    .A(net3512),
    .B(net8030));
 sg13g2_o21ai_1 _31838_ (.B1(_08903_),
    .Y(_02474_),
    .A1(net7568),
    .A2(net8030));
 sg13g2_nand2_1 _31839_ (.Y(_08904_),
    .A(net3973),
    .B(net8037));
 sg13g2_o21ai_1 _31840_ (.B1(_08904_),
    .Y(_02475_),
    .A1(net7543),
    .A2(net8037));
 sg13g2_nand2_1 _31841_ (.Y(_08905_),
    .A(net2946),
    .B(net8039));
 sg13g2_o21ai_1 _31842_ (.B1(_08905_),
    .Y(_02476_),
    .A1(net7552),
    .A2(net8039));
 sg13g2_nand2_1 _31843_ (.Y(_08906_),
    .A(net3332),
    .B(net8034));
 sg13g2_o21ai_1 _31844_ (.B1(_08906_),
    .Y(_02477_),
    .A1(net7585),
    .A2(net8034));
 sg13g2_nand2_1 _31845_ (.Y(_08907_),
    .A(net3635),
    .B(net8031));
 sg13g2_o21ai_1 _31846_ (.B1(_08907_),
    .Y(_02478_),
    .A1(net7563),
    .A2(net8031));
 sg13g2_nand2_1 _31847_ (.Y(_08908_),
    .A(net3764),
    .B(net8030));
 sg13g2_o21ai_1 _31848_ (.B1(_08908_),
    .Y(_02479_),
    .A1(net7522),
    .A2(net8030));
 sg13g2_nand2_1 _31849_ (.Y(_08909_),
    .A(net3290),
    .B(net8030));
 sg13g2_o21ai_1 _31850_ (.B1(_08909_),
    .Y(_02480_),
    .A1(net7534),
    .A2(net8030));
 sg13g2_nand2_1 _31851_ (.Y(_08910_),
    .A(net3659),
    .B(net8031));
 sg13g2_o21ai_1 _31852_ (.B1(_08910_),
    .Y(_02481_),
    .A1(net7529),
    .A2(net8031));
 sg13g2_nand2_1 _31853_ (.Y(_08911_),
    .A(net3422),
    .B(net8033));
 sg13g2_o21ai_1 _31854_ (.B1(_08911_),
    .Y(_02482_),
    .A1(net7518),
    .A2(net8033));
 sg13g2_nand2_1 _31855_ (.Y(_08912_),
    .A(net3842),
    .B(net8036));
 sg13g2_o21ai_1 _31856_ (.B1(_08912_),
    .Y(_02483_),
    .A1(net7509),
    .A2(net8036));
 sg13g2_nand2_1 _31857_ (.Y(_08913_),
    .A(net3681),
    .B(net8035));
 sg13g2_o21ai_1 _31858_ (.B1(_08913_),
    .Y(_02484_),
    .A1(net7514),
    .A2(net8035));
 sg13g2_nand2_1 _31859_ (.Y(_08914_),
    .A(net3901),
    .B(net8038));
 sg13g2_o21ai_1 _31860_ (.B1(_08914_),
    .Y(_02485_),
    .A1(net7496),
    .A2(net8038));
 sg13g2_nand2_1 _31861_ (.Y(_08915_),
    .A(net3734),
    .B(net8031));
 sg13g2_o21ai_1 _31862_ (.B1(_08915_),
    .Y(_02486_),
    .A1(net7500),
    .A2(net8031));
 sg13g2_nand2_1 _31863_ (.Y(_08916_),
    .A(net3079),
    .B(net8035));
 sg13g2_o21ai_1 _31864_ (.B1(_08916_),
    .Y(_02487_),
    .A1(net7643),
    .A2(net8035));
 sg13g2_nand2_1 _31865_ (.Y(_08917_),
    .A(net3123),
    .B(net8040));
 sg13g2_o21ai_1 _31866_ (.B1(_08917_),
    .Y(_02488_),
    .A1(net7650),
    .A2(net8040));
 sg13g2_nand2_1 _31867_ (.Y(_08918_),
    .A(net3217),
    .B(net8037));
 sg13g2_o21ai_1 _31868_ (.B1(_08918_),
    .Y(_02489_),
    .A1(net7655),
    .A2(net8037));
 sg13g2_nand2_1 _31869_ (.Y(_08919_),
    .A(net3816),
    .B(net8033));
 sg13g2_o21ai_1 _31870_ (.B1(_08919_),
    .Y(_02490_),
    .A1(net7659),
    .A2(net8033));
 sg13g2_nand2_1 _31871_ (.Y(_08920_),
    .A(net3382),
    .B(net8033));
 sg13g2_o21ai_1 _31872_ (.B1(_08920_),
    .Y(_02491_),
    .A1(net7638),
    .A2(net8033));
 sg13g2_nand2_1 _31873_ (.Y(_08921_),
    .A(net3879),
    .B(net8035));
 sg13g2_o21ai_1 _31874_ (.B1(_08921_),
    .Y(_02492_),
    .A1(net7628),
    .A2(net8035));
 sg13g2_nand2_1 _31875_ (.Y(_08922_),
    .A(net3888),
    .B(net8033));
 sg13g2_o21ai_1 _31876_ (.B1(_08922_),
    .Y(_02493_),
    .A1(net7622),
    .A2(net8033));
 sg13g2_nand2_1 _31877_ (.Y(_08923_),
    .A(net3487),
    .B(net8032));
 sg13g2_o21ai_1 _31878_ (.B1(_08923_),
    .Y(_02494_),
    .A1(net7633),
    .A2(net8032));
 sg13g2_and3_1 _31879_ (.X(_08924_),
    .A(net9710),
    .B(net8371),
    .C(_02848_));
 sg13g2_nand2_2 _31880_ (.Y(_08925_),
    .A(_14199_),
    .B(_08924_));
 sg13g2_nand2_1 _31881_ (.Y(_08926_),
    .A(net3565),
    .B(net7968));
 sg13g2_o21ai_1 _31882_ (.B1(_08926_),
    .Y(_02495_),
    .A1(net7485),
    .A2(net7968));
 sg13g2_nand2_1 _31883_ (.Y(_08927_),
    .A(net3328),
    .B(net7967));
 sg13g2_o21ai_1 _31884_ (.B1(_08927_),
    .Y(_02496_),
    .A1(net7664),
    .A2(net7967));
 sg13g2_nand2_1 _31885_ (.Y(_08928_),
    .A(net3749),
    .B(net7965));
 sg13g2_o21ai_1 _31886_ (.B1(_08928_),
    .Y(_02497_),
    .A1(net7614),
    .A2(net7965));
 sg13g2_nand2_1 _31887_ (.Y(_08929_),
    .A(net3277),
    .B(net7966));
 sg13g2_o21ai_1 _31888_ (.B1(_08929_),
    .Y(_02498_),
    .A1(net7608),
    .A2(net7966));
 sg13g2_nand2_1 _31889_ (.Y(_08930_),
    .A(net3562),
    .B(net7963));
 sg13g2_o21ai_1 _31890_ (.B1(_08930_),
    .Y(_02499_),
    .A1(net7588),
    .A2(net7963));
 sg13g2_nand2_1 _31891_ (.Y(_08931_),
    .A(net3844),
    .B(net7963));
 sg13g2_o21ai_1 _31892_ (.B1(_08931_),
    .Y(_02500_),
    .A1(net7599),
    .A2(net7963));
 sg13g2_nand2_1 _31893_ (.Y(_08932_),
    .A(net2990),
    .B(net7966));
 sg13g2_o21ai_1 _31894_ (.B1(_08932_),
    .Y(_02501_),
    .A1(net7592),
    .A2(net7966));
 sg13g2_nand2_1 _31895_ (.Y(_08933_),
    .A(net2722),
    .B(net7961));
 sg13g2_o21ai_1 _31896_ (.B1(_08933_),
    .Y(_02502_),
    .A1(net7605),
    .A2(net7961));
 sg13g2_nand2_1 _31897_ (.Y(_08934_),
    .A(net2639),
    .B(net7964));
 sg13g2_o21ai_1 _31898_ (.B1(_08934_),
    .Y(_02503_),
    .A1(net7561),
    .A2(net7964));
 sg13g2_nand2_1 _31899_ (.Y(_08935_),
    .A(net3349),
    .B(net7965));
 sg13g2_o21ai_1 _31900_ (.B1(_08935_),
    .Y(_02504_),
    .A1(net7578),
    .A2(net7965));
 sg13g2_nand2_1 _31901_ (.Y(_08936_),
    .A(net3998),
    .B(net7967));
 sg13g2_o21ai_1 _31902_ (.B1(_08936_),
    .Y(_02505_),
    .A1(net7546),
    .A2(net7967));
 sg13g2_nand2_1 _31903_ (.Y(_08937_),
    .A(net3880),
    .B(net7959));
 sg13g2_o21ai_1 _31904_ (.B1(_08937_),
    .Y(_02506_),
    .A1(net7571),
    .A2(net7959));
 sg13g2_nand2_1 _31905_ (.Y(_08938_),
    .A(net3718),
    .B(net7965));
 sg13g2_o21ai_1 _31906_ (.B1(_08938_),
    .Y(_02507_),
    .A1(net7540),
    .A2(net7965));
 sg13g2_nand2_1 _31907_ (.Y(_08939_),
    .A(net3544),
    .B(net7965));
 sg13g2_o21ai_1 _31908_ (.B1(_08939_),
    .Y(_02508_),
    .A1(net7554),
    .A2(net7965));
 sg13g2_nand2_1 _31909_ (.Y(_08940_),
    .A(net2644),
    .B(net7962));
 sg13g2_o21ai_1 _31910_ (.B1(_08940_),
    .Y(_02509_),
    .A1(net7583),
    .A2(net7962));
 sg13g2_nand2_1 _31911_ (.Y(_08941_),
    .A(net3424),
    .B(net7960));
 sg13g2_o21ai_1 _31912_ (.B1(_08941_),
    .Y(_02510_),
    .A1(net7565),
    .A2(net7960));
 sg13g2_nand2_1 _31913_ (.Y(_08942_),
    .A(net3087),
    .B(net7959));
 sg13g2_o21ai_1 _31914_ (.B1(_08942_),
    .Y(_02511_),
    .A1(net7525),
    .A2(net7959));
 sg13g2_nand2_1 _31915_ (.Y(_08943_),
    .A(net3089),
    .B(net7959));
 sg13g2_o21ai_1 _31916_ (.B1(_08943_),
    .Y(_02512_),
    .A1(net7537),
    .A2(net7959));
 sg13g2_nand2_1 _31917_ (.Y(_08944_),
    .A(net3736),
    .B(net7960));
 sg13g2_o21ai_1 _31918_ (.B1(_08944_),
    .Y(_02513_),
    .A1(net7532),
    .A2(net7960));
 sg13g2_nand2_1 _31919_ (.Y(_08945_),
    .A(net4352),
    .B(net7960));
 sg13g2_o21ai_1 _31920_ (.B1(_08945_),
    .Y(_02514_),
    .A1(net7516),
    .A2(net7960));
 sg13g2_nand2_1 _31921_ (.Y(_08946_),
    .A(net3007),
    .B(net7968));
 sg13g2_o21ai_1 _31922_ (.B1(_08946_),
    .Y(_02515_),
    .A1(net7506),
    .A2(net7968));
 sg13g2_nand2_1 _31923_ (.Y(_08947_),
    .A(net3906),
    .B(net7963));
 sg13g2_o21ai_1 _31924_ (.B1(_08947_),
    .Y(_02516_),
    .A1(net7513),
    .A2(net7963));
 sg13g2_nand2_1 _31925_ (.Y(_08948_),
    .A(net3655),
    .B(net7966));
 sg13g2_o21ai_1 _31926_ (.B1(_08948_),
    .Y(_02517_),
    .A1(net7497),
    .A2(net7966));
 sg13g2_nand2_1 _31927_ (.Y(_08949_),
    .A(net3189),
    .B(net7959));
 sg13g2_o21ai_1 _31928_ (.B1(_08949_),
    .Y(_02518_),
    .A1(net7501),
    .A2(net7959));
 sg13g2_nand2_1 _31929_ (.Y(_08950_),
    .A(net3582),
    .B(net7963));
 sg13g2_o21ai_1 _31930_ (.B1(_08950_),
    .Y(_02519_),
    .A1(net7642),
    .A2(net7963));
 sg13g2_nand2_1 _31931_ (.Y(_08951_),
    .A(net3915),
    .B(net7968));
 sg13g2_o21ai_1 _31932_ (.B1(_08951_),
    .Y(_02520_),
    .A1(net7652),
    .A2(net7968));
 sg13g2_nand2_1 _31933_ (.Y(_08952_),
    .A(net3647),
    .B(net7966));
 sg13g2_o21ai_1 _31934_ (.B1(_08952_),
    .Y(_02521_),
    .A1(net7653),
    .A2(net7966));
 sg13g2_nand2_1 _31935_ (.Y(_08953_),
    .A(net3853),
    .B(net7961));
 sg13g2_o21ai_1 _31936_ (.B1(_08953_),
    .Y(_02522_),
    .A1(net7659),
    .A2(net7961));
 sg13g2_nand2_1 _31937_ (.Y(_08954_),
    .A(net3685),
    .B(net7962));
 sg13g2_o21ai_1 _31938_ (.B1(_08954_),
    .Y(_02523_),
    .A1(net7637),
    .A2(net7961));
 sg13g2_nand2_1 _31939_ (.Y(_08955_),
    .A(net3696),
    .B(net7964));
 sg13g2_o21ai_1 _31940_ (.B1(_08955_),
    .Y(_02524_),
    .A1(net7627),
    .A2(net7964));
 sg13g2_nand2_1 _31941_ (.Y(_08956_),
    .A(net3663),
    .B(net7962));
 sg13g2_o21ai_1 _31942_ (.B1(_08956_),
    .Y(_02525_),
    .A1(net7619),
    .A2(net7961));
 sg13g2_nand2_1 _31943_ (.Y(_08957_),
    .A(net2903),
    .B(net7961));
 sg13g2_o21ai_1 _31944_ (.B1(_08957_),
    .Y(_02526_),
    .A1(net7634),
    .A2(net7960));
 sg13g2_nand2b_1 _31945_ (.Y(_08958_),
    .B(net8938),
    .A_N(_06967_));
 sg13g2_o21ai_1 _31946_ (.B1(_07036_),
    .Y(_08959_),
    .A1(net3927),
    .A2(net8935));
 sg13g2_a21oi_1 _31947_ (.A1(_08958_),
    .A2(_08959_),
    .Y(_02527_),
    .B1(net9006));
 sg13g2_o21ai_1 _31948_ (.B1(_07036_),
    .Y(_08960_),
    .A1(net5289),
    .A2(net8935));
 sg13g2_a21oi_1 _31949_ (.A1(_08958_),
    .A2(_08960_),
    .Y(_02528_),
    .B1(net9006));
 sg13g2_nand2b_1 _31950_ (.Y(_08961_),
    .B(_07301_),
    .A_N(_07208_));
 sg13g2_a21oi_1 _31951_ (.A1(net8683),
    .A2(_07185_),
    .Y(_08962_),
    .B1(_08961_));
 sg13g2_inv_1 _31952_ (.Y(_08963_),
    .A(net8319));
 sg13g2_o21ai_1 _31953_ (.B1(net8603),
    .Y(_08964_),
    .A1(_13971_),
    .A2(_14297_));
 sg13g2_nor2b_1 _31954_ (.A(net9255),
    .B_N(\soc_I.qqspi_I.spi_buf[7] ),
    .Y(_08965_));
 sg13g2_a21oi_1 _31955_ (.A1(\soc_I.qqspi_I.spi_buf[4] ),
    .A2(net9258),
    .Y(_08966_),
    .B1(_08965_));
 sg13g2_a221oi_1 _31956_ (.B2(net8680),
    .C1(_08963_),
    .B1(_08966_),
    .A1(_13979_),
    .Y(_08967_),
    .A2(net8582));
 sg13g2_a22oi_1 _31957_ (.Y(_08968_),
    .B1(_08964_),
    .B2(_08967_),
    .A2(_08963_),
    .A1(net5191));
 sg13g2_nor2_1 _31958_ (.A(net9021),
    .B(_08968_),
    .Y(_02529_));
 sg13g2_nor2b_1 _31959_ (.A(net9264),
    .B_N(\soc_I.qqspi_I.spi_buf[8] ),
    .Y(_08969_));
 sg13g2_a21oi_1 _31960_ (.A1(net5198),
    .A2(net9259),
    .Y(_08970_),
    .B1(_08969_));
 sg13g2_a22oi_1 _31961_ (.Y(_08971_),
    .B1(_08970_),
    .B2(net8680),
    .A2(net8582),
    .A1(_13988_));
 sg13g2_o21ai_1 _31962_ (.B1(_08971_),
    .Y(_08972_),
    .A1(_14274_),
    .A2(_07323_));
 sg13g2_o21ai_1 _31963_ (.B1(net9344),
    .Y(_08973_),
    .A1(net5435),
    .A2(net8319));
 sg13g2_a21oi_1 _31964_ (.A1(net8319),
    .A2(_08972_),
    .Y(_02530_),
    .B1(_08973_));
 sg13g2_nand2b_1 _31965_ (.Y(_08974_),
    .B(net9255),
    .A_N(\soc_I.qqspi_I.spi_buf[6] ));
 sg13g2_o21ai_1 _31966_ (.B1(_08974_),
    .Y(_08975_),
    .A1(\soc_I.qqspi_I.spi_buf[9] ),
    .A2(net9255));
 sg13g2_o21ai_1 _31967_ (.B1(net8322),
    .Y(_08976_),
    .A1(net8686),
    .A2(_08975_));
 sg13g2_a221oi_1 _31968_ (.B2(_13994_),
    .C1(_08976_),
    .B1(net8582),
    .A1(net7493),
    .Y(_08977_),
    .A2(net8603));
 sg13g2_o21ai_1 _31969_ (.B1(net9342),
    .Y(_08978_),
    .A1(net5365),
    .A2(net8322));
 sg13g2_nor2_1 _31970_ (.A(_08977_),
    .B(_08978_),
    .Y(_02531_));
 sg13g2_nand2b_1 _31971_ (.Y(_08979_),
    .B(net9255),
    .A_N(\soc_I.qqspi_I.spi_buf[7] ));
 sg13g2_o21ai_1 _31972_ (.B1(_08979_),
    .Y(_08980_),
    .A1(\soc_I.qqspi_I.spi_buf[10] ),
    .A2(net9257));
 sg13g2_o21ai_1 _31973_ (.B1(net8319),
    .Y(_08981_),
    .A1(net8686),
    .A2(_08980_));
 sg13g2_a221oi_1 _31974_ (.B2(_14002_),
    .C1(_08981_),
    .B1(net8582),
    .A1(_12906_),
    .Y(_08982_),
    .A2(net8603));
 sg13g2_o21ai_1 _31975_ (.B1(net9342),
    .Y(_08983_),
    .A1(net5407),
    .A2(net8319));
 sg13g2_nor2_1 _31976_ (.A(_08982_),
    .B(_08983_),
    .Y(_02532_));
 sg13g2_nand2b_1 _31977_ (.Y(_08984_),
    .B(net9260),
    .A_N(\soc_I.qqspi_I.spi_buf[8] ));
 sg13g2_o21ai_1 _31978_ (.B1(_08984_),
    .Y(_08985_),
    .A1(\soc_I.qqspi_I.spi_buf[11] ),
    .A2(net9260));
 sg13g2_o21ai_1 _31979_ (.B1(net8320),
    .Y(_08986_),
    .A1(net8687),
    .A2(_08985_));
 sg13g2_a221oi_1 _31980_ (.B2(_14006_),
    .C1(_08986_),
    .B1(_07186_),
    .A1(_12953_),
    .Y(_08987_),
    .A2(net8601));
 sg13g2_o21ai_1 _31981_ (.B1(net9337),
    .Y(_08988_),
    .A1(net5355),
    .A2(net8318));
 sg13g2_nor2_1 _31982_ (.A(_08987_),
    .B(_08988_),
    .Y(_02533_));
 sg13g2_nand2b_1 _31983_ (.Y(_08989_),
    .B(net9260),
    .A_N(\soc_I.qqspi_I.spi_buf[9] ));
 sg13g2_o21ai_1 _31984_ (.B1(_08989_),
    .Y(_08990_),
    .A1(\soc_I.qqspi_I.spi_buf[12] ),
    .A2(net9260));
 sg13g2_o21ai_1 _31985_ (.B1(net8321),
    .Y(_08991_),
    .A1(net8687),
    .A2(_08990_));
 sg13g2_a221oi_1 _31986_ (.B2(_14013_),
    .C1(_08991_),
    .B1(net8582),
    .A1(_12930_),
    .Y(_08992_),
    .A2(net8601));
 sg13g2_o21ai_1 _31987_ (.B1(net9338),
    .Y(_08993_),
    .A1(net5347),
    .A2(net8318));
 sg13g2_nor2_1 _31988_ (.A(_08992_),
    .B(_08993_),
    .Y(_02534_));
 sg13g2_nand2b_1 _31989_ (.Y(_08994_),
    .B(net9260),
    .A_N(\soc_I.qqspi_I.spi_buf[10] ));
 sg13g2_o21ai_1 _31990_ (.B1(_08994_),
    .Y(_08995_),
    .A1(\soc_I.qqspi_I.spi_buf[13] ),
    .A2(net9260));
 sg13g2_o21ai_1 _31991_ (.B1(net8320),
    .Y(_08996_),
    .A1(net8687),
    .A2(_08995_));
 sg13g2_a221oi_1 _31992_ (.B2(_14019_),
    .C1(_08996_),
    .B1(net8582),
    .A1(_12941_),
    .Y(_08997_),
    .A2(net8601));
 sg13g2_o21ai_1 _31993_ (.B1(net9338),
    .Y(_08998_),
    .A1(net5380),
    .A2(net8319));
 sg13g2_nor2_1 _31994_ (.A(_08997_),
    .B(_08998_),
    .Y(_02535_));
 sg13g2_nand2b_1 _31995_ (.Y(_08999_),
    .B(net9263),
    .A_N(\soc_I.qqspi_I.spi_buf[11] ));
 sg13g2_o21ai_1 _31996_ (.B1(_08999_),
    .Y(_09000_),
    .A1(\soc_I.qqspi_I.spi_buf[14] ),
    .A2(net9260));
 sg13g2_o21ai_1 _31997_ (.B1(net8320),
    .Y(_09001_),
    .A1(net8687),
    .A2(_09000_));
 sg13g2_a221oi_1 _31998_ (.B2(_14030_),
    .C1(_09001_),
    .B1(net8582),
    .A1(_12919_),
    .Y(_09002_),
    .A2(net8602));
 sg13g2_o21ai_1 _31999_ (.B1(net9337),
    .Y(_09003_),
    .A1(net5277),
    .A2(net8318));
 sg13g2_nor2_1 _32000_ (.A(_09002_),
    .B(_09003_),
    .Y(_02536_));
 sg13g2_and2_1 _32001_ (.A(net9707),
    .B(_07323_),
    .X(_09004_));
 sg13g2_nand2_1 _32002_ (.Y(_09005_),
    .A(net9707),
    .B(_07323_));
 sg13g2_a21oi_1 _32003_ (.A1(_14037_),
    .A2(net7469),
    .Y(_09006_),
    .B1(_07187_));
 sg13g2_o21ai_1 _32004_ (.B1(_09006_),
    .Y(_09007_),
    .A1(_13977_),
    .A2(net7469));
 sg13g2_mux2_1 _32005_ (.A0(\soc_I.qqspi_I.spi_buf[15] ),
    .A1(\soc_I.qqspi_I.spi_buf[12] ),
    .S(net9261),
    .X(_09008_));
 sg13g2_a22oi_1 _32006_ (.Y(_09009_),
    .B1(_09008_),
    .B2(net8682),
    .A2(net8601),
    .A1(_13008_));
 sg13g2_nand3_1 _32007_ (.B(_09007_),
    .C(_09009_),
    .A(net8320),
    .Y(_09010_));
 sg13g2_o21ai_1 _32008_ (.B1(_09010_),
    .Y(_09011_),
    .A1(net5273),
    .A2(net8318));
 sg13g2_nor2_1 _32009_ (.A(net9021),
    .B(_09011_),
    .Y(_02537_));
 sg13g2_nand2b_1 _32010_ (.Y(_09012_),
    .B(net9261),
    .A_N(\soc_I.qqspi_I.spi_buf[13] ));
 sg13g2_o21ai_1 _32011_ (.B1(_09012_),
    .Y(_09013_),
    .A1(\soc_I.qqspi_I.spi_buf[16] ),
    .A2(net9262));
 sg13g2_o21ai_1 _32012_ (.B1(net8321),
    .Y(_09014_),
    .A1(net8688),
    .A2(_09013_));
 sg13g2_nand2_1 _32013_ (.Y(_09015_),
    .A(net8613),
    .B(_09004_));
 sg13g2_a21oi_1 _32014_ (.A1(_14041_),
    .A2(net7469),
    .Y(_09016_),
    .B1(_07187_));
 sg13g2_a221oi_1 _32015_ (.B2(_09016_),
    .C1(_09014_),
    .B1(_09015_),
    .A1(_12977_),
    .Y(_09017_),
    .A2(net8601));
 sg13g2_o21ai_1 _32016_ (.B1(net9337),
    .Y(_09018_),
    .A1(net5300),
    .A2(net8318));
 sg13g2_nor2_1 _32017_ (.A(_09017_),
    .B(_09018_),
    .Y(_02538_));
 sg13g2_nand2_1 _32018_ (.Y(_09019_),
    .A(net8611),
    .B(_09004_));
 sg13g2_a21oi_1 _32019_ (.A1(_14046_),
    .A2(net7469),
    .Y(_09020_),
    .B1(_07187_));
 sg13g2_nand2b_1 _32020_ (.Y(_09021_),
    .B(net9261),
    .A_N(\soc_I.qqspi_I.spi_buf[14] ));
 sg13g2_o21ai_1 _32021_ (.B1(_09021_),
    .Y(_09022_),
    .A1(\soc_I.qqspi_I.spi_buf[17] ),
    .A2(net9261));
 sg13g2_o21ai_1 _32022_ (.B1(net8320),
    .Y(_09023_),
    .A1(net8688),
    .A2(_09022_));
 sg13g2_a221oi_1 _32023_ (.B2(_09020_),
    .C1(_09023_),
    .B1(_09019_),
    .A1(_13030_),
    .Y(_09024_),
    .A2(net8601));
 sg13g2_o21ai_1 _32024_ (.B1(net9338),
    .Y(_09025_),
    .A1(net5286),
    .A2(net8320));
 sg13g2_nor2_1 _32025_ (.A(_09024_),
    .B(_09025_),
    .Y(_02539_));
 sg13g2_nand2b_1 _32026_ (.Y(_09026_),
    .B(net9261),
    .A_N(\soc_I.qqspi_I.spi_buf[15] ));
 sg13g2_o21ai_1 _32027_ (.B1(_09026_),
    .Y(_09027_),
    .A1(\soc_I.qqspi_I.spi_buf[18] ),
    .A2(net9261));
 sg13g2_o21ai_1 _32028_ (.B1(net8321),
    .Y(_09028_),
    .A1(net8687),
    .A2(_09027_));
 sg13g2_a221oi_1 _32029_ (.B2(_14050_),
    .C1(_09028_),
    .B1(net8582),
    .A1(_12987_),
    .Y(_09029_),
    .A2(net8601));
 sg13g2_o21ai_1 _32030_ (.B1(net9338),
    .Y(_09030_),
    .A1(net5351),
    .A2(net8318));
 sg13g2_nor2_1 _32031_ (.A(_09029_),
    .B(_09030_),
    .Y(_02540_));
 sg13g2_nand2_1 _32032_ (.Y(_09031_),
    .A(net8609),
    .B(_09004_));
 sg13g2_a21oi_1 _32033_ (.A1(_14056_),
    .A2(net7469),
    .Y(_09032_),
    .B1(_07187_));
 sg13g2_nand2b_1 _32034_ (.Y(_09033_),
    .B(net9262),
    .A_N(\soc_I.qqspi_I.spi_buf[16] ));
 sg13g2_o21ai_1 _32035_ (.B1(_09033_),
    .Y(_09034_),
    .A1(\soc_I.qqspi_I.spi_buf[19] ),
    .A2(net9262));
 sg13g2_o21ai_1 _32036_ (.B1(net8320),
    .Y(_09035_),
    .A1(net8687),
    .A2(_09034_));
 sg13g2_a221oi_1 _32037_ (.B2(_09032_),
    .C1(_09035_),
    .B1(_09031_),
    .A1(_13041_),
    .Y(_09036_),
    .A2(net8601));
 sg13g2_o21ai_1 _32038_ (.B1(net9337),
    .Y(_09037_),
    .A1(net5406),
    .A2(net8318));
 sg13g2_nor2_1 _32039_ (.A(_09036_),
    .B(_09037_),
    .Y(_02541_));
 sg13g2_nand2_1 _32040_ (.Y(_09038_),
    .A(net8607),
    .B(_09004_));
 sg13g2_a21oi_1 _32041_ (.A1(_14060_),
    .A2(net7469),
    .Y(_09039_),
    .B1(_07187_));
 sg13g2_nand2b_1 _32042_ (.Y(_09040_),
    .B(net9261),
    .A_N(\soc_I.qqspi_I.spi_buf[17] ));
 sg13g2_o21ai_1 _32043_ (.B1(_09040_),
    .Y(_09041_),
    .A1(\soc_I.qqspi_I.spi_buf[20] ),
    .A2(net9261));
 sg13g2_o21ai_1 _32044_ (.B1(net8320),
    .Y(_09042_),
    .A1(net8687),
    .A2(_09041_));
 sg13g2_a221oi_1 _32045_ (.B2(_09039_),
    .C1(_09042_),
    .B1(_09038_),
    .A1(_13019_),
    .Y(_09043_),
    .A2(net8602));
 sg13g2_o21ai_1 _32046_ (.B1(net9344),
    .Y(_09044_),
    .A1(net5485),
    .A2(net8318));
 sg13g2_nor2_1 _32047_ (.A(_09043_),
    .B(_09044_),
    .Y(_02542_));
 sg13g2_nand2_1 _32048_ (.Y(_09045_),
    .A(net8605),
    .B(_09004_));
 sg13g2_a21oi_1 _32049_ (.A1(_14065_),
    .A2(_09005_),
    .Y(_09046_),
    .B1(_07187_));
 sg13g2_nand2b_1 _32050_ (.Y(_09047_),
    .B(net9262),
    .A_N(\soc_I.qqspi_I.spi_buf[18] ));
 sg13g2_o21ai_1 _32051_ (.B1(_09047_),
    .Y(_09048_),
    .A1(\soc_I.qqspi_I.spi_buf[21] ),
    .A2(net9262));
 sg13g2_o21ai_1 _32052_ (.B1(net8321),
    .Y(_09049_),
    .A1(net8687),
    .A2(_09048_));
 sg13g2_a221oi_1 _32053_ (.B2(_09046_),
    .C1(_09049_),
    .B1(_09045_),
    .A1(_12966_),
    .Y(_09050_),
    .A2(net8603));
 sg13g2_o21ai_1 _32054_ (.B1(net9344),
    .Y(_09051_),
    .A1(net5419),
    .A2(net8319));
 sg13g2_nor2_1 _32055_ (.A(_09050_),
    .B(_09051_),
    .Y(_02543_));
 sg13g2_a21oi_1 _32056_ (.A1(_14070_),
    .A2(net7469),
    .Y(_09052_),
    .B1(_07187_));
 sg13g2_o21ai_1 _32057_ (.B1(_09052_),
    .Y(_09053_),
    .A1(_14025_),
    .A2(net7469));
 sg13g2_mux2_1 _32058_ (.A0(\soc_I.qqspi_I.spi_buf[22] ),
    .A1(\soc_I.qqspi_I.spi_buf[19] ),
    .S(net9260),
    .X(_09054_));
 sg13g2_a221oi_1 _32059_ (.B2(net8680),
    .C1(_08963_),
    .B1(_09054_),
    .A1(_12998_),
    .Y(_09055_),
    .A2(net8602));
 sg13g2_a221oi_1 _32060_ (.B2(_09055_),
    .C1(net9021),
    .B1(_09053_),
    .A1(_10375_),
    .Y(_02544_),
    .A2(_08963_));
 sg13g2_nor2_1 _32061_ (.A(_14273_),
    .B(_08961_),
    .Y(_09056_));
 sg13g2_nor2b_1 _32062_ (.A(net9256),
    .B_N(net11),
    .Y(_09057_));
 sg13g2_a21oi_1 _32063_ (.A1(net9256),
    .A2(net10),
    .Y(_09058_),
    .B1(_09057_));
 sg13g2_nor2_1 _32064_ (.A(net8685),
    .B(_09058_),
    .Y(_09059_));
 sg13g2_a21oi_1 _32065_ (.A1(net8685),
    .A2(_13977_),
    .Y(_09060_),
    .B1(_09059_));
 sg13g2_o21ai_1 _32066_ (.B1(net9341),
    .Y(_09061_),
    .A1(net5466),
    .A2(net8317));
 sg13g2_a21oi_1 _32067_ (.A1(net8317),
    .A2(_09060_),
    .Y(_02545_),
    .B1(_09061_));
 sg13g2_mux2_1 _32068_ (.A0(\soc_I.qqspi_I.spi_buf[0] ),
    .A1(net11),
    .S(net9256),
    .X(_09062_));
 sg13g2_nor2_1 _32069_ (.A(net8677),
    .B(net8613),
    .Y(_09063_));
 sg13g2_a21oi_1 _32070_ (.A1(net8677),
    .A2(_09062_),
    .Y(_09064_),
    .B1(_09063_));
 sg13g2_o21ai_1 _32071_ (.B1(net9341),
    .Y(_09065_),
    .A1(net5468),
    .A2(net8317));
 sg13g2_a21oi_1 _32072_ (.A1(net8317),
    .A2(_09064_),
    .Y(_02546_),
    .B1(_09065_));
 sg13g2_mux2_1 _32073_ (.A0(\soc_I.qqspi_I.spi_buf[1] ),
    .A1(net12),
    .S(net9256),
    .X(_09066_));
 sg13g2_nor2_1 _32074_ (.A(net8677),
    .B(net8611),
    .Y(_09067_));
 sg13g2_a21oi_1 _32075_ (.A1(net8677),
    .A2(_09066_),
    .Y(_09068_),
    .B1(_09067_));
 sg13g2_o21ai_1 _32076_ (.B1(net9341),
    .Y(_09069_),
    .A1(net5459),
    .A2(net8317));
 sg13g2_a21oi_1 _32077_ (.A1(net8317),
    .A2(_09068_),
    .Y(_02547_),
    .B1(_09069_));
 sg13g2_mux2_1 _32078_ (.A0(\soc_I.qqspi_I.spi_buf[2] ),
    .A1(net13),
    .S(net9256),
    .X(_09070_));
 sg13g2_nor2_1 _32079_ (.A(net8677),
    .B(net8550),
    .Y(_09071_));
 sg13g2_a21oi_1 _32080_ (.A1(net8677),
    .A2(_09070_),
    .Y(_09072_),
    .B1(_09071_));
 sg13g2_o21ai_1 _32081_ (.B1(net9341),
    .Y(_09073_),
    .A1(net5413),
    .A2(net8317));
 sg13g2_a21oi_1 _32082_ (.A1(net8317),
    .A2(_09072_),
    .Y(_02548_),
    .B1(_09073_));
 sg13g2_mux2_1 _32083_ (.A0(\soc_I.qqspi_I.spi_buf[3] ),
    .A1(\soc_I.qqspi_I.spi_buf[0] ),
    .S(net9255),
    .X(_09074_));
 sg13g2_nor2_1 _32084_ (.A(net8679),
    .B(net8609),
    .Y(_09075_));
 sg13g2_a21oi_1 _32085_ (.A1(net8679),
    .A2(_09074_),
    .Y(_09076_),
    .B1(_09075_));
 sg13g2_o21ai_1 _32086_ (.B1(net9344),
    .Y(_09077_),
    .A1(net5287),
    .A2(net8316));
 sg13g2_a21oi_1 _32087_ (.A1(net8316),
    .A2(_09076_),
    .Y(_02549_),
    .B1(_09077_));
 sg13g2_mux2_1 _32088_ (.A0(\soc_I.qqspi_I.spi_buf[4] ),
    .A1(\soc_I.qqspi_I.spi_buf[1] ),
    .S(net9255),
    .X(_09078_));
 sg13g2_nor2_1 _32089_ (.A(net8679),
    .B(net8607),
    .Y(_09079_));
 sg13g2_a21oi_1 _32090_ (.A1(net8679),
    .A2(_09078_),
    .Y(_09080_),
    .B1(_09079_));
 sg13g2_o21ai_1 _32091_ (.B1(net9342),
    .Y(_09081_),
    .A1(net5198),
    .A2(net8316));
 sg13g2_a21oi_1 _32092_ (.A1(net8316),
    .A2(_09080_),
    .Y(_02550_),
    .B1(_09081_));
 sg13g2_mux2_1 _32093_ (.A0(\soc_I.qqspi_I.spi_buf[5] ),
    .A1(\soc_I.qqspi_I.spi_buf[2] ),
    .S(net9257),
    .X(_09082_));
 sg13g2_nor2_1 _32094_ (.A(net8679),
    .B(net8605),
    .Y(_09083_));
 sg13g2_a21oi_1 _32095_ (.A1(net8679),
    .A2(_09082_),
    .Y(_09084_),
    .B1(_09083_));
 sg13g2_o21ai_1 _32096_ (.B1(net9339),
    .Y(_09085_),
    .A1(net5320),
    .A2(net8316));
 sg13g2_a21oi_1 _32097_ (.A1(net8316),
    .A2(_09084_),
    .Y(_02551_),
    .B1(_09085_));
 sg13g2_nor2b_1 _32098_ (.A(net9255),
    .B_N(\soc_I.qqspi_I.spi_buf[6] ),
    .Y(_09086_));
 sg13g2_a21oi_1 _32099_ (.A1(\soc_I.qqspi_I.spi_buf[3] ),
    .A2(net9255),
    .Y(_09087_),
    .B1(_09086_));
 sg13g2_nor2_1 _32100_ (.A(net8686),
    .B(_09087_),
    .Y(_09088_));
 sg13g2_a21oi_1 _32101_ (.A1(net8686),
    .A2(_14025_),
    .Y(_09089_),
    .B1(_09088_));
 sg13g2_o21ai_1 _32102_ (.B1(net9339),
    .Y(_09090_),
    .A1(net5348),
    .A2(net8316));
 sg13g2_a21oi_1 _32103_ (.A1(net8316),
    .A2(_09089_),
    .Y(_02552_),
    .B1(_09090_));
 sg13g2_nand2_2 _32104_ (.Y(_09091_),
    .A(_14199_),
    .B(_06463_));
 sg13g2_nand2_1 _32105_ (.Y(_09092_),
    .A(net2679),
    .B(net8028));
 sg13g2_o21ai_1 _32106_ (.B1(_09092_),
    .Y(_02553_),
    .A1(net7485),
    .A2(net8028));
 sg13g2_nand2_1 _32107_ (.Y(_09093_),
    .A(net3119),
    .B(net8026));
 sg13g2_o21ai_1 _32108_ (.B1(_09093_),
    .Y(_02554_),
    .A1(net7665),
    .A2(net8026));
 sg13g2_nand2_1 _32109_ (.Y(_09094_),
    .A(net3768),
    .B(net8026));
 sg13g2_o21ai_1 _32110_ (.B1(_09094_),
    .Y(_02555_),
    .A1(net7615),
    .A2(net8026));
 sg13g2_nand2_1 _32111_ (.Y(_09095_),
    .A(net3439),
    .B(net8025));
 sg13g2_o21ai_1 _32112_ (.B1(_09095_),
    .Y(_02556_),
    .A1(net7607),
    .A2(net8025));
 sg13g2_nand2_1 _32113_ (.Y(_09096_),
    .A(net3380),
    .B(net8028));
 sg13g2_o21ai_1 _32114_ (.B1(_09096_),
    .Y(_02557_),
    .A1(net7587),
    .A2(net8028));
 sg13g2_nand2_1 _32115_ (.Y(_09097_),
    .A(net3140),
    .B(net8024));
 sg13g2_o21ai_1 _32116_ (.B1(_09097_),
    .Y(_02558_),
    .A1(net7597),
    .A2(net8024));
 sg13g2_nand2_1 _32117_ (.Y(_09098_),
    .A(net2936),
    .B(net8027));
 sg13g2_o21ai_1 _32118_ (.B1(_09098_),
    .Y(_02559_),
    .A1(net7593),
    .A2(net8027));
 sg13g2_nand2_1 _32119_ (.Y(_09099_),
    .A(net3765),
    .B(net8022));
 sg13g2_o21ai_1 _32120_ (.B1(_09099_),
    .Y(_02560_),
    .A1(net7604),
    .A2(net8022));
 sg13g2_nand2_1 _32121_ (.Y(_09100_),
    .A(net3732),
    .B(net8029));
 sg13g2_o21ai_1 _32122_ (.B1(_09100_),
    .Y(_02561_),
    .A1(net7561),
    .A2(net8029));
 sg13g2_nand2_1 _32123_ (.Y(_09101_),
    .A(net2942),
    .B(net8025));
 sg13g2_o21ai_1 _32124_ (.B1(_09101_),
    .Y(_02562_),
    .A1(net7576),
    .A2(net8025));
 sg13g2_nand2_1 _32125_ (.Y(_09102_),
    .A(net3156),
    .B(net8027));
 sg13g2_o21ai_1 _32126_ (.B1(_09102_),
    .Y(_02563_),
    .A1(net7546),
    .A2(net8027));
 sg13g2_nand2_1 _32127_ (.Y(_09103_),
    .A(net2956),
    .B(net8020));
 sg13g2_o21ai_1 _32128_ (.B1(_09103_),
    .Y(_02564_),
    .A1(net7570),
    .A2(net8020));
 sg13g2_nand2_1 _32129_ (.Y(_09104_),
    .A(net3704),
    .B(net8027));
 sg13g2_o21ai_1 _32130_ (.B1(_09104_),
    .Y(_02565_),
    .A1(net7540),
    .A2(net8027));
 sg13g2_nand2_1 _32131_ (.Y(_09105_),
    .A(net3733),
    .B(net8027));
 sg13g2_o21ai_1 _32132_ (.B1(_09105_),
    .Y(_02566_),
    .A1(net7551),
    .A2(net8027));
 sg13g2_nand2_1 _32133_ (.Y(_09106_),
    .A(net3822),
    .B(net8023));
 sg13g2_o21ai_1 _32134_ (.B1(_09106_),
    .Y(_02567_),
    .A1(net7580),
    .A2(net8023));
 sg13g2_nand2_1 _32135_ (.Y(_09107_),
    .A(net3507),
    .B(net8021));
 sg13g2_o21ai_1 _32136_ (.B1(_09107_),
    .Y(_02568_),
    .A1(net7566),
    .A2(net8021));
 sg13g2_nand2_1 _32137_ (.Y(_09108_),
    .A(net3601),
    .B(net8020));
 sg13g2_o21ai_1 _32138_ (.B1(_09108_),
    .Y(_02569_),
    .A1(net7524),
    .A2(net8020));
 sg13g2_nand2_1 _32139_ (.Y(_09109_),
    .A(net3083),
    .B(net8020));
 sg13g2_o21ai_1 _32140_ (.B1(_09109_),
    .Y(_02570_),
    .A1(net7537),
    .A2(net8020));
 sg13g2_nand2_1 _32141_ (.Y(_09110_),
    .A(net3561),
    .B(net8021));
 sg13g2_o21ai_1 _32142_ (.B1(_09110_),
    .Y(_02571_),
    .A1(net7530),
    .A2(net8021));
 sg13g2_nand2_1 _32143_ (.Y(_09111_),
    .A(net3896),
    .B(net8021));
 sg13g2_o21ai_1 _32144_ (.B1(_09111_),
    .Y(_02572_),
    .A1(net7518),
    .A2(net8021));
 sg13g2_nand2_1 _32145_ (.Y(_09112_),
    .A(net3742),
    .B(net8028));
 sg13g2_o21ai_1 _32146_ (.B1(_09112_),
    .Y(_02573_),
    .A1(net7504),
    .A2(net8028));
 sg13g2_nand2_1 _32147_ (.Y(_09113_),
    .A(net3863),
    .B(net8024));
 sg13g2_o21ai_1 _32148_ (.B1(_09113_),
    .Y(_02574_),
    .A1(net7512),
    .A2(net8024));
 sg13g2_nand2_1 _32149_ (.Y(_09114_),
    .A(net2979),
    .B(net8025));
 sg13g2_o21ai_1 _32150_ (.B1(_09114_),
    .Y(_02575_),
    .A1(net7494),
    .A2(net8025));
 sg13g2_nand2_1 _32151_ (.Y(_09115_),
    .A(net3668),
    .B(net8020));
 sg13g2_o21ai_1 _32152_ (.B1(_09115_),
    .Y(_02576_),
    .A1(net7503),
    .A2(net8020));
 sg13g2_nand2_1 _32153_ (.Y(_09116_),
    .A(net3508),
    .B(net8024));
 sg13g2_o21ai_1 _32154_ (.B1(_09116_),
    .Y(_02577_),
    .A1(net7646),
    .A2(net8024));
 sg13g2_nand2_1 _32155_ (.Y(_09117_),
    .A(net3154),
    .B(net8028));
 sg13g2_o21ai_1 _32156_ (.B1(_09117_),
    .Y(_02578_),
    .A1(net7648),
    .A2(net8028));
 sg13g2_nand2_1 _32157_ (.Y(_09118_),
    .A(net3367),
    .B(net8025));
 sg13g2_o21ai_1 _32158_ (.B1(_09118_),
    .Y(_02579_),
    .A1(net7657),
    .A2(net8025));
 sg13g2_nand2_1 _32159_ (.Y(_09119_),
    .A(net3727),
    .B(net8022));
 sg13g2_o21ai_1 _32160_ (.B1(_09119_),
    .Y(_02580_),
    .A1(net7660),
    .A2(net8022));
 sg13g2_nand2_1 _32161_ (.Y(_09120_),
    .A(net4007),
    .B(net8022));
 sg13g2_o21ai_1 _32162_ (.B1(_09120_),
    .Y(_02581_),
    .A1(net7636),
    .A2(net8022));
 sg13g2_nand2_1 _32163_ (.Y(_09121_),
    .A(net3475),
    .B(net8024));
 sg13g2_o21ai_1 _32164_ (.B1(_09121_),
    .Y(_02582_),
    .A1(net7626),
    .A2(net8024));
 sg13g2_nand2_1 _32165_ (.Y(_09122_),
    .A(net3618),
    .B(net8023));
 sg13g2_o21ai_1 _32166_ (.B1(_09122_),
    .Y(_02583_),
    .A1(net7621),
    .A2(net8023));
 sg13g2_nand2_1 _32167_ (.Y(_09123_),
    .A(net3686),
    .B(net8022));
 sg13g2_o21ai_1 _32168_ (.B1(_09123_),
    .Y(_02584_),
    .A1(net7630),
    .A2(net8021));
 sg13g2_nand2_1 _32169_ (.Y(_09124_),
    .A(_14126_),
    .B(_14370_));
 sg13g2_nand2_1 _32170_ (.Y(_09125_),
    .A(net3563),
    .B(net7817));
 sg13g2_o21ai_1 _32171_ (.B1(_09125_),
    .Y(_02585_),
    .A1(net7486),
    .A2(net7817));
 sg13g2_nand2_1 _32172_ (.Y(_09126_),
    .A(net3972),
    .B(net7818));
 sg13g2_o21ai_1 _32173_ (.B1(_09126_),
    .Y(_02586_),
    .A1(net7665),
    .A2(net7818));
 sg13g2_nand2_1 _32174_ (.Y(_09127_),
    .A(net2902),
    .B(net7818));
 sg13g2_o21ai_1 _32175_ (.B1(_09127_),
    .Y(_02587_),
    .A1(net7614),
    .A2(net7818));
 sg13g2_nand2_1 _32176_ (.Y(_09128_),
    .A(net3142),
    .B(net7819));
 sg13g2_o21ai_1 _32177_ (.B1(_09128_),
    .Y(_02588_),
    .A1(net7607),
    .A2(net7819));
 sg13g2_nand2_1 _32178_ (.Y(_09129_),
    .A(net3318),
    .B(net7817));
 sg13g2_o21ai_1 _32179_ (.B1(_09129_),
    .Y(_02589_),
    .A1(net7589),
    .A2(net7817));
 sg13g2_nand2_1 _32180_ (.Y(_09130_),
    .A(net3343),
    .B(net7822));
 sg13g2_o21ai_1 _32181_ (.B1(_09130_),
    .Y(_02590_),
    .A1(net7599),
    .A2(net7822));
 sg13g2_nand2_1 _32182_ (.Y(_09131_),
    .A(net3700),
    .B(net7820));
 sg13g2_o21ai_1 _32183_ (.B1(_09131_),
    .Y(_02591_),
    .A1(net7592),
    .A2(net7820));
 sg13g2_nand2_1 _32184_ (.Y(_09132_),
    .A(net3628),
    .B(net7815));
 sg13g2_o21ai_1 _32185_ (.B1(_09132_),
    .Y(_02592_),
    .A1(net7604),
    .A2(net7815));
 sg13g2_nand2_1 _32186_ (.Y(_09133_),
    .A(net3375),
    .B(net7822));
 sg13g2_o21ai_1 _32187_ (.B1(_09133_),
    .Y(_02593_),
    .A1(net7558),
    .A2(net7822));
 sg13g2_nand2_1 _32188_ (.Y(_09134_),
    .A(net2685),
    .B(net7820));
 sg13g2_o21ai_1 _32189_ (.B1(_09134_),
    .Y(_02594_),
    .A1(net7578),
    .A2(net7820));
 sg13g2_nand2_1 _32190_ (.Y(_09135_),
    .A(net2984),
    .B(net7819));
 sg13g2_o21ai_1 _32191_ (.B1(_09135_),
    .Y(_02595_),
    .A1(net7546),
    .A2(net7819));
 sg13g2_nand2_1 _32192_ (.Y(_09136_),
    .A(net4224),
    .B(net7813));
 sg13g2_o21ai_1 _32193_ (.B1(_09136_),
    .Y(_02596_),
    .A1(net7570),
    .A2(net7813));
 sg13g2_nand2_1 _32194_ (.Y(_09137_),
    .A(net3617),
    .B(net7820));
 sg13g2_o21ai_1 _32195_ (.B1(_09137_),
    .Y(_02597_),
    .A1(net7540),
    .A2(net7817));
 sg13g2_nand2_1 _32196_ (.Y(_09138_),
    .A(net3823),
    .B(net7820));
 sg13g2_o21ai_1 _32197_ (.B1(_09138_),
    .Y(_02598_),
    .A1(net7551),
    .A2(net7820));
 sg13g2_nand2_1 _32198_ (.Y(_09139_),
    .A(net3581),
    .B(net7815));
 sg13g2_o21ai_1 _32199_ (.B1(_09139_),
    .Y(_02599_),
    .A1(net7583),
    .A2(net7815));
 sg13g2_nand2_1 _32200_ (.Y(_09140_),
    .A(net3075),
    .B(net7814));
 sg13g2_o21ai_1 _32201_ (.B1(_09140_),
    .Y(_02600_),
    .A1(net7565),
    .A2(net7814));
 sg13g2_nand2_1 _32202_ (.Y(_09141_),
    .A(net3410),
    .B(net7813));
 sg13g2_o21ai_1 _32203_ (.B1(_09141_),
    .Y(_02601_),
    .A1(net7526),
    .A2(net7813));
 sg13g2_nand2_1 _32204_ (.Y(_09142_),
    .A(net2952),
    .B(net7813));
 sg13g2_o21ai_1 _32205_ (.B1(_09142_),
    .Y(_02602_),
    .A1(net7538),
    .A2(net7813));
 sg13g2_nand2_1 _32206_ (.Y(_09143_),
    .A(net4342),
    .B(net7813));
 sg13g2_o21ai_1 _32207_ (.B1(_09143_),
    .Y(_02603_),
    .A1(net7530),
    .A2(net7813));
 sg13g2_nand2_1 _32208_ (.Y(_09144_),
    .A(net3418),
    .B(net7815));
 sg13g2_o21ai_1 _32209_ (.B1(_09144_),
    .Y(_02604_),
    .A1(net7516),
    .A2(net7815));
 sg13g2_nand2_1 _32210_ (.Y(_09145_),
    .A(net3728),
    .B(net7817));
 sg13g2_o21ai_1 _32211_ (.B1(_09145_),
    .Y(_02605_),
    .A1(net7506),
    .A2(net7817));
 sg13g2_nand2_1 _32212_ (.Y(_09146_),
    .A(net2997),
    .B(net7823));
 sg13g2_o21ai_1 _32213_ (.B1(_09146_),
    .Y(_02606_),
    .A1(net7511),
    .A2(net7816));
 sg13g2_nand2_1 _32214_ (.Y(_09147_),
    .A(net3502),
    .B(net7818));
 sg13g2_o21ai_1 _32215_ (.B1(_09147_),
    .Y(_02607_),
    .A1(net7497),
    .A2(net7818));
 sg13g2_nand2_1 _32216_ (.Y(_09148_),
    .A(net3210),
    .B(net7814));
 sg13g2_o21ai_1 _32217_ (.B1(_09148_),
    .Y(_02608_),
    .A1(net7500),
    .A2(net7814));
 sg13g2_nand2_1 _32218_ (.Y(_09149_),
    .A(net3321),
    .B(net7822));
 sg13g2_o21ai_1 _32219_ (.B1(_09149_),
    .Y(_02609_),
    .A1(net7642),
    .A2(net7822));
 sg13g2_nand2_1 _32220_ (.Y(_09150_),
    .A(net3824),
    .B(net7821));
 sg13g2_o21ai_1 _32221_ (.B1(_09150_),
    .Y(_02610_),
    .A1(net7651),
    .A2(net7817));
 sg13g2_nand2_1 _32222_ (.Y(_09151_),
    .A(net3161),
    .B(net7818));
 sg13g2_o21ai_1 _32223_ (.B1(_09151_),
    .Y(_02611_),
    .A1(net7653),
    .A2(net7818));
 sg13g2_nand2_1 _32224_ (.Y(_09152_),
    .A(net3481),
    .B(net7816));
 sg13g2_o21ai_1 _32225_ (.B1(_09152_),
    .Y(_02612_),
    .A1(net7660),
    .A2(net7816));
 sg13g2_nand2_1 _32226_ (.Y(_09153_),
    .A(net3346),
    .B(net7816));
 sg13g2_o21ai_1 _32227_ (.B1(_09153_),
    .Y(_02613_),
    .A1(net7636),
    .A2(net7816));
 sg13g2_nand2_1 _32228_ (.Y(_09154_),
    .A(net3403),
    .B(net7822));
 sg13g2_o21ai_1 _32229_ (.B1(_09154_),
    .Y(_02614_),
    .A1(net7626),
    .A2(net7822));
 sg13g2_nand2_1 _32230_ (.Y(_09155_),
    .A(net3295),
    .B(net7816));
 sg13g2_o21ai_1 _32231_ (.B1(_09155_),
    .Y(_02615_),
    .A1(net7619),
    .A2(net7816));
 sg13g2_nand2_1 _32232_ (.Y(_09156_),
    .A(net2914),
    .B(net7814));
 sg13g2_o21ai_1 _32233_ (.B1(_09156_),
    .Y(_02616_),
    .A1(net7632),
    .A2(net7814));
 sg13g2_nand3_1 _32234_ (.B(_14126_),
    .C(net8372),
    .A(_12607_),
    .Y(_09157_));
 sg13g2_nand2_1 _32235_ (.Y(_09158_),
    .A(net2967),
    .B(net8018));
 sg13g2_o21ai_1 _32236_ (.B1(_09158_),
    .Y(_02649_),
    .A1(net7486),
    .A2(net8018));
 sg13g2_nand2_1 _32237_ (.Y(_09159_),
    .A(net3157),
    .B(net8018));
 sg13g2_o21ai_1 _32238_ (.B1(_09159_),
    .Y(_02650_),
    .A1(net7663),
    .A2(net8018));
 sg13g2_nand2_1 _32239_ (.Y(_09160_),
    .A(net2983),
    .B(net8018));
 sg13g2_o21ai_1 _32240_ (.B1(_09160_),
    .Y(_02651_),
    .A1(net7617),
    .A2(net8018));
 sg13g2_nand2_1 _32241_ (.Y(_09161_),
    .A(net3028),
    .B(net8016));
 sg13g2_o21ai_1 _32242_ (.B1(_09161_),
    .Y(_02652_),
    .A1(net7611),
    .A2(net8016));
 sg13g2_nand2_1 _32243_ (.Y(_09162_),
    .A(net3317),
    .B(net8014));
 sg13g2_o21ai_1 _32244_ (.B1(_09162_),
    .Y(_02653_),
    .A1(net7586),
    .A2(net8014));
 sg13g2_nand2_1 _32245_ (.Y(_09163_),
    .A(net2964),
    .B(net8013));
 sg13g2_o21ai_1 _32246_ (.B1(_09163_),
    .Y(_02654_),
    .A1(net7600),
    .A2(net8013));
 sg13g2_nand2_1 _32247_ (.Y(_09164_),
    .A(net3164),
    .B(net8015));
 sg13g2_o21ai_1 _32248_ (.B1(_09164_),
    .Y(_02655_),
    .A1(net7594),
    .A2(net8015));
 sg13g2_nand2_1 _32249_ (.Y(_09165_),
    .A(net2894),
    .B(net8009));
 sg13g2_o21ai_1 _32250_ (.B1(_09165_),
    .Y(_02656_),
    .A1(net7603),
    .A2(net8009));
 sg13g2_nand2_1 _32251_ (.Y(_09166_),
    .A(net3453),
    .B(net8014));
 sg13g2_o21ai_1 _32252_ (.B1(_09166_),
    .Y(_02657_),
    .A1(net7562),
    .A2(net8013));
 sg13g2_nand2_1 _32253_ (.Y(_09167_),
    .A(net2820),
    .B(net8017));
 sg13g2_o21ai_1 _32254_ (.B1(_09167_),
    .Y(_02658_),
    .A1(net7576),
    .A2(net8017));
 sg13g2_nand2_1 _32255_ (.Y(_09168_),
    .A(net3166),
    .B(net8015));
 sg13g2_o21ai_1 _32256_ (.B1(_09168_),
    .Y(_02659_),
    .A1(net7548),
    .A2(net8015));
 sg13g2_nand2_1 _32257_ (.Y(_09169_),
    .A(net3858),
    .B(net8009));
 sg13g2_o21ai_1 _32258_ (.B1(_09169_),
    .Y(_02660_),
    .A1(net7568),
    .A2(net8009));
 sg13g2_nand2_1 _32259_ (.Y(_09170_),
    .A(net3539),
    .B(net8015));
 sg13g2_o21ai_1 _32260_ (.B1(_09170_),
    .Y(_02661_),
    .A1(net7543),
    .A2(net8015));
 sg13g2_nand2_1 _32261_ (.Y(_09171_),
    .A(net3478),
    .B(net8017));
 sg13g2_o21ai_1 _32262_ (.B1(_09171_),
    .Y(_02662_),
    .A1(net7552),
    .A2(net8017));
 sg13g2_nand2_1 _32263_ (.Y(_09172_),
    .A(net3097),
    .B(net8012));
 sg13g2_o21ai_1 _32264_ (.B1(_09172_),
    .Y(_02663_),
    .A1(net7585),
    .A2(net8012));
 sg13g2_nand2_1 _32265_ (.Y(_09173_),
    .A(net2624),
    .B(net8010));
 sg13g2_o21ai_1 _32266_ (.B1(_09173_),
    .Y(_02664_),
    .A1(net7563),
    .A2(net8010));
 sg13g2_nand2_1 _32267_ (.Y(_09174_),
    .A(net3248),
    .B(net8009));
 sg13g2_o21ai_1 _32268_ (.B1(_09174_),
    .Y(_02665_),
    .A1(net7522),
    .A2(net8009));
 sg13g2_nand2_1 _32269_ (.Y(_09175_),
    .A(net2977),
    .B(net8009));
 sg13g2_o21ai_1 _32270_ (.B1(_09175_),
    .Y(_02666_),
    .A1(net7534),
    .A2(net8009));
 sg13g2_nand2_1 _32271_ (.Y(_09176_),
    .A(net3223),
    .B(net8010));
 sg13g2_o21ai_1 _32272_ (.B1(_09176_),
    .Y(_02667_),
    .A1(net7529),
    .A2(net8010));
 sg13g2_nand2_1 _32273_ (.Y(_09177_),
    .A(net3891),
    .B(net8011));
 sg13g2_o21ai_1 _32274_ (.B1(_09177_),
    .Y(_02668_),
    .A1(net7518),
    .A2(net8011));
 sg13g2_nand2_1 _32275_ (.Y(_09178_),
    .A(net3559),
    .B(net8014));
 sg13g2_o21ai_1 _32276_ (.B1(_09178_),
    .Y(_02669_),
    .A1(net7509),
    .A2(net8014));
 sg13g2_nand2_1 _32277_ (.Y(_09179_),
    .A(net3334),
    .B(net8013));
 sg13g2_o21ai_1 _32278_ (.B1(_09179_),
    .Y(_02670_),
    .A1(net7514),
    .A2(net8013));
 sg13g2_nand2_1 _32279_ (.Y(_09180_),
    .A(net3665),
    .B(net8016));
 sg13g2_o21ai_1 _32280_ (.B1(_09180_),
    .Y(_02671_),
    .A1(net7497),
    .A2(net8016));
 sg13g2_nand2_1 _32281_ (.Y(_09181_),
    .A(net3493),
    .B(net8010));
 sg13g2_o21ai_1 _32282_ (.B1(_09181_),
    .Y(_02672_),
    .A1(net7499),
    .A2(net8010));
 sg13g2_nand2_1 _32283_ (.Y(_09182_),
    .A(net3348),
    .B(net8013));
 sg13g2_o21ai_1 _32284_ (.B1(_09182_),
    .Y(_02673_),
    .A1(net7643),
    .A2(net8013));
 sg13g2_nand2_1 _32285_ (.Y(_09183_),
    .A(net3071),
    .B(net8018));
 sg13g2_o21ai_1 _32286_ (.B1(_09183_),
    .Y(_02674_),
    .A1(net7650),
    .A2(net8018));
 sg13g2_nand2_1 _32287_ (.Y(_09184_),
    .A(net3257),
    .B(net8015));
 sg13g2_o21ai_1 _32288_ (.B1(_09184_),
    .Y(_02675_),
    .A1(net7655),
    .A2(net8015));
 sg13g2_nand2_1 _32289_ (.Y(_09185_),
    .A(net3849),
    .B(net8011));
 sg13g2_o21ai_1 _32290_ (.B1(_09185_),
    .Y(_02676_),
    .A1(net7660),
    .A2(net8011));
 sg13g2_nand2_1 _32291_ (.Y(_09186_),
    .A(net2945),
    .B(net8011));
 sg13g2_o21ai_1 _32292_ (.B1(_09186_),
    .Y(_02677_),
    .A1(net7638),
    .A2(net8011));
 sg13g2_nand2_1 _32293_ (.Y(_09187_),
    .A(net2999),
    .B(net8014));
 sg13g2_o21ai_1 _32294_ (.B1(_09187_),
    .Y(_02678_),
    .A1(net7625),
    .A2(net8013));
 sg13g2_nand2_1 _32295_ (.Y(_09188_),
    .A(net3059),
    .B(net8011));
 sg13g2_o21ai_1 _32296_ (.B1(_09188_),
    .Y(_02679_),
    .A1(net7621),
    .A2(net8011));
 sg13g2_nand2_1 _32297_ (.Y(_09189_),
    .A(net2890),
    .B(net8012));
 sg13g2_o21ai_1 _32298_ (.B1(_09189_),
    .Y(_02680_),
    .A1(net7633),
    .A2(net8012));
 sg13g2_a21o_1 _32299_ (.A2(net8888),
    .A1(net8927),
    .B1(net9438),
    .X(_09190_));
 sg13g2_a21oi_1 _32300_ (.A1(net9143),
    .A2(_10695_),
    .Y(_09191_),
    .B1(net9168));
 sg13g2_o21ai_1 _32301_ (.B1(_09191_),
    .Y(_09192_),
    .A1(net9143),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][0] ));
 sg13g2_a22oi_1 _32302_ (.Y(_09193_),
    .B1(net8890),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][0] ),
    .A2(net8781),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][0] ));
 sg13g2_nand3_1 _32303_ (.B(_09192_),
    .C(_09193_),
    .A(net9468),
    .Y(_09194_));
 sg13g2_nor2_1 _32304_ (.A(net9536),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][0] ),
    .Y(_09195_));
 sg13g2_o21ai_1 _32305_ (.B1(net9499),
    .Y(_09196_),
    .A1(net9143),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][0] ));
 sg13g2_a221oi_1 _32306_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][0] ),
    .C1(net9468),
    .B1(net8890),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][0] ),
    .Y(_09197_),
    .A2(net8781));
 sg13g2_o21ai_1 _32307_ (.B1(_09197_),
    .Y(_09198_),
    .A1(_09195_),
    .A2(_09196_));
 sg13g2_and3_1 _32308_ (.X(_09199_),
    .A(net9449),
    .B(_09194_),
    .C(_09198_));
 sg13g2_nor2_1 _32309_ (.A(net9143),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][0] ),
    .Y(_09200_));
 sg13g2_o21ai_1 _32310_ (.B1(net9499),
    .Y(_09201_),
    .A1(net9536),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][0] ));
 sg13g2_a22oi_1 _32311_ (.Y(_09202_),
    .B1(net8890),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][0] ),
    .A2(net8781),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][0] ));
 sg13g2_o21ai_1 _32312_ (.B1(_09202_),
    .Y(_09203_),
    .A1(_09200_),
    .A2(_09201_));
 sg13g2_nor2_1 _32313_ (.A(net9533),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][0] ),
    .Y(_09204_));
 sg13g2_o21ai_1 _32314_ (.B1(net9497),
    .Y(_09205_),
    .A1(net9141),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][0] ));
 sg13g2_a22oi_1 _32315_ (.Y(_09206_),
    .B1(net8888),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][0] ),
    .A2(net8779),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][0] ));
 sg13g2_o21ai_1 _32316_ (.B1(_09206_),
    .Y(_09207_),
    .A1(_09204_),
    .A2(_09205_));
 sg13g2_a221oi_1 _32317_ (.B2(_08542_),
    .C1(_09199_),
    .B1(_09207_),
    .A1(net8927),
    .Y(_09208_),
    .A2(_09203_));
 sg13g2_a21oi_1 _32318_ (.A1(net9142),
    .A2(_10698_),
    .Y(_09209_),
    .B1(net9164));
 sg13g2_o21ai_1 _32319_ (.B1(_09209_),
    .Y(_09210_),
    .A1(net9142),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][0] ));
 sg13g2_a22oi_1 _32320_ (.Y(_09211_),
    .B1(net8888),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][0] ),
    .A2(net8779),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][0] ));
 sg13g2_nand3_1 _32321_ (.B(_09210_),
    .C(_09211_),
    .A(net9467),
    .Y(_09212_));
 sg13g2_nor2_1 _32322_ (.A(net9536),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][0] ),
    .Y(_09213_));
 sg13g2_o21ai_1 _32323_ (.B1(net9499),
    .Y(_09214_),
    .A1(net9141),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][0] ));
 sg13g2_a221oi_1 _32324_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][0] ),
    .C1(net9468),
    .B1(net8888),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][0] ),
    .Y(_09215_),
    .A2(net8779));
 sg13g2_o21ai_1 _32325_ (.B1(_09215_),
    .Y(_09216_),
    .A1(_09213_),
    .A2(_09214_));
 sg13g2_nand3_1 _32326_ (.B(_09212_),
    .C(_09216_),
    .A(net9449),
    .Y(_09217_));
 sg13g2_o21ai_1 _32327_ (.B1(net9496),
    .Y(_09218_),
    .A1(net9533),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][0] ));
 sg13g2_a21oi_1 _32328_ (.A1(net9532),
    .A2(_10696_),
    .Y(_09219_),
    .B1(_09218_));
 sg13g2_a221oi_1 _32329_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][0] ),
    .C1(_09219_),
    .B1(net8888),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][0] ),
    .Y(_09220_),
    .A2(net8779));
 sg13g2_nor2_1 _32330_ (.A(net8919),
    .B(_09220_),
    .Y(_09221_));
 sg13g2_o21ai_1 _32331_ (.B1(net9496),
    .Y(_09222_),
    .A1(net9533),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][0] ));
 sg13g2_a21oi_1 _32332_ (.A1(net9533),
    .A2(_10697_),
    .Y(_09223_),
    .B1(_09222_));
 sg13g2_a221oi_1 _32333_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][0] ),
    .C1(_09223_),
    .B1(net8888),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][0] ),
    .Y(_09224_),
    .A2(net8780));
 sg13g2_o21ai_1 _32334_ (.B1(_09217_),
    .Y(_09225_),
    .A1(net8915),
    .A2(_09224_));
 sg13g2_o21ai_1 _32335_ (.B1(net9438),
    .Y(_09226_),
    .A1(_09221_),
    .A2(_09225_));
 sg13g2_o21ai_1 _32336_ (.B1(_09226_),
    .Y(_02681_),
    .A1(net8747),
    .A2(_09208_));
 sg13g2_mux2_1 _32337_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][1] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][1] ),
    .S(net9535),
    .X(_09227_));
 sg13g2_a22oi_1 _32338_ (.Y(_09228_),
    .B1(net8892),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][1] ),
    .A2(net8783),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][1] ));
 sg13g2_nand2_1 _32339_ (.Y(_09229_),
    .A(net9468),
    .B(_09228_));
 sg13g2_a21oi_1 _32340_ (.A1(net9498),
    .A2(_09227_),
    .Y(_09230_),
    .B1(_09229_));
 sg13g2_a21oi_1 _32341_ (.A1(net9145),
    .A2(_10699_),
    .Y(_09231_),
    .B1(net9164));
 sg13g2_o21ai_1 _32342_ (.B1(_09231_),
    .Y(_09232_),
    .A1(net9145),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][1] ));
 sg13g2_a221oi_1 _32343_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][1] ),
    .C1(net9468),
    .B1(net8891),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][1] ),
    .Y(_09233_),
    .A2(net8782));
 sg13g2_a21oi_1 _32344_ (.A1(_09232_),
    .A2(_09233_),
    .Y(_09234_),
    .B1(_09230_));
 sg13g2_nor2_1 _32345_ (.A(net9535),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][1] ),
    .Y(_09235_));
 sg13g2_o21ai_1 _32346_ (.B1(net9498),
    .Y(_09236_),
    .A1(net9145),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][1] ));
 sg13g2_a22oi_1 _32347_ (.Y(_09237_),
    .B1(net8891),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][1] ),
    .A2(net8782),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][1] ));
 sg13g2_o21ai_1 _32348_ (.B1(_09237_),
    .Y(_09238_),
    .A1(_09235_),
    .A2(_09236_));
 sg13g2_mux2_1 _32349_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][1] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][1] ),
    .S(net9535),
    .X(_09239_));
 sg13g2_nand2_1 _32350_ (.Y(_09240_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][1] ),
    .B(net8891));
 sg13g2_a22oi_1 _32351_ (.Y(_09241_),
    .B1(_09239_),
    .B2(net9498),
    .A2(net8782),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][1] ));
 sg13g2_a21oi_1 _32352_ (.A1(_09240_),
    .A2(_09241_),
    .Y(_09242_),
    .B1(net8915));
 sg13g2_a221oi_1 _32353_ (.B2(net8927),
    .C1(_09242_),
    .B1(_09238_),
    .A1(net9449),
    .Y(_09243_),
    .A2(_09234_));
 sg13g2_nor2_1 _32354_ (.A(net9539),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][1] ),
    .Y(_09244_));
 sg13g2_o21ai_1 _32355_ (.B1(net9502),
    .Y(_09245_),
    .A1(net9148),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][1] ));
 sg13g2_a221oi_1 _32356_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][1] ),
    .C1(net9471),
    .B1(net8892),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][1] ),
    .Y(_09246_),
    .A2(net8783));
 sg13g2_o21ai_1 _32357_ (.B1(_09246_),
    .Y(_09247_),
    .A1(_09244_),
    .A2(_09245_));
 sg13g2_a21oi_1 _32358_ (.A1(net9148),
    .A2(_10702_),
    .Y(_09248_),
    .B1(net9167));
 sg13g2_o21ai_1 _32359_ (.B1(_09248_),
    .Y(_09249_),
    .A1(net9148),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][1] ));
 sg13g2_a22oi_1 _32360_ (.Y(_09250_),
    .B1(net8897),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][1] ),
    .A2(net8787),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][1] ));
 sg13g2_nand3_1 _32361_ (.B(_09249_),
    .C(_09250_),
    .A(net9471),
    .Y(_09251_));
 sg13g2_nand3_1 _32362_ (.B(_09247_),
    .C(_09251_),
    .A(net9448),
    .Y(_09252_));
 sg13g2_mux2_1 _32363_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][1] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][1] ),
    .S(net9535),
    .X(_09253_));
 sg13g2_nand2_1 _32364_ (.Y(_09254_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][1] ),
    .B(net8892));
 sg13g2_a22oi_1 _32365_ (.Y(_09255_),
    .B1(_09253_),
    .B2(net9500),
    .A2(net8783),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][1] ));
 sg13g2_a21oi_1 _32366_ (.A1(_09254_),
    .A2(_09255_),
    .Y(_09256_),
    .B1(net8919));
 sg13g2_o21ai_1 _32367_ (.B1(net9502),
    .Y(_09257_),
    .A1(net9148),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][1] ));
 sg13g2_a21oi_1 _32368_ (.A1(net9148),
    .A2(_10700_),
    .Y(_09258_),
    .B1(_09257_));
 sg13g2_a221oi_1 _32369_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][1] ),
    .C1(_09258_),
    .B1(net8897),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][1] ),
    .Y(_09259_),
    .A2(net8787));
 sg13g2_o21ai_1 _32370_ (.B1(_09252_),
    .Y(_09260_),
    .A1(net8913),
    .A2(_09259_));
 sg13g2_o21ai_1 _32371_ (.B1(net9438),
    .Y(_09261_),
    .A1(_09256_),
    .A2(_09260_));
 sg13g2_o21ai_1 _32372_ (.B1(_09261_),
    .Y(_02682_),
    .A1(net8747),
    .A2(_09243_));
 sg13g2_a21oi_1 _32373_ (.A1(net9143),
    .A2(_10703_),
    .Y(_09262_),
    .B1(net9164));
 sg13g2_o21ai_1 _32374_ (.B1(_09262_),
    .Y(_09263_),
    .A1(net9143),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][2] ));
 sg13g2_a22oi_1 _32375_ (.Y(_09264_),
    .B1(net8891),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][2] ),
    .A2(net8782),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][2] ));
 sg13g2_nand3_1 _32376_ (.B(_09263_),
    .C(_09264_),
    .A(net9469),
    .Y(_09265_));
 sg13g2_nor2_1 _32377_ (.A(net9535),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][2] ),
    .Y(_09266_));
 sg13g2_o21ai_1 _32378_ (.B1(net9498),
    .Y(_09267_),
    .A1(net9145),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][2] ));
 sg13g2_a221oi_1 _32379_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][2] ),
    .C1(net9468),
    .B1(net8891),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][2] ),
    .Y(_09268_),
    .A2(net8782));
 sg13g2_o21ai_1 _32380_ (.B1(_09268_),
    .Y(_09269_),
    .A1(_09266_),
    .A2(_09267_));
 sg13g2_and3_1 _32381_ (.X(_09270_),
    .A(net9449),
    .B(_09265_),
    .C(_09269_));
 sg13g2_nor2_1 _32382_ (.A(net9535),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][2] ),
    .Y(_09271_));
 sg13g2_o21ai_1 _32383_ (.B1(net9498),
    .Y(_09272_),
    .A1(net9145),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][2] ));
 sg13g2_a22oi_1 _32384_ (.Y(_09273_),
    .B1(net8891),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][2] ),
    .A2(net8782),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][2] ));
 sg13g2_o21ai_1 _32385_ (.B1(_09273_),
    .Y(_09274_),
    .A1(_09271_),
    .A2(_09272_));
 sg13g2_nor2_1 _32386_ (.A(net9535),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][2] ),
    .Y(_09275_));
 sg13g2_o21ai_1 _32387_ (.B1(net9498),
    .Y(_09276_),
    .A1(net9145),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][2] ));
 sg13g2_a22oi_1 _32388_ (.Y(_09277_),
    .B1(net8891),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][2] ),
    .A2(net8782),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][2] ));
 sg13g2_o21ai_1 _32389_ (.B1(_09277_),
    .Y(_09278_),
    .A1(_09275_),
    .A2(_09276_));
 sg13g2_a221oi_1 _32390_ (.B2(_08542_),
    .C1(_09270_),
    .B1(_09278_),
    .A1(net8927),
    .Y(_09279_),
    .A2(_09274_));
 sg13g2_nor2_1 _32391_ (.A(net9536),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][2] ),
    .Y(_09280_));
 sg13g2_o21ai_1 _32392_ (.B1(net9498),
    .Y(_09281_),
    .A1(net9146),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][2] ));
 sg13g2_a221oi_1 _32393_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][2] ),
    .C1(net9469),
    .B1(net8890),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][2] ),
    .Y(_09282_),
    .A2(net8781));
 sg13g2_o21ai_1 _32394_ (.B1(_09282_),
    .Y(_09283_),
    .A1(_09280_),
    .A2(_09281_));
 sg13g2_a21oi_1 _32395_ (.A1(net9146),
    .A2(_10706_),
    .Y(_09284_),
    .B1(net9164));
 sg13g2_o21ai_1 _32396_ (.B1(_09284_),
    .Y(_09285_),
    .A1(net9146),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][2] ));
 sg13g2_a22oi_1 _32397_ (.Y(_09286_),
    .B1(net8892),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][2] ),
    .A2(net8783),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][2] ));
 sg13g2_nand3_1 _32398_ (.B(_09285_),
    .C(_09286_),
    .A(net9469),
    .Y(_09287_));
 sg13g2_nand3_1 _32399_ (.B(_09283_),
    .C(_09287_),
    .A(net9449),
    .Y(_09288_));
 sg13g2_mux2_1 _32400_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][2] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][2] ),
    .S(net9535),
    .X(_09289_));
 sg13g2_nand2_1 _32401_ (.Y(_09290_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][2] ),
    .B(net8891));
 sg13g2_a22oi_1 _32402_ (.Y(_09291_),
    .B1(_09289_),
    .B2(net9498),
    .A2(net8783),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][2] ));
 sg13g2_a21oi_1 _32403_ (.A1(_09290_),
    .A2(_09291_),
    .Y(_09292_),
    .B1(net8919));
 sg13g2_o21ai_1 _32404_ (.B1(net9500),
    .Y(_09293_),
    .A1(net9145),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][2] ));
 sg13g2_a21oi_1 _32405_ (.A1(net9145),
    .A2(_10704_),
    .Y(_09294_),
    .B1(_09293_));
 sg13g2_a221oi_1 _32406_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][2] ),
    .C1(_09294_),
    .B1(net8892),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][2] ),
    .Y(_09295_),
    .A2(net8782));
 sg13g2_o21ai_1 _32407_ (.B1(_09288_),
    .Y(_09296_),
    .A1(net8915),
    .A2(_09295_));
 sg13g2_o21ai_1 _32408_ (.B1(net9438),
    .Y(_09297_),
    .A1(_09292_),
    .A2(_09296_));
 sg13g2_o21ai_1 _32409_ (.B1(_09297_),
    .Y(_02683_),
    .A1(net8746),
    .A2(_09279_));
 sg13g2_nor2_1 _32410_ (.A(net9539),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][3] ),
    .Y(_09298_));
 sg13g2_o21ai_1 _32411_ (.B1(net9503),
    .Y(_09299_),
    .A1(net9149),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][3] ));
 sg13g2_a221oi_1 _32412_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][3] ),
    .C1(net9471),
    .B1(net8897),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][3] ),
    .Y(_09300_),
    .A2(net8787));
 sg13g2_o21ai_1 _32413_ (.B1(_09300_),
    .Y(_09301_),
    .A1(_09298_),
    .A2(_09299_));
 sg13g2_a21oi_1 _32414_ (.A1(net9148),
    .A2(_10709_),
    .Y(_09302_),
    .B1(net9167));
 sg13g2_o21ai_1 _32415_ (.B1(_09302_),
    .Y(_09303_),
    .A1(net9148),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][3] ));
 sg13g2_a22oi_1 _32416_ (.Y(_09304_),
    .B1(net8898),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][3] ),
    .A2(net8788),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][3] ));
 sg13g2_nand3_1 _32417_ (.B(_09303_),
    .C(_09304_),
    .A(net9471),
    .Y(_09305_));
 sg13g2_nand3_1 _32418_ (.B(_09301_),
    .C(_09305_),
    .A(net9446),
    .Y(_09306_));
 sg13g2_nor2_1 _32419_ (.A(net9149),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][3] ),
    .Y(_09307_));
 sg13g2_o21ai_1 _32420_ (.B1(net9507),
    .Y(_09308_),
    .A1(net9542),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][3] ));
 sg13g2_a22oi_1 _32421_ (.Y(_09309_),
    .B1(net8898),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][3] ),
    .A2(net8788),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][3] ));
 sg13g2_o21ai_1 _32422_ (.B1(_09309_),
    .Y(_09310_),
    .A1(_09307_),
    .A2(_09308_));
 sg13g2_o21ai_1 _32423_ (.B1(net9502),
    .Y(_09311_),
    .A1(net9538),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][3] ));
 sg13g2_a21oi_1 _32424_ (.A1(net9538),
    .A2(_10708_),
    .Y(_09312_),
    .B1(_09311_));
 sg13g2_a221oi_1 _32425_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][3] ),
    .C1(_09312_),
    .B1(net8898),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][3] ),
    .Y(_09313_),
    .A2(net8788));
 sg13g2_o21ai_1 _32426_ (.B1(net9436),
    .Y(_09314_),
    .A1(net8913),
    .A2(_09313_));
 sg13g2_a21oi_1 _32427_ (.A1(net8926),
    .A2(_09310_),
    .Y(_09315_),
    .B1(_09314_));
 sg13g2_nor4_2 _32428_ (.A(net9436),
    .B(net9503),
    .C(net9538),
    .Y(_09316_),
    .D(net8920));
 sg13g2_nor2_1 _32429_ (.A(net9542),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][3] ),
    .Y(_09317_));
 sg13g2_o21ai_1 _32430_ (.B1(net9507),
    .Y(_09318_),
    .A1(net9153),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][3] ));
 sg13g2_a221oi_1 _32431_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][3] ),
    .C1(net9472),
    .B1(net8904),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][3] ),
    .Y(_09319_),
    .A2(net8793));
 sg13g2_o21ai_1 _32432_ (.B1(_09319_),
    .Y(_09320_),
    .A1(_09317_),
    .A2(_09318_));
 sg13g2_a21oi_1 _32433_ (.A1(net9156),
    .A2(_10707_),
    .Y(_09321_),
    .B1(net9165));
 sg13g2_o21ai_1 _32434_ (.B1(_09321_),
    .Y(_09322_),
    .A1(net9153),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][3] ));
 sg13g2_a22oi_1 _32435_ (.Y(_09323_),
    .B1(net8904),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][3] ),
    .A2(net8793),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][3] ));
 sg13g2_nand3_1 _32436_ (.B(_09322_),
    .C(_09323_),
    .A(net9472),
    .Y(_09324_));
 sg13g2_nand3_1 _32437_ (.B(_09320_),
    .C(_09324_),
    .A(net9448),
    .Y(_09325_));
 sg13g2_nor2_1 _32438_ (.A(net9542),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][3] ),
    .Y(_09326_));
 sg13g2_o21ai_1 _32439_ (.B1(net9507),
    .Y(_09327_),
    .A1(net9154),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][3] ));
 sg13g2_a22oi_1 _32440_ (.Y(_09328_),
    .B1(net8903),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][3] ),
    .A2(net8792),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][3] ));
 sg13g2_o21ai_1 _32441_ (.B1(_09328_),
    .Y(_09329_),
    .A1(_09326_),
    .A2(_09327_));
 sg13g2_nor2_1 _32442_ (.A(net9543),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][3] ),
    .Y(_09330_));
 sg13g2_o21ai_1 _32443_ (.B1(net9507),
    .Y(_09331_),
    .A1(net9154),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][3] ));
 sg13g2_a22oi_1 _32444_ (.Y(_09332_),
    .B1(net8903),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][3] ),
    .A2(net8792),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][3] ));
 sg13g2_o21ai_1 _32445_ (.B1(_09332_),
    .Y(_09333_),
    .A1(_09330_),
    .A2(_09331_));
 sg13g2_a221oi_1 _32446_ (.B2(net8926),
    .C1(net9437),
    .B1(_09333_),
    .A1(_08542_),
    .Y(_09334_),
    .A2(_09329_));
 sg13g2_a221oi_1 _32447_ (.B2(_09334_),
    .C1(_09316_),
    .B1(_09325_),
    .A1(_09306_),
    .Y(_02684_),
    .A2(_09315_));
 sg13g2_mux2_1 _32448_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][4] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][4] ),
    .S(net9532),
    .X(_09335_));
 sg13g2_a22oi_1 _32449_ (.Y(_09336_),
    .B1(net8885),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][4] ),
    .A2(net8776),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][4] ));
 sg13g2_nand2_1 _32450_ (.Y(_09337_),
    .A(net9467),
    .B(_09336_));
 sg13g2_a21oi_1 _32451_ (.A1(net9494),
    .A2(_09335_),
    .Y(_09338_),
    .B1(_09337_));
 sg13g2_a21oi_1 _32452_ (.A1(net9138),
    .A2(_10710_),
    .Y(_09339_),
    .B1(net9163));
 sg13g2_o21ai_1 _32453_ (.B1(_09339_),
    .Y(_09340_),
    .A1(net9139),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][4] ));
 sg13g2_a221oi_1 _32454_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][4] ),
    .C1(net9465),
    .B1(net8885),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][4] ),
    .Y(_09341_),
    .A2(net8776));
 sg13g2_a21oi_1 _32455_ (.A1(_09340_),
    .A2(_09341_),
    .Y(_09342_),
    .B1(_09338_));
 sg13g2_nor2_1 _32456_ (.A(net9531),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][4] ),
    .Y(_09343_));
 sg13g2_o21ai_1 _32457_ (.B1(net9493),
    .Y(_09344_),
    .A1(net9138),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][4] ));
 sg13g2_a22oi_1 _32458_ (.Y(_09345_),
    .B1(net8884),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][4] ),
    .A2(net8775),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][4] ));
 sg13g2_o21ai_1 _32459_ (.B1(_09345_),
    .Y(_09346_),
    .A1(_09343_),
    .A2(_09344_));
 sg13g2_mux2_1 _32460_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][4] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][4] ),
    .S(net9530),
    .X(_09347_));
 sg13g2_nand2_1 _32461_ (.Y(_09348_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][4] ),
    .B(net8884));
 sg13g2_a22oi_1 _32462_ (.Y(_09349_),
    .B1(_09347_),
    .B2(net9493),
    .A2(net8775),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][4] ));
 sg13g2_a21oi_1 _32463_ (.A1(_09348_),
    .A2(_09349_),
    .Y(_09350_),
    .B1(net8912));
 sg13g2_a221oi_1 _32464_ (.B2(net8925),
    .C1(_09350_),
    .B1(_09346_),
    .A1(net9445),
    .Y(_09351_),
    .A2(_09342_));
 sg13g2_a21oi_1 _32465_ (.A1(net9139),
    .A2(_10712_),
    .Y(_09352_),
    .B1(net9163));
 sg13g2_o21ai_1 _32466_ (.B1(_09352_),
    .Y(_09353_),
    .A1(net9139),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][4] ));
 sg13g2_a22oi_1 _32467_ (.Y(_09354_),
    .B1(net8885),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][4] ),
    .A2(net8776),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][4] ));
 sg13g2_nand3_1 _32468_ (.B(_09353_),
    .C(_09354_),
    .A(net9465),
    .Y(_09355_));
 sg13g2_nor2_1 _32469_ (.A(net9532),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][4] ),
    .Y(_09356_));
 sg13g2_o21ai_1 _32470_ (.B1(net9496),
    .Y(_09357_),
    .A1(net9141),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][4] ));
 sg13g2_a221oi_1 _32471_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][4] ),
    .C1(net9467),
    .B1(net8889),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][4] ),
    .Y(_09358_),
    .A2(net8779));
 sg13g2_o21ai_1 _32472_ (.B1(_09358_),
    .Y(_09359_),
    .A1(_09356_),
    .A2(_09357_));
 sg13g2_nand3_1 _32473_ (.B(_09355_),
    .C(_09359_),
    .A(net9445),
    .Y(_09360_));
 sg13g2_mux2_1 _32474_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][4] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][4] ),
    .S(net9530),
    .X(_09361_));
 sg13g2_nand2_1 _32475_ (.Y(_09362_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][4] ),
    .B(net8884));
 sg13g2_a22oi_1 _32476_ (.Y(_09363_),
    .B1(_09361_),
    .B2(net9493),
    .A2(net8775),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][4] ));
 sg13g2_a21oi_1 _32477_ (.A1(_09362_),
    .A2(_09363_),
    .Y(_09364_),
    .B1(net8921));
 sg13g2_o21ai_1 _32478_ (.B1(net9493),
    .Y(_09365_),
    .A1(net9138),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][4] ));
 sg13g2_a21oi_1 _32479_ (.A1(net9138),
    .A2(_10711_),
    .Y(_09366_),
    .B1(_09365_));
 sg13g2_a221oi_1 _32480_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][4] ),
    .C1(_09366_),
    .B1(net8884),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][4] ),
    .Y(_09367_),
    .A2(net8775));
 sg13g2_o21ai_1 _32481_ (.B1(_09360_),
    .Y(_09368_),
    .A1(net8912),
    .A2(_09367_));
 sg13g2_o21ai_1 _32482_ (.B1(net9439),
    .Y(_09369_),
    .A1(_09364_),
    .A2(_09368_));
 sg13g2_o21ai_1 _32483_ (.B1(_09369_),
    .Y(_02685_),
    .A1(net8747),
    .A2(_09351_));
 sg13g2_mux2_1 _32484_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][5] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][5] ),
    .S(net9525),
    .X(_09370_));
 sg13g2_a22oi_1 _32485_ (.Y(_09371_),
    .B1(net8880),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][5] ),
    .A2(net8769),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][5] ));
 sg13g2_nand2_1 _32486_ (.Y(_09372_),
    .A(net9463),
    .B(_09371_));
 sg13g2_a21oi_1 _32487_ (.A1(net9490),
    .A2(_09370_),
    .Y(_09373_),
    .B1(_09372_));
 sg13g2_mux2_1 _32488_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][5] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][5] ),
    .S(net9525),
    .X(_09374_));
 sg13g2_nand2_1 _32489_ (.Y(_09375_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][5] ),
    .B(net8880));
 sg13g2_a221oi_1 _32490_ (.B2(net9490),
    .C1(net9463),
    .B1(_09374_),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][5] ),
    .Y(_09376_),
    .A2(net8771));
 sg13g2_a21oi_1 _32491_ (.A1(_09375_),
    .A2(_09376_),
    .Y(_09377_),
    .B1(_09373_));
 sg13g2_nor2_1 _32492_ (.A(net9526),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][5] ),
    .Y(_09378_));
 sg13g2_o21ai_1 _32493_ (.B1(net9491),
    .Y(_09379_),
    .A1(net9135),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][5] ));
 sg13g2_a22oi_1 _32494_ (.Y(_09380_),
    .B1(net8881),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][5] ),
    .A2(net8772),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][5] ));
 sg13g2_o21ai_1 _32495_ (.B1(_09380_),
    .Y(_09381_),
    .A1(_09378_),
    .A2(_09379_));
 sg13g2_mux2_1 _32496_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][5] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][5] ),
    .S(net9526),
    .X(_09382_));
 sg13g2_nand2_1 _32497_ (.Y(_09383_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][5] ),
    .B(net8881));
 sg13g2_a22oi_1 _32498_ (.Y(_09384_),
    .B1(_09382_),
    .B2(net9491),
    .A2(net8772),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][5] ));
 sg13g2_a21oi_1 _32499_ (.A1(_09383_),
    .A2(_09384_),
    .Y(_09385_),
    .B1(net8911));
 sg13g2_a221oi_1 _32500_ (.B2(net8925),
    .C1(_09385_),
    .B1(_09381_),
    .A1(net9444),
    .Y(_09386_),
    .A2(_09377_));
 sg13g2_a21oi_1 _32501_ (.A1(net9134),
    .A2(_10714_),
    .Y(_09387_),
    .B1(net9163));
 sg13g2_o21ai_1 _32502_ (.B1(_09387_),
    .Y(_09388_),
    .A1(net9134),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][5] ));
 sg13g2_a22oi_1 _32503_ (.Y(_09389_),
    .B1(net8881),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][5] ),
    .A2(net8772),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][5] ));
 sg13g2_nand3_1 _32504_ (.B(_09388_),
    .C(_09389_),
    .A(net9463),
    .Y(_09390_));
 sg13g2_nor2_1 _32505_ (.A(net9526),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][5] ),
    .Y(_09391_));
 sg13g2_o21ai_1 _32506_ (.B1(net9490),
    .Y(_09392_),
    .A1(net9134),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][5] ));
 sg13g2_a221oi_1 _32507_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][5] ),
    .C1(net9463),
    .B1(net8881),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][5] ),
    .Y(_09393_),
    .A2(net8771));
 sg13g2_o21ai_1 _32508_ (.B1(_09393_),
    .Y(_09394_),
    .A1(_09391_),
    .A2(_09392_));
 sg13g2_nand3_1 _32509_ (.B(_09390_),
    .C(_09394_),
    .A(net9444),
    .Y(_09395_));
 sg13g2_mux2_1 _32510_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][5] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][5] ),
    .S(net9525),
    .X(_09396_));
 sg13g2_nand2_1 _32511_ (.Y(_09397_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][5] ),
    .B(net8878));
 sg13g2_a22oi_1 _32512_ (.Y(_09398_),
    .B1(_09396_),
    .B2(net9489),
    .A2(net8769),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][5] ));
 sg13g2_a21oi_1 _32513_ (.A1(_09397_),
    .A2(_09398_),
    .Y(_09399_),
    .B1(net8918));
 sg13g2_o21ai_1 _32514_ (.B1(net9490),
    .Y(_09400_),
    .A1(net9134),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][5] ));
 sg13g2_a21oi_1 _32515_ (.A1(net9134),
    .A2(_10713_),
    .Y(_09401_),
    .B1(_09400_));
 sg13g2_a221oi_1 _32516_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][5] ),
    .C1(_09401_),
    .B1(net8880),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][5] ),
    .Y(_09402_),
    .A2(net8771));
 sg13g2_o21ai_1 _32517_ (.B1(_09395_),
    .Y(_09403_),
    .A1(net8911),
    .A2(_09402_));
 sg13g2_o21ai_1 _32518_ (.B1(net9434),
    .Y(_09404_),
    .A1(_09399_),
    .A2(_09403_));
 sg13g2_o21ai_1 _32519_ (.B1(_09404_),
    .Y(_02686_),
    .A1(net8746),
    .A2(_09386_));
 sg13g2_a21oi_1 _32520_ (.A1(net9152),
    .A2(_10717_),
    .Y(_09405_),
    .B1(net9166));
 sg13g2_o21ai_1 _32521_ (.B1(_09405_),
    .Y(_09406_),
    .A1(net9152),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][6] ));
 sg13g2_a22oi_1 _32522_ (.Y(_09407_),
    .B1(net8902),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][6] ),
    .A2(net8791),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][6] ));
 sg13g2_nand3_1 _32523_ (.B(_09406_),
    .C(_09407_),
    .A(net9474),
    .Y(_09408_));
 sg13g2_nor2_1 _32524_ (.A(net9540),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][6] ),
    .Y(_09409_));
 sg13g2_o21ai_1 _32525_ (.B1(net9505),
    .Y(_09410_),
    .A1(net9152),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][6] ));
 sg13g2_a221oi_1 _32526_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][6] ),
    .C1(net9474),
    .B1(net8902),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][6] ),
    .Y(_09411_),
    .A2(net8791));
 sg13g2_o21ai_1 _32527_ (.B1(_09411_),
    .Y(_09412_),
    .A1(_09409_),
    .A2(_09410_));
 sg13g2_nand3_1 _32528_ (.B(_09408_),
    .C(_09412_),
    .A(net9447),
    .Y(_09413_));
 sg13g2_o21ai_1 _32529_ (.B1(net9505),
    .Y(_09414_),
    .A1(net9540),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][6] ));
 sg13g2_a21oi_1 _32530_ (.A1(net9540),
    .A2(_10716_),
    .Y(_09415_),
    .B1(_09414_));
 sg13g2_a221oi_1 _32531_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][6] ),
    .C1(_09415_),
    .B1(net8896),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][6] ),
    .Y(_09416_),
    .A2(net8785));
 sg13g2_nor2_1 _32532_ (.A(net9152),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][6] ),
    .Y(_09417_));
 sg13g2_o21ai_1 _32533_ (.B1(net9505),
    .Y(_09418_),
    .A1(net9540),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][6] ));
 sg13g2_a22oi_1 _32534_ (.Y(_09419_),
    .B1(net8902),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][6] ),
    .A2(net8791),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][6] ));
 sg13g2_o21ai_1 _32535_ (.B1(_09419_),
    .Y(_09420_),
    .A1(_09417_),
    .A2(_09418_));
 sg13g2_o21ai_1 _32536_ (.B1(net9437),
    .Y(_09421_),
    .A1(net8914),
    .A2(_09416_));
 sg13g2_a21oi_1 _32537_ (.A1(net8927),
    .A2(_09420_),
    .Y(_09422_),
    .B1(_09421_));
 sg13g2_nor2_1 _32538_ (.A(net9541),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][6] ),
    .Y(_09423_));
 sg13g2_o21ai_1 _32539_ (.B1(net9506),
    .Y(_09424_),
    .A1(net9151),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][6] ));
 sg13g2_a221oi_1 _32540_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][6] ),
    .C1(net9474),
    .B1(net8900),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][6] ),
    .Y(_09425_),
    .A2(net8791));
 sg13g2_o21ai_1 _32541_ (.B1(_09425_),
    .Y(_09426_),
    .A1(_09423_),
    .A2(_09424_));
 sg13g2_a21oi_1 _32542_ (.A1(net9151),
    .A2(_10715_),
    .Y(_09427_),
    .B1(net9166));
 sg13g2_o21ai_1 _32543_ (.B1(_09427_),
    .Y(_09428_),
    .A1(net9151),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][6] ));
 sg13g2_a22oi_1 _32544_ (.Y(_09429_),
    .B1(net8900),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][6] ),
    .A2(net8790),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][6] ));
 sg13g2_nand3_1 _32545_ (.B(_09428_),
    .C(_09429_),
    .A(net9474),
    .Y(_09430_));
 sg13g2_nand3_1 _32546_ (.B(_09426_),
    .C(_09430_),
    .A(net9447),
    .Y(_09431_));
 sg13g2_mux2_1 _32547_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][6] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][6] ),
    .S(net9541),
    .X(_09432_));
 sg13g2_nand2_1 _32548_ (.Y(_09433_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][6] ),
    .B(net8900));
 sg13g2_a22oi_1 _32549_ (.Y(_09434_),
    .B1(_09432_),
    .B2(net9506),
    .A2(net8790),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][6] ));
 sg13g2_a21oi_1 _32550_ (.A1(_09433_),
    .A2(_09434_),
    .Y(_09435_),
    .B1(net8914));
 sg13g2_mux2_1 _32551_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][6] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][6] ),
    .S(net9541),
    .X(_09436_));
 sg13g2_a22oi_1 _32552_ (.Y(_09437_),
    .B1(_09436_),
    .B2(net9505),
    .A2(net8790),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][6] ));
 sg13g2_nor3_1 _32553_ (.A(net8920),
    .B(net8900),
    .C(_09437_),
    .Y(_09438_));
 sg13g2_nor3_2 _32554_ (.A(net9437),
    .B(_09435_),
    .C(_09438_),
    .Y(_09439_));
 sg13g2_a22oi_1 _32555_ (.Y(_02687_),
    .B1(_09431_),
    .B2(_09439_),
    .A2(_09422_),
    .A1(_09413_));
 sg13g2_mux2_1 _32556_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][7] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][7] ),
    .S(net9511),
    .X(_09440_));
 sg13g2_a22oi_1 _32557_ (.Y(_09441_),
    .B1(net8862),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][7] ),
    .A2(net8751),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][7] ));
 sg13g2_nand2_1 _32558_ (.Y(_09442_),
    .A(net9452),
    .B(_09441_));
 sg13g2_a21oi_1 _32559_ (.A1(net9477),
    .A2(_09440_),
    .Y(_09443_),
    .B1(_09442_));
 sg13g2_a21oi_1 _32560_ (.A1(net9116),
    .A2(_10718_),
    .Y(_09444_),
    .B1(net9158));
 sg13g2_o21ai_1 _32561_ (.B1(_09444_),
    .Y(_09445_),
    .A1(net9116),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][7] ));
 sg13g2_a221oi_1 _32562_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][7] ),
    .C1(net9451),
    .B1(net8860),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][7] ),
    .Y(_09446_),
    .A2(net8749));
 sg13g2_a21oi_1 _32563_ (.A1(_09445_),
    .A2(_09446_),
    .Y(_09447_),
    .B1(_09443_));
 sg13g2_nor2_1 _32564_ (.A(net9510),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][7] ),
    .Y(_09448_));
 sg13g2_o21ai_1 _32565_ (.B1(net9476),
    .Y(_09449_),
    .A1(net9116),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][7] ));
 sg13g2_a22oi_1 _32566_ (.Y(_09450_),
    .B1(net8860),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][7] ),
    .A2(net8749),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][7] ));
 sg13g2_o21ai_1 _32567_ (.B1(_09450_),
    .Y(_09451_),
    .A1(_09448_),
    .A2(_09449_));
 sg13g2_mux2_1 _32568_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][7] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][7] ),
    .S(net9510),
    .X(_09452_));
 sg13g2_nand2_1 _32569_ (.Y(_09453_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][7] ),
    .B(net8860));
 sg13g2_a22oi_1 _32570_ (.Y(_09454_),
    .B1(_09452_),
    .B2(net9476),
    .A2(net8749),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][7] ));
 sg13g2_a21oi_1 _32571_ (.A1(_09453_),
    .A2(_09454_),
    .Y(_09455_),
    .B1(net8908));
 sg13g2_a221oi_1 _32572_ (.B2(net8922),
    .C1(_09455_),
    .B1(_09451_),
    .A1(net9440),
    .Y(_09456_),
    .A2(_09447_));
 sg13g2_a21oi_1 _32573_ (.A1(net9123),
    .A2(_10719_),
    .Y(_09457_),
    .B1(net9159));
 sg13g2_o21ai_1 _32574_ (.B1(_09457_),
    .Y(_09458_),
    .A1(net9123),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][7] ));
 sg13g2_a221oi_1 _32575_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][7] ),
    .C1(net9455),
    .B1(net8869),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][7] ),
    .Y(_09459_),
    .A2(net8759));
 sg13g2_o21ai_1 _32576_ (.B1(net9484),
    .Y(_09460_),
    .A1(net9518),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][7] ));
 sg13g2_a21oi_1 _32577_ (.A1(net9518),
    .A2(_10721_),
    .Y(_09461_),
    .B1(_09460_));
 sg13g2_a221oi_1 _32578_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][7] ),
    .C1(_09461_),
    .B1(net8869),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][7] ),
    .Y(_09462_),
    .A2(net8759));
 sg13g2_a22oi_1 _32579_ (.Y(_09463_),
    .B1(_09462_),
    .B2(net9455),
    .A2(_09459_),
    .A1(_09458_));
 sg13g2_nor2_1 _32580_ (.A(net9515),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][7] ),
    .Y(_09464_));
 sg13g2_o21ai_1 _32581_ (.B1(net9481),
    .Y(_09465_),
    .A1(net9122),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][7] ));
 sg13g2_a22oi_1 _32582_ (.Y(_09466_),
    .B1(net8866),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][7] ),
    .A2(net8757),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][7] ));
 sg13g2_o21ai_1 _32583_ (.B1(_09466_),
    .Y(_09467_),
    .A1(_09464_),
    .A2(_09465_));
 sg13g2_mux2_1 _32584_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][7] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][7] ),
    .S(net9515),
    .X(_09468_));
 sg13g2_nand2_1 _32585_ (.Y(_09469_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][7] ),
    .B(net8866));
 sg13g2_a22oi_1 _32586_ (.Y(_09470_),
    .B1(_09468_),
    .B2(net9481),
    .A2(net8757),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][7] ));
 sg13g2_a21oi_1 _32587_ (.A1(_09469_),
    .A2(_09470_),
    .Y(_09471_),
    .B1(net8907));
 sg13g2_a221oi_1 _32588_ (.B2(net8923),
    .C1(_09471_),
    .B1(_09467_),
    .A1(net9441),
    .Y(_09472_),
    .A2(_09463_));
 sg13g2_nand2b_1 _32589_ (.Y(_09473_),
    .B(net9432),
    .A_N(_09472_));
 sg13g2_o21ai_1 _32590_ (.B1(_09473_),
    .Y(_02688_),
    .A1(net8745),
    .A2(_09456_));
 sg13g2_a21oi_1 _32591_ (.A1(net9136),
    .A2(_10722_),
    .Y(_09474_),
    .B1(net9169));
 sg13g2_o21ai_1 _32592_ (.B1(_09474_),
    .Y(_09475_),
    .A1(net9136),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][8] ));
 sg13g2_a221oi_1 _32593_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][8] ),
    .C1(net9464),
    .B1(net8882),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][8] ),
    .Y(_09476_),
    .A2(net8773));
 sg13g2_o21ai_1 _32594_ (.B1(net9495),
    .Y(_09477_),
    .A1(net9529),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][8] ));
 sg13g2_a21oi_1 _32595_ (.A1(net9529),
    .A2(_10724_),
    .Y(_09478_),
    .B1(_09477_));
 sg13g2_a221oi_1 _32596_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][8] ),
    .C1(_09478_),
    .B1(net8883),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][8] ),
    .Y(_09479_),
    .A2(net8774));
 sg13g2_a22oi_1 _32597_ (.Y(_09480_),
    .B1(_09479_),
    .B2(net9464),
    .A2(_09476_),
    .A1(_09475_));
 sg13g2_nor2_1 _32598_ (.A(net9525),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][8] ),
    .Y(_09481_));
 sg13g2_o21ai_1 _32599_ (.B1(net9490),
    .Y(_09482_),
    .A1(net9135),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][8] ));
 sg13g2_a22oi_1 _32600_ (.Y(_09483_),
    .B1(net8880),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][8] ),
    .A2(net8771),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][8] ));
 sg13g2_o21ai_1 _32601_ (.B1(_09483_),
    .Y(_09484_),
    .A1(_09481_),
    .A2(_09482_));
 sg13g2_mux2_1 _32602_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][8] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][8] ),
    .S(net9528),
    .X(_09485_));
 sg13g2_nand2_1 _32603_ (.Y(_09486_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][8] ),
    .B(net8882));
 sg13g2_a22oi_1 _32604_ (.Y(_09487_),
    .B1(_09485_),
    .B2(net9492),
    .A2(net8773),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][8] ));
 sg13g2_a21oi_1 _32605_ (.A1(_09486_),
    .A2(_09487_),
    .Y(_09488_),
    .B1(net8912));
 sg13g2_a221oi_1 _32606_ (.B2(net8928),
    .C1(_09488_),
    .B1(_09484_),
    .A1(net9445),
    .Y(_09489_),
    .A2(_09480_));
 sg13g2_a21oi_1 _32607_ (.A1(net9136),
    .A2(_10725_),
    .Y(_09490_),
    .B1(net9169));
 sg13g2_o21ai_1 _32608_ (.B1(_09490_),
    .Y(_09491_),
    .A1(net9136),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][8] ));
 sg13g2_a221oi_1 _32609_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][8] ),
    .C1(net9464),
    .B1(net8883),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][8] ),
    .Y(_09492_),
    .A2(net8773));
 sg13g2_o21ai_1 _32610_ (.B1(net9495),
    .Y(_09493_),
    .A1(net9529),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][8] ));
 sg13g2_a21oi_1 _32611_ (.A1(net9529),
    .A2(_10727_),
    .Y(_09494_),
    .B1(_09493_));
 sg13g2_a221oi_1 _32612_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][8] ),
    .C1(_09494_),
    .B1(net8883),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][8] ),
    .Y(_09495_),
    .A2(net8774));
 sg13g2_a22oi_1 _32613_ (.Y(_09496_),
    .B1(_09495_),
    .B2(net9464),
    .A2(_09492_),
    .A1(_09491_));
 sg13g2_nor2_1 _32614_ (.A(net9528),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][8] ),
    .Y(_09497_));
 sg13g2_o21ai_1 _32615_ (.B1(net9492),
    .Y(_09498_),
    .A1(net9136),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][8] ));
 sg13g2_a22oi_1 _32616_ (.Y(_09499_),
    .B1(net8882),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][8] ),
    .A2(net8773),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][8] ));
 sg13g2_o21ai_1 _32617_ (.B1(_09499_),
    .Y(_09500_),
    .A1(_09497_),
    .A2(_09498_));
 sg13g2_mux2_1 _32618_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][8] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][8] ),
    .S(net9528),
    .X(_09501_));
 sg13g2_nand2_1 _32619_ (.Y(_09502_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][8] ),
    .B(net8883));
 sg13g2_a22oi_1 _32620_ (.Y(_09503_),
    .B1(_09501_),
    .B2(net9492),
    .A2(net8774),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][8] ));
 sg13g2_a21oi_1 _32621_ (.A1(_09502_),
    .A2(_09503_),
    .Y(_09504_),
    .B1(net8911));
 sg13g2_a221oi_1 _32622_ (.B2(net8925),
    .C1(_09504_),
    .B1(_09500_),
    .A1(net9445),
    .Y(_09505_),
    .A2(_09496_));
 sg13g2_nand2b_1 _32623_ (.Y(_09506_),
    .B(net9439),
    .A_N(_09505_));
 sg13g2_o21ai_1 _32624_ (.B1(_09506_),
    .Y(_02689_),
    .A1(net8746),
    .A2(_09489_));
 sg13g2_nor2_1 _32625_ (.A(net9537),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][9] ),
    .Y(_09507_));
 sg13g2_o21ai_1 _32626_ (.B1(net9501),
    .Y(_09508_),
    .A1(net9147),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][9] ));
 sg13g2_a221oi_1 _32627_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][9] ),
    .C1(net9470),
    .B1(net8895),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][9] ),
    .Y(_09509_),
    .A2(net8785));
 sg13g2_o21ai_1 _32628_ (.B1(_09509_),
    .Y(_09510_),
    .A1(_09507_),
    .A2(_09508_));
 sg13g2_a21oi_1 _32629_ (.A1(net9144),
    .A2(_10731_),
    .Y(_09511_),
    .B1(net9164));
 sg13g2_o21ai_1 _32630_ (.B1(_09511_),
    .Y(_09512_),
    .A1(net9144),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][9] ));
 sg13g2_a22oi_1 _32631_ (.Y(_09513_),
    .B1(net8890),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][9] ),
    .A2(net8781),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][9] ));
 sg13g2_nand3_1 _32632_ (.B(_09512_),
    .C(_09513_),
    .A(net9470),
    .Y(_09514_));
 sg13g2_nand3_1 _32633_ (.B(_09510_),
    .C(_09514_),
    .A(net9446),
    .Y(_09515_));
 sg13g2_o21ai_1 _32634_ (.B1(net9502),
    .Y(_09516_),
    .A1(net9539),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][9] ));
 sg13g2_a21oi_1 _32635_ (.A1(net9539),
    .A2(_10729_),
    .Y(_09517_),
    .B1(_09516_));
 sg13g2_a221oi_1 _32636_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][9] ),
    .C1(_09517_),
    .B1(net8897),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][9] ),
    .Y(_09518_),
    .A2(net8787));
 sg13g2_nor2_1 _32637_ (.A(net9539),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][9] ),
    .Y(_09519_));
 sg13g2_o21ai_1 _32638_ (.B1(net9502),
    .Y(_09520_),
    .A1(net9148),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][9] ));
 sg13g2_a22oi_1 _32639_ (.Y(_09521_),
    .B1(net8895),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][9] ),
    .A2(net8785),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][9] ));
 sg13g2_o21ai_1 _32640_ (.B1(_09521_),
    .Y(_09522_),
    .A1(_09519_),
    .A2(_09520_));
 sg13g2_o21ai_1 _32641_ (.B1(net9438),
    .Y(_09523_),
    .A1(net8913),
    .A2(_09518_));
 sg13g2_a21oi_1 _32642_ (.A1(net8926),
    .A2(_09522_),
    .Y(_09524_),
    .B1(_09523_));
 sg13g2_nor2_1 _32643_ (.A(net9537),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][9] ),
    .Y(_09525_));
 sg13g2_o21ai_1 _32644_ (.B1(net9501),
    .Y(_09526_),
    .A1(net9147),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][9] ));
 sg13g2_a221oi_1 _32645_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][9] ),
    .C1(net9471),
    .B1(net8895),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][9] ),
    .Y(_09527_),
    .A2(net8785));
 sg13g2_o21ai_1 _32646_ (.B1(_09527_),
    .Y(_09528_),
    .A1(_09525_),
    .A2(_09526_));
 sg13g2_a21oi_1 _32647_ (.A1(net9147),
    .A2(_10728_),
    .Y(_09529_),
    .B1(net9167));
 sg13g2_o21ai_1 _32648_ (.B1(_09529_),
    .Y(_09530_),
    .A1(net9147),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][9] ));
 sg13g2_a22oi_1 _32649_ (.Y(_09531_),
    .B1(net8896),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][9] ),
    .A2(net8786),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][9] ));
 sg13g2_nand3_1 _32650_ (.B(_09530_),
    .C(_09531_),
    .A(net9471),
    .Y(_09532_));
 sg13g2_nand3_1 _32651_ (.B(_09528_),
    .C(_09532_),
    .A(net9446),
    .Y(_09533_));
 sg13g2_mux2_1 _32652_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][9] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][9] ),
    .S(net9539),
    .X(_09534_));
 sg13g2_nand2_1 _32653_ (.Y(_09535_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][9] ),
    .B(net8895));
 sg13g2_a22oi_1 _32654_ (.Y(_09536_),
    .B1(_09534_),
    .B2(net9502),
    .A2(net8787),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][9] ));
 sg13g2_a21oi_1 _32655_ (.A1(_09535_),
    .A2(_09536_),
    .Y(_09537_),
    .B1(net8913));
 sg13g2_mux2_1 _32656_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][9] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][9] ),
    .S(net9538),
    .X(_09538_));
 sg13g2_a22oi_1 _32657_ (.Y(_09539_),
    .B1(_09538_),
    .B2(net9503),
    .A2(net8788),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][9] ));
 sg13g2_nor3_1 _32658_ (.A(net8920),
    .B(net8897),
    .C(_09539_),
    .Y(_09540_));
 sg13g2_nor3_1 _32659_ (.A(net9436),
    .B(_09537_),
    .C(_09540_),
    .Y(_09541_));
 sg13g2_a22oi_1 _32660_ (.Y(_02690_),
    .B1(_09533_),
    .B2(_09541_),
    .A2(_09524_),
    .A1(_09515_));
 sg13g2_o21ai_1 _32661_ (.B1(net9505),
    .Y(_09542_),
    .A1(net9543),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][10] ));
 sg13g2_a21oi_1 _32662_ (.A1(net9540),
    .A2(_10734_),
    .Y(_09543_),
    .B1(_09542_));
 sg13g2_a221oi_1 _32663_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][10] ),
    .C1(_09543_),
    .B1(net8901),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][10] ),
    .Y(_09544_),
    .A2(net8794));
 sg13g2_nor2_1 _32664_ (.A(net9540),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][10] ),
    .Y(_09545_));
 sg13g2_o21ai_1 _32665_ (.B1(net9505),
    .Y(_09546_),
    .A1(net9151),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][10] ));
 sg13g2_a221oi_1 _32666_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][10] ),
    .C1(net9474),
    .B1(net8900),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][10] ),
    .Y(_09547_),
    .A2(net8790));
 sg13g2_o21ai_1 _32667_ (.B1(_09547_),
    .Y(_09548_),
    .A1(_09545_),
    .A2(_09546_));
 sg13g2_nand2_1 _32668_ (.Y(_09549_),
    .A(net9447),
    .B(_09548_));
 sg13g2_a21oi_1 _32669_ (.A1(net9472),
    .A2(_09544_),
    .Y(_09550_),
    .B1(_09549_));
 sg13g2_a21oi_1 _32670_ (.A1(net9151),
    .A2(_10732_),
    .Y(_09551_),
    .B1(net9166));
 sg13g2_o21ai_1 _32671_ (.B1(_09551_),
    .Y(_09552_),
    .A1(net9151),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][10] ));
 sg13g2_a22oi_1 _32672_ (.Y(_09553_),
    .B1(net8900),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][10] ),
    .A2(net8790),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][10] ));
 sg13g2_a21oi_1 _32673_ (.A1(_09552_),
    .A2(_09553_),
    .Y(_09554_),
    .B1(net8919));
 sg13g2_a21oi_1 _32674_ (.A1(net9155),
    .A2(_10733_),
    .Y(_09555_),
    .B1(net9166));
 sg13g2_o21ai_1 _32675_ (.B1(_09555_),
    .Y(_09556_),
    .A1(net9155),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][10] ));
 sg13g2_a22oi_1 _32676_ (.Y(_09557_),
    .B1(net8900),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][10] ),
    .A2(net8790),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][10] ));
 sg13g2_a21oi_1 _32677_ (.A1(_09556_),
    .A2(_09557_),
    .Y(_09558_),
    .B1(net8914));
 sg13g2_nor4_2 _32678_ (.A(net9437),
    .B(_09550_),
    .C(_09554_),
    .Y(_09559_),
    .D(_09558_));
 sg13g2_a21oi_1 _32679_ (.A1(net9153),
    .A2(_10736_),
    .Y(_09560_),
    .B1(net9165));
 sg13g2_o21ai_1 _32680_ (.B1(_09560_),
    .Y(_09561_),
    .A1(net9153),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][10] ));
 sg13g2_a221oi_1 _32681_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][10] ),
    .C1(net9472),
    .B1(net8902),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][10] ),
    .Y(_09562_),
    .A2(net8791));
 sg13g2_mux2_1 _32682_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][10] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][10] ),
    .S(net9542),
    .X(_09563_));
 sg13g2_a22oi_1 _32683_ (.Y(_09564_),
    .B1(net8902),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][10] ),
    .A2(net8791),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][10] ));
 sg13g2_nand2_1 _32684_ (.Y(_09565_),
    .A(net9473),
    .B(_09564_));
 sg13g2_a21oi_1 _32685_ (.A1(net9505),
    .A2(_09563_),
    .Y(_09566_),
    .B1(_09565_));
 sg13g2_a21oi_1 _32686_ (.A1(_09561_),
    .A2(_09562_),
    .Y(_09567_),
    .B1(_09566_));
 sg13g2_nor2_1 _32687_ (.A(net9152),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][10] ),
    .Y(_09568_));
 sg13g2_o21ai_1 _32688_ (.B1(net9505),
    .Y(_09569_),
    .A1(net9540),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][10] ));
 sg13g2_a22oi_1 _32689_ (.Y(_09570_),
    .B1(net8902),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][10] ),
    .A2(net8791),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][10] ));
 sg13g2_o21ai_1 _32690_ (.B1(_09570_),
    .Y(_09571_),
    .A1(_09568_),
    .A2(_09569_));
 sg13g2_o21ai_1 _32691_ (.B1(net9501),
    .Y(_09572_),
    .A1(net9537),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][10] ));
 sg13g2_a21oi_1 _32692_ (.A1(net9540),
    .A2(_10735_),
    .Y(_09573_),
    .B1(_09572_));
 sg13g2_a221oi_1 _32693_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][10] ),
    .C1(_09573_),
    .B1(net8895),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][10] ),
    .Y(_09574_),
    .A2(net8785));
 sg13g2_o21ai_1 _32694_ (.B1(net9436),
    .Y(_09575_),
    .A1(net8914),
    .A2(_09574_));
 sg13g2_a221oi_1 _32695_ (.B2(net8926),
    .C1(_09575_),
    .B1(_09571_),
    .A1(net9447),
    .Y(_09576_),
    .A2(_09567_));
 sg13g2_nor3_2 _32696_ (.A(_09316_),
    .B(_09559_),
    .C(_09576_),
    .Y(_02691_));
 sg13g2_a21oi_1 _32697_ (.A1(net9116),
    .A2(_10737_),
    .Y(_09577_),
    .B1(net9158));
 sg13g2_o21ai_1 _32698_ (.B1(_09577_),
    .Y(_09578_),
    .A1(net9116),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][11] ));
 sg13g2_a221oi_1 _32699_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][11] ),
    .C1(net9451),
    .B1(net8860),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][11] ),
    .Y(_09579_),
    .A2(net8750));
 sg13g2_mux2_1 _32700_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][11] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][11] ),
    .S(net9511),
    .X(_09580_));
 sg13g2_a22oi_1 _32701_ (.Y(_09581_),
    .B1(net8862),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][11] ),
    .A2(net8751),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][11] ));
 sg13g2_nand2_1 _32702_ (.Y(_09582_),
    .A(net9451),
    .B(_09581_));
 sg13g2_a21oi_1 _32703_ (.A1(net9477),
    .A2(_09580_),
    .Y(_09583_),
    .B1(_09582_));
 sg13g2_a21oi_1 _32704_ (.A1(_09578_),
    .A2(_09579_),
    .Y(_09584_),
    .B1(_09583_));
 sg13g2_nor2_1 _32705_ (.A(net9510),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][11] ),
    .Y(_09585_));
 sg13g2_o21ai_1 _32706_ (.B1(net9476),
    .Y(_09586_),
    .A1(net9116),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][11] ));
 sg13g2_a22oi_1 _32707_ (.Y(_09587_),
    .B1(net8860),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][11] ),
    .A2(net8749),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][11] ));
 sg13g2_o21ai_1 _32708_ (.B1(_09587_),
    .Y(_09588_),
    .A1(_09585_),
    .A2(_09586_));
 sg13g2_mux2_1 _32709_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][11] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][11] ),
    .S(net9510),
    .X(_09589_));
 sg13g2_nand2_1 _32710_ (.Y(_09590_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][11] ),
    .B(net8860));
 sg13g2_a22oi_1 _32711_ (.Y(_09591_),
    .B1(_09589_),
    .B2(net9476),
    .A2(net8749),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][11] ));
 sg13g2_a21oi_1 _32712_ (.A1(_09590_),
    .A2(_09591_),
    .Y(_09592_),
    .B1(net8908));
 sg13g2_a221oi_1 _32713_ (.B2(net8922),
    .C1(_09592_),
    .B1(_09588_),
    .A1(net9440),
    .Y(_09593_),
    .A2(_09584_));
 sg13g2_a21oi_1 _32714_ (.A1(net9122),
    .A2(_10739_),
    .Y(_09594_),
    .B1(net9158));
 sg13g2_o21ai_1 _32715_ (.B1(_09594_),
    .Y(_09595_),
    .A1(net9122),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][11] ));
 sg13g2_a22oi_1 _32716_ (.Y(_09596_),
    .B1(net8867),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][11] ),
    .A2(net8756),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][11] ));
 sg13g2_nand3_1 _32717_ (.B(_09595_),
    .C(_09596_),
    .A(net9455),
    .Y(_09597_));
 sg13g2_nor2_1 _32718_ (.A(net9514),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][11] ),
    .Y(_09598_));
 sg13g2_o21ai_1 _32719_ (.B1(net9480),
    .Y(_09599_),
    .A1(net9120),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][11] ));
 sg13g2_a221oi_1 _32720_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][11] ),
    .C1(net9453),
    .B1(net8863),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][11] ),
    .Y(_09600_),
    .A2(net8753));
 sg13g2_o21ai_1 _32721_ (.B1(_09600_),
    .Y(_09601_),
    .A1(_09598_),
    .A2(_09599_));
 sg13g2_nand3_1 _32722_ (.B(_09597_),
    .C(_09601_),
    .A(net9441),
    .Y(_09602_));
 sg13g2_mux2_1 _32723_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][11] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][11] ),
    .S(net9513),
    .X(_09603_));
 sg13g2_nand2_1 _32724_ (.Y(_09604_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][11] ),
    .B(net8864));
 sg13g2_a22oi_1 _32725_ (.Y(_09605_),
    .B1(_09603_),
    .B2(net9480),
    .A2(net8753),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][11] ));
 sg13g2_a21oi_1 _32726_ (.A1(_09604_),
    .A2(_09605_),
    .Y(_09606_),
    .B1(net8917));
 sg13g2_o21ai_1 _32727_ (.B1(net9479),
    .Y(_09607_),
    .A1(net9119),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][11] ));
 sg13g2_a21oi_1 _32728_ (.A1(net9119),
    .A2(_10738_),
    .Y(_09608_),
    .B1(_09607_));
 sg13g2_a221oi_1 _32729_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][11] ),
    .C1(_09608_),
    .B1(net8863),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][11] ),
    .Y(_09609_),
    .A2(net8752));
 sg13g2_o21ai_1 _32730_ (.B1(_09602_),
    .Y(_09610_),
    .A1(net8907),
    .A2(_09609_));
 sg13g2_o21ai_1 _32731_ (.B1(net9432),
    .Y(_09611_),
    .A1(_09606_),
    .A2(_09610_));
 sg13g2_o21ai_1 _32732_ (.B1(_09611_),
    .Y(_02692_),
    .A1(net8745),
    .A2(_09593_));
 sg13g2_mux2_1 _32733_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][12] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][12] ),
    .S(net9541),
    .X(_09612_));
 sg13g2_a22oi_1 _32734_ (.Y(_09613_),
    .B1(net8900),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][12] ),
    .A2(net8790),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][12] ));
 sg13g2_nand2_1 _32735_ (.Y(_09614_),
    .A(net9474),
    .B(_09613_));
 sg13g2_a21oi_1 _32736_ (.A1(net9506),
    .A2(_09612_),
    .Y(_09615_),
    .B1(_09614_));
 sg13g2_a21oi_1 _32737_ (.A1(net9151),
    .A2(_10740_),
    .Y(_09616_),
    .B1(net9166));
 sg13g2_o21ai_1 _32738_ (.B1(_09616_),
    .Y(_09617_),
    .A1(net9151),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][12] ));
 sg13g2_a221oi_1 _32739_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][12] ),
    .C1(net9474),
    .B1(net8901),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][12] ),
    .Y(_09618_),
    .A2(net8794));
 sg13g2_a21oi_1 _32740_ (.A1(_09617_),
    .A2(_09618_),
    .Y(_09619_),
    .B1(_09615_));
 sg13g2_nor2_1 _32741_ (.A(net9541),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][12] ),
    .Y(_09620_));
 sg13g2_o21ai_1 _32742_ (.B1(net9506),
    .Y(_09621_),
    .A1(net9152),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][12] ));
 sg13g2_a22oi_1 _32743_ (.Y(_09622_),
    .B1(net8901),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][12] ),
    .A2(net8794),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][12] ));
 sg13g2_o21ai_1 _32744_ (.B1(_09622_),
    .Y(_09623_),
    .A1(_09620_),
    .A2(_09621_));
 sg13g2_mux2_1 _32745_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][12] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][12] ),
    .S(net9541),
    .X(_09624_));
 sg13g2_nand2_1 _32746_ (.Y(_09625_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][12] ),
    .B(net8901));
 sg13g2_a22oi_1 _32747_ (.Y(_09626_),
    .B1(_09624_),
    .B2(net9506),
    .A2(net8790),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][12] ));
 sg13g2_a21oi_1 _32748_ (.A1(_09625_),
    .A2(_09626_),
    .Y(_09627_),
    .B1(net8914));
 sg13g2_a221oi_1 _32749_ (.B2(net8926),
    .C1(_09627_),
    .B1(_09623_),
    .A1(net9447),
    .Y(_09628_),
    .A2(_09619_));
 sg13g2_a21oi_1 _32750_ (.A1(net9144),
    .A2(_10743_),
    .Y(_09629_),
    .B1(net9168));
 sg13g2_o21ai_1 _32751_ (.B1(_09629_),
    .Y(_09630_),
    .A1(net9144),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][12] ));
 sg13g2_a22oi_1 _32752_ (.Y(_09631_),
    .B1(net8893),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][12] ),
    .A2(net8784),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][12] ));
 sg13g2_nand3_1 _32753_ (.B(_09630_),
    .C(_09631_),
    .A(net9468),
    .Y(_09632_));
 sg13g2_nor2_1 _32754_ (.A(net9536),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][12] ),
    .Y(_09633_));
 sg13g2_o21ai_1 _32755_ (.B1(net9499),
    .Y(_09634_),
    .A1(net9143),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][12] ));
 sg13g2_a221oi_1 _32756_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][12] ),
    .C1(net9468),
    .B1(net8890),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][12] ),
    .Y(_09635_),
    .A2(net8781));
 sg13g2_o21ai_1 _32757_ (.B1(_09635_),
    .Y(_09636_),
    .A1(_09633_),
    .A2(_09634_));
 sg13g2_nand3_1 _32758_ (.B(_09632_),
    .C(_09636_),
    .A(net9449),
    .Y(_09637_));
 sg13g2_mux2_1 _32759_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][12] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][12] ),
    .S(net9536),
    .X(_09638_));
 sg13g2_nand2_1 _32760_ (.Y(_09639_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][12] ),
    .B(net8890));
 sg13g2_a22oi_1 _32761_ (.Y(_09640_),
    .B1(_09638_),
    .B2(net9499),
    .A2(net8781),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][12] ));
 sg13g2_a21oi_1 _32762_ (.A1(_09639_),
    .A2(_09640_),
    .Y(_09641_),
    .B1(net8919));
 sg13g2_o21ai_1 _32763_ (.B1(net9499),
    .Y(_09642_),
    .A1(net9144),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][12] ));
 sg13g2_a21oi_1 _32764_ (.A1(net9144),
    .A2(_10741_),
    .Y(_09643_),
    .B1(_09642_));
 sg13g2_a221oi_1 _32765_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][12] ),
    .C1(_09643_),
    .B1(net8893),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][12] ),
    .Y(_09644_),
    .A2(net8784));
 sg13g2_o21ai_1 _32766_ (.B1(_09637_),
    .Y(_09645_),
    .A1(net8915),
    .A2(_09644_));
 sg13g2_o21ai_1 _32767_ (.B1(net9438),
    .Y(_09646_),
    .A1(_09641_),
    .A2(_09645_));
 sg13g2_o21ai_1 _32768_ (.B1(_09646_),
    .Y(_02693_),
    .A1(net8746),
    .A2(_09628_));
 sg13g2_mux2_1 _32769_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][13] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][13] ),
    .S(net9544),
    .X(_09647_));
 sg13g2_a22oi_1 _32770_ (.Y(_09648_),
    .B1(net8896),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][13] ),
    .A2(net8786),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][13] ));
 sg13g2_nand2_1 _32771_ (.Y(_09649_),
    .A(net9470),
    .B(_09648_));
 sg13g2_a21oi_1 _32772_ (.A1(net9504),
    .A2(_09647_),
    .Y(_09650_),
    .B1(_09649_));
 sg13g2_a21oi_1 _32773_ (.A1(net9150),
    .A2(_10744_),
    .Y(_09651_),
    .B1(net9167));
 sg13g2_o21ai_1 _32774_ (.B1(_09651_),
    .Y(_09652_),
    .A1(net9150),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][13] ));
 sg13g2_a221oi_1 _32775_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][13] ),
    .C1(net9470),
    .B1(net8896),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][13] ),
    .Y(_09653_),
    .A2(net8786));
 sg13g2_a21oi_1 _32776_ (.A1(_09652_),
    .A2(_09653_),
    .Y(_09654_),
    .B1(_09650_));
 sg13g2_nor2_1 _32777_ (.A(net9537),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][13] ),
    .Y(_09655_));
 sg13g2_o21ai_1 _32778_ (.B1(net9501),
    .Y(_09656_),
    .A1(net9147),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][13] ));
 sg13g2_a22oi_1 _32779_ (.Y(_09657_),
    .B1(net8896),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][13] ),
    .A2(net8786),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][13] ));
 sg13g2_o21ai_1 _32780_ (.B1(_09657_),
    .Y(_09658_),
    .A1(_09655_),
    .A2(_09656_));
 sg13g2_mux2_1 _32781_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][13] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][13] ),
    .S(net9537),
    .X(_09659_));
 sg13g2_nand2_1 _32782_ (.Y(_09660_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][13] ),
    .B(net8896));
 sg13g2_a22oi_1 _32783_ (.Y(_09661_),
    .B1(_09659_),
    .B2(net9501),
    .A2(net8786),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][13] ));
 sg13g2_a21oi_1 _32784_ (.A1(_09660_),
    .A2(_09661_),
    .Y(_09662_),
    .B1(net8913));
 sg13g2_a221oi_1 _32785_ (.B2(net8926),
    .C1(_09662_),
    .B1(_09658_),
    .A1(net9446),
    .Y(_09663_),
    .A2(_09654_));
 sg13g2_a21oi_1 _32786_ (.A1(net9147),
    .A2(_10747_),
    .Y(_09664_),
    .B1(net9167));
 sg13g2_o21ai_1 _32787_ (.B1(_09664_),
    .Y(_09665_),
    .A1(net9147),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][13] ));
 sg13g2_a22oi_1 _32788_ (.Y(_09666_),
    .B1(net8895),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][13] ),
    .A2(net8785),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][13] ));
 sg13g2_nand3_1 _32789_ (.B(_09665_),
    .C(_09666_),
    .A(net9470),
    .Y(_09667_));
 sg13g2_nor2_1 _32790_ (.A(net9537),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][13] ),
    .Y(_09668_));
 sg13g2_o21ai_1 _32791_ (.B1(net9501),
    .Y(_09669_),
    .A1(net9147),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][13] ));
 sg13g2_a221oi_1 _32792_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][13] ),
    .C1(net9470),
    .B1(net8890),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][13] ),
    .Y(_09670_),
    .A2(net8781));
 sg13g2_o21ai_1 _32793_ (.B1(_09670_),
    .Y(_09671_),
    .A1(_09668_),
    .A2(_09669_));
 sg13g2_nand3_1 _32794_ (.B(_09667_),
    .C(_09671_),
    .A(net9446),
    .Y(_09672_));
 sg13g2_mux2_1 _32795_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][13] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][13] ),
    .S(net9537),
    .X(_09673_));
 sg13g2_nand2_1 _32796_ (.Y(_09674_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][13] ),
    .B(net8895));
 sg13g2_a22oi_1 _32797_ (.Y(_09675_),
    .B1(_09673_),
    .B2(net9501),
    .A2(net8785),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][13] ));
 sg13g2_a21oi_1 _32798_ (.A1(_09674_),
    .A2(_09675_),
    .Y(_09676_),
    .B1(net8919));
 sg13g2_o21ai_1 _32799_ (.B1(net9501),
    .Y(_09677_),
    .A1(net9144),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][13] ));
 sg13g2_a21oi_1 _32800_ (.A1(net9143),
    .A2(_10745_),
    .Y(_09678_),
    .B1(_09677_));
 sg13g2_a221oi_1 _32801_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][13] ),
    .C1(_09678_),
    .B1(net8895),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][13] ),
    .Y(_09679_),
    .A2(net8785));
 sg13g2_o21ai_1 _32802_ (.B1(_09672_),
    .Y(_09680_),
    .A1(net8913),
    .A2(_09679_));
 sg13g2_o21ai_1 _32803_ (.B1(net9438),
    .Y(_09681_),
    .A1(_09676_),
    .A2(_09680_));
 sg13g2_o21ai_1 _32804_ (.B1(_09681_),
    .Y(_02694_),
    .A1(net8747),
    .A2(_09663_));
 sg13g2_mux2_1 _32805_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][14] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][14] ),
    .S(net9519),
    .X(_09682_));
 sg13g2_a22oi_1 _32806_ (.Y(_09683_),
    .B1(net8872),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][14] ),
    .A2(net8761),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][14] ));
 sg13g2_nand2_1 _32807_ (.Y(_09684_),
    .A(net9457),
    .B(_09683_));
 sg13g2_a21oi_1 _32808_ (.A1(net9488),
    .A2(_09682_),
    .Y(_09685_),
    .B1(_09684_));
 sg13g2_a21oi_1 _32809_ (.A1(net9127),
    .A2(_10748_),
    .Y(_09686_),
    .B1(net9160));
 sg13g2_o21ai_1 _32810_ (.B1(_09686_),
    .Y(_09687_),
    .A1(net9128),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][14] ));
 sg13g2_a221oi_1 _32811_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][14] ),
    .C1(net9457),
    .B1(net8877),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][14] ),
    .Y(_09688_),
    .A2(net8767));
 sg13g2_a21oi_1 _32812_ (.A1(_09687_),
    .A2(_09688_),
    .Y(_09689_),
    .B1(_09685_));
 sg13g2_nor2_1 _32813_ (.A(net9521),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][14] ),
    .Y(_09690_));
 sg13g2_o21ai_1 _32814_ (.B1(net9486),
    .Y(_09691_),
    .A1(net9129),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][14] ));
 sg13g2_a22oi_1 _32815_ (.Y(_09692_),
    .B1(net8874),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][14] ),
    .A2(net8763),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][14] ));
 sg13g2_o21ai_1 _32816_ (.B1(_09692_),
    .Y(_09693_),
    .A1(_09690_),
    .A2(_09691_));
 sg13g2_mux2_1 _32817_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][14] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][14] ),
    .S(net9521),
    .X(_09694_));
 sg13g2_nand2_1 _32818_ (.Y(_09695_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][14] ),
    .B(net8874));
 sg13g2_a22oi_1 _32819_ (.Y(_09696_),
    .B1(_09694_),
    .B2(net9486),
    .A2(net8763),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][14] ));
 sg13g2_a21oi_1 _32820_ (.A1(_09695_),
    .A2(_09696_),
    .Y(_09697_),
    .B1(net8910));
 sg13g2_a221oi_1 _32821_ (.B2(net8924),
    .C1(_09697_),
    .B1(_09693_),
    .A1(net9442),
    .Y(_09698_),
    .A2(_09689_));
 sg13g2_a21oi_1 _32822_ (.A1(net9127),
    .A2(_10750_),
    .Y(_09699_),
    .B1(net9160));
 sg13g2_o21ai_1 _32823_ (.B1(_09699_),
    .Y(_09700_),
    .A1(net9127),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][14] ));
 sg13g2_a221oi_1 _32824_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][14] ),
    .C1(net9457),
    .B1(net8873),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][14] ),
    .Y(_09701_),
    .A2(net8762));
 sg13g2_o21ai_1 _32825_ (.B1(net9488),
    .Y(_09702_),
    .A1(net9519),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][14] ));
 sg13g2_a21oi_1 _32826_ (.A1(net9519),
    .A2(_10752_),
    .Y(_09703_),
    .B1(_09702_));
 sg13g2_a221oi_1 _32827_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][14] ),
    .C1(_09703_),
    .B1(net8872),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][14] ),
    .Y(_09704_),
    .A2(net8761));
 sg13g2_a22oi_1 _32828_ (.Y(_09705_),
    .B1(_09704_),
    .B2(net9457),
    .A2(_09701_),
    .A1(_09700_));
 sg13g2_nor2_1 _32829_ (.A(net9520),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][14] ),
    .Y(_09706_));
 sg13g2_o21ai_1 _32830_ (.B1(net9485),
    .Y(_09707_),
    .A1(net9127),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][14] ));
 sg13g2_a22oi_1 _32831_ (.Y(_09708_),
    .B1(net8872),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][14] ),
    .A2(net8761),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][14] ));
 sg13g2_o21ai_1 _32832_ (.B1(_09708_),
    .Y(_09709_),
    .A1(_09706_),
    .A2(_09707_));
 sg13g2_mux2_1 _32833_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][14] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][14] ),
    .S(net9520),
    .X(_09710_));
 sg13g2_nand2_1 _32834_ (.Y(_09711_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][14] ),
    .B(net8872));
 sg13g2_a22oi_1 _32835_ (.Y(_09712_),
    .B1(_09710_),
    .B2(net9485),
    .A2(net8761),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][14] ));
 sg13g2_a21oi_1 _32836_ (.A1(_09711_),
    .A2(_09712_),
    .Y(_09713_),
    .B1(net8909));
 sg13g2_a221oi_1 _32837_ (.B2(net8924),
    .C1(_09713_),
    .B1(_09709_),
    .A1(net9442),
    .Y(_09714_),
    .A2(_09705_));
 sg13g2_nand2b_1 _32838_ (.Y(_09715_),
    .B(net9435),
    .A_N(_09714_));
 sg13g2_o21ai_1 _32839_ (.B1(_09715_),
    .Y(_02695_),
    .A1(net8748),
    .A2(_09698_));
 sg13g2_nor2_1 _32840_ (.A(net9514),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][15] ),
    .Y(_09716_));
 sg13g2_o21ai_1 _32841_ (.B1(net9480),
    .Y(_09717_),
    .A1(net9121),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][15] ));
 sg13g2_a221oi_1 _32842_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][15] ),
    .C1(net9453),
    .B1(net8865),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][15] ),
    .Y(_09718_),
    .A2(net8754));
 sg13g2_o21ai_1 _32843_ (.B1(_09718_),
    .Y(_09719_),
    .A1(_09716_),
    .A2(_09717_));
 sg13g2_a21oi_1 _32844_ (.A1(net9124),
    .A2(_10755_),
    .Y(_09720_),
    .B1(net9159));
 sg13g2_o21ai_1 _32845_ (.B1(_09720_),
    .Y(_09721_),
    .A1(net9124),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][15] ));
 sg13g2_a22oi_1 _32846_ (.Y(_09722_),
    .B1(net8867),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][15] ),
    .A2(net8757),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][15] ));
 sg13g2_nand3_1 _32847_ (.B(_09721_),
    .C(_09722_),
    .A(net9455),
    .Y(_09723_));
 sg13g2_nand3_1 _32848_ (.B(_09719_),
    .C(_09723_),
    .A(net9443),
    .Y(_09724_));
 sg13g2_nor2_1 _32849_ (.A(net9124),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][15] ),
    .Y(_09725_));
 sg13g2_o21ai_1 _32850_ (.B1(net9482),
    .Y(_09726_),
    .A1(net9516),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][15] ));
 sg13g2_a22oi_1 _32851_ (.Y(_09727_),
    .B1(net8868),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][15] ),
    .A2(net8758),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][15] ));
 sg13g2_o21ai_1 _32852_ (.B1(_09727_),
    .Y(_09728_),
    .A1(_09725_),
    .A2(_09726_));
 sg13g2_o21ai_1 _32853_ (.B1(net9482),
    .Y(_09729_),
    .A1(net9516),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][15] ));
 sg13g2_a21oi_1 _32854_ (.A1(net9516),
    .A2(_10754_),
    .Y(_09730_),
    .B1(_09729_));
 sg13g2_a221oi_1 _32855_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][15] ),
    .C1(_09730_),
    .B1(net8868),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][15] ),
    .Y(_09731_),
    .A2(net8758));
 sg13g2_o21ai_1 _32856_ (.B1(net9432),
    .Y(_09732_),
    .A1(net8907),
    .A2(_09731_));
 sg13g2_a21oi_1 _32857_ (.A1(net8923),
    .A2(_09728_),
    .Y(_09733_),
    .B1(_09732_));
 sg13g2_nor2_1 _32858_ (.A(net9513),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][15] ),
    .Y(_09734_));
 sg13g2_o21ai_1 _32859_ (.B1(net9479),
    .Y(_09735_),
    .A1(net9120),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][15] ));
 sg13g2_a221oi_1 _32860_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][15] ),
    .C1(net9453),
    .B1(net8863),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][15] ),
    .Y(_09736_),
    .A2(net8752));
 sg13g2_o21ai_1 _32861_ (.B1(_09736_),
    .Y(_09737_),
    .A1(_09734_),
    .A2(_09735_));
 sg13g2_a21oi_1 _32862_ (.A1(net9120),
    .A2(_10753_),
    .Y(_09738_),
    .B1(net9158));
 sg13g2_o21ai_1 _32863_ (.B1(_09738_),
    .Y(_09739_),
    .A1(net9120),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][15] ));
 sg13g2_a22oi_1 _32864_ (.Y(_09740_),
    .B1(net8864),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][15] ),
    .A2(net8753),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][15] ));
 sg13g2_nand3_1 _32865_ (.B(_09739_),
    .C(_09740_),
    .A(net9453),
    .Y(_09741_));
 sg13g2_nand3_1 _32866_ (.B(_09737_),
    .C(_09741_),
    .A(net9440),
    .Y(_09742_));
 sg13g2_mux2_1 _32867_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][15] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][15] ),
    .S(net9514),
    .X(_09743_));
 sg13g2_nand2_1 _32868_ (.Y(_09744_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][15] ),
    .B(net8865));
 sg13g2_a22oi_1 _32869_ (.Y(_09745_),
    .B1(_09743_),
    .B2(net9480),
    .A2(net8752),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][15] ));
 sg13g2_a21oi_1 _32870_ (.A1(_09744_),
    .A2(_09745_),
    .Y(_09746_),
    .B1(net8908));
 sg13g2_mux2_1 _32871_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][15] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][15] ),
    .S(net9513),
    .X(_09747_));
 sg13g2_a22oi_1 _32872_ (.Y(_09748_),
    .B1(_09747_),
    .B2(net9479),
    .A2(net8752),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][15] ));
 sg13g2_nor3_1 _32873_ (.A(net8917),
    .B(net8866),
    .C(_09748_),
    .Y(_09749_));
 sg13g2_nor3_2 _32874_ (.A(net9432),
    .B(_09746_),
    .C(_09749_),
    .Y(_09750_));
 sg13g2_a22oi_1 _32875_ (.Y(_02696_),
    .B1(_09742_),
    .B2(_09750_),
    .A2(_09733_),
    .A1(_09724_));
 sg13g2_mux2_1 _32876_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][16] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][16] ),
    .S(net9511),
    .X(_09751_));
 sg13g2_a22oi_1 _32877_ (.Y(_09752_),
    .B1(net8862),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][16] ),
    .A2(net8749),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][16] ));
 sg13g2_nand2_1 _32878_ (.Y(_09753_),
    .A(net9451),
    .B(_09752_));
 sg13g2_a21oi_1 _32879_ (.A1(net9477),
    .A2(_09751_),
    .Y(_09754_),
    .B1(_09753_));
 sg13g2_a21oi_1 _32880_ (.A1(net9117),
    .A2(_10756_),
    .Y(_09755_),
    .B1(net9158));
 sg13g2_o21ai_1 _32881_ (.B1(_09755_),
    .Y(_09756_),
    .A1(net9117),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][16] ));
 sg13g2_a221oi_1 _32882_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][16] ),
    .C1(net9451),
    .B1(net8860),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][16] ),
    .Y(_09757_),
    .A2(net8749));
 sg13g2_a21oi_1 _32883_ (.A1(_09756_),
    .A2(_09757_),
    .Y(_09758_),
    .B1(_09754_));
 sg13g2_nor2_1 _32884_ (.A(net9511),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][16] ),
    .Y(_09759_));
 sg13g2_o21ai_1 _32885_ (.B1(net9476),
    .Y(_09760_),
    .A1(net9117),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][16] ));
 sg13g2_a22oi_1 _32886_ (.Y(_09761_),
    .B1(net8860),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][16] ),
    .A2(net8749),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][16] ));
 sg13g2_o21ai_1 _32887_ (.B1(_09761_),
    .Y(_09762_),
    .A1(_09759_),
    .A2(_09760_));
 sg13g2_mux2_1 _32888_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][16] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][16] ),
    .S(net9510),
    .X(_09763_));
 sg13g2_nand2_1 _32889_ (.Y(_09764_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][16] ),
    .B(net8861));
 sg13g2_a22oi_1 _32890_ (.Y(_09765_),
    .B1(_09763_),
    .B2(net9476),
    .A2(net8750),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][16] ));
 sg13g2_a21oi_1 _32891_ (.A1(_09764_),
    .A2(_09765_),
    .Y(_09766_),
    .B1(net8908));
 sg13g2_a221oi_1 _32892_ (.B2(net8922),
    .C1(_09766_),
    .B1(_09762_),
    .A1(net9440),
    .Y(_09767_),
    .A2(_09758_));
 sg13g2_a21oi_1 _32893_ (.A1(net9122),
    .A2(_10759_),
    .Y(_09768_),
    .B1(net9159));
 sg13g2_o21ai_1 _32894_ (.B1(_09768_),
    .Y(_09769_),
    .A1(net9122),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][16] ));
 sg13g2_a22oi_1 _32895_ (.Y(_09770_),
    .B1(net8867),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][16] ),
    .A2(net8756),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][16] ));
 sg13g2_nand3_1 _32896_ (.B(_09769_),
    .C(_09770_),
    .A(net9455),
    .Y(_09771_));
 sg13g2_nor2_1 _32897_ (.A(net9513),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][16] ),
    .Y(_09772_));
 sg13g2_o21ai_1 _32898_ (.B1(net9479),
    .Y(_09773_),
    .A1(net9120),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][16] ));
 sg13g2_a221oi_1 _32899_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][16] ),
    .C1(net9453),
    .B1(net8863),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][16] ),
    .Y(_09774_),
    .A2(net8752));
 sg13g2_o21ai_1 _32900_ (.B1(_09774_),
    .Y(_09775_),
    .A1(_09772_),
    .A2(_09773_));
 sg13g2_nand3_1 _32901_ (.B(_09771_),
    .C(_09775_),
    .A(net9441),
    .Y(_09776_));
 sg13g2_mux2_1 _32902_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][16] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][16] ),
    .S(net9513),
    .X(_09777_));
 sg13g2_nand2_1 _32903_ (.Y(_09778_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][16] ),
    .B(net8864));
 sg13g2_a22oi_1 _32904_ (.Y(_09779_),
    .B1(_09777_),
    .B2(net9479),
    .A2(net8753),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][16] ));
 sg13g2_a21oi_1 _32905_ (.A1(_09778_),
    .A2(_09779_),
    .Y(_09780_),
    .B1(net8917));
 sg13g2_o21ai_1 _32906_ (.B1(net9477),
    .Y(_09781_),
    .A1(net9118),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][16] ));
 sg13g2_a21oi_1 _32907_ (.A1(net9118),
    .A2(_10757_),
    .Y(_09782_),
    .B1(_09781_));
 sg13g2_a221oi_1 _32908_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][16] ),
    .C1(_09782_),
    .B1(net8862),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][16] ),
    .Y(_09783_),
    .A2(net8751));
 sg13g2_o21ai_1 _32909_ (.B1(_09776_),
    .Y(_09784_),
    .A1(net8907),
    .A2(_09783_));
 sg13g2_o21ai_1 _32910_ (.B1(net9432),
    .Y(_09785_),
    .A1(_09780_),
    .A2(_09784_));
 sg13g2_o21ai_1 _32911_ (.B1(_09785_),
    .Y(_02697_),
    .A1(net8745),
    .A2(_09767_));
 sg13g2_mux2_1 _32912_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][17] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][17] ),
    .S(net9510),
    .X(_09786_));
 sg13g2_a22oi_1 _32913_ (.Y(_09787_),
    .B1(net8861),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][17] ),
    .A2(net8750),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][17] ));
 sg13g2_nand2_1 _32914_ (.Y(_09788_),
    .A(net9451),
    .B(_09787_));
 sg13g2_a21oi_1 _32915_ (.A1(net9477),
    .A2(_09786_),
    .Y(_09789_),
    .B1(_09788_));
 sg13g2_a21oi_1 _32916_ (.A1(net9116),
    .A2(_10760_),
    .Y(_09790_),
    .B1(net9158));
 sg13g2_o21ai_1 _32917_ (.B1(_09790_),
    .Y(_09791_),
    .A1(net9116),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][17] ));
 sg13g2_a221oi_1 _32918_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][17] ),
    .C1(net9451),
    .B1(net8861),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][17] ),
    .Y(_09792_),
    .A2(net8750));
 sg13g2_a21oi_1 _32919_ (.A1(_09791_),
    .A2(_09792_),
    .Y(_09793_),
    .B1(_09789_));
 sg13g2_nor2_1 _32920_ (.A(net9510),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][17] ),
    .Y(_09794_));
 sg13g2_o21ai_1 _32921_ (.B1(net9476),
    .Y(_09795_),
    .A1(net9117),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][17] ));
 sg13g2_a22oi_1 _32922_ (.Y(_09796_),
    .B1(net8861),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][17] ),
    .A2(net8750),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][17] ));
 sg13g2_o21ai_1 _32923_ (.B1(_09796_),
    .Y(_09797_),
    .A1(_09794_),
    .A2(_09795_));
 sg13g2_mux2_1 _32924_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][17] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][17] ),
    .S(net9510),
    .X(_09798_));
 sg13g2_nand2_1 _32925_ (.Y(_09799_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][17] ),
    .B(net8861));
 sg13g2_a22oi_1 _32926_ (.Y(_09800_),
    .B1(_09798_),
    .B2(net9476),
    .A2(net8750),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][17] ));
 sg13g2_a21oi_1 _32927_ (.A1(_09799_),
    .A2(_09800_),
    .Y(_09801_),
    .B1(net8908));
 sg13g2_a221oi_1 _32928_ (.B2(net8922),
    .C1(_09801_),
    .B1(_09797_),
    .A1(net9440),
    .Y(_09802_),
    .A2(_09793_));
 sg13g2_nor2_1 _32929_ (.A(net9513),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][17] ),
    .Y(_09803_));
 sg13g2_o21ai_1 _32930_ (.B1(net9479),
    .Y(_09804_),
    .A1(net9120),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][17] ));
 sg13g2_a221oi_1 _32931_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][17] ),
    .C1(net9453),
    .B1(net8863),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][17] ),
    .Y(_09805_),
    .A2(net8752));
 sg13g2_o21ai_1 _32932_ (.B1(_09805_),
    .Y(_09806_),
    .A1(_09803_),
    .A2(_09804_));
 sg13g2_a21oi_1 _32933_ (.A1(net9123),
    .A2(_10763_),
    .Y(_09807_),
    .B1(net9158));
 sg13g2_o21ai_1 _32934_ (.B1(_09807_),
    .Y(_09808_),
    .A1(net9120),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][17] ));
 sg13g2_a22oi_1 _32935_ (.Y(_09809_),
    .B1(net8867),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][17] ),
    .A2(net8756),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][17] ));
 sg13g2_nand3_1 _32936_ (.B(_09808_),
    .C(_09809_),
    .A(net9453),
    .Y(_09810_));
 sg13g2_nand3_1 _32937_ (.B(_09806_),
    .C(_09810_),
    .A(net9440),
    .Y(_09811_));
 sg13g2_mux2_1 _32938_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][17] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][17] ),
    .S(net9513),
    .X(_09812_));
 sg13g2_nand2_1 _32939_ (.Y(_09813_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][17] ),
    .B(net8864));
 sg13g2_a22oi_1 _32940_ (.Y(_09814_),
    .B1(_09812_),
    .B2(net9479),
    .A2(net8753),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][17] ));
 sg13g2_a21oi_1 _32941_ (.A1(_09813_),
    .A2(_09814_),
    .Y(_09815_),
    .B1(net8917));
 sg13g2_o21ai_1 _32942_ (.B1(net9477),
    .Y(_09816_),
    .A1(net9118),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][17] ));
 sg13g2_a21oi_1 _32943_ (.A1(net9118),
    .A2(_10762_),
    .Y(_09817_),
    .B1(_09816_));
 sg13g2_a221oi_1 _32944_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][17] ),
    .C1(_09817_),
    .B1(net8862),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][17] ),
    .Y(_09818_),
    .A2(net8751));
 sg13g2_o21ai_1 _32945_ (.B1(_09811_),
    .Y(_09819_),
    .A1(net8908),
    .A2(_09818_));
 sg13g2_o21ai_1 _32946_ (.B1(net9432),
    .Y(_09820_),
    .A1(_09815_),
    .A2(_09819_));
 sg13g2_o21ai_1 _32947_ (.B1(_09820_),
    .Y(_02698_),
    .A1(net8745),
    .A2(_09802_));
 sg13g2_mux2_1 _32948_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][18] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][18] ),
    .S(net9512),
    .X(_09821_));
 sg13g2_a22oi_1 _32949_ (.Y(_09822_),
    .B1(net8861),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][18] ),
    .A2(net8750),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][18] ));
 sg13g2_nand2_1 _32950_ (.Y(_09823_),
    .A(net9452),
    .B(_09822_));
 sg13g2_a21oi_1 _32951_ (.A1(net9478),
    .A2(_09821_),
    .Y(_09824_),
    .B1(_09823_));
 sg13g2_mux2_1 _32952_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][18] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][18] ),
    .S(net9511),
    .X(_09825_));
 sg13g2_nand2_1 _32953_ (.Y(_09826_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][18] ),
    .B(net8862));
 sg13g2_a221oi_1 _32954_ (.B2(net9477),
    .C1(net9452),
    .B1(_09825_),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][18] ),
    .Y(_09827_),
    .A2(net8751));
 sg13g2_a21oi_1 _32955_ (.A1(_09826_),
    .A2(_09827_),
    .Y(_09828_),
    .B1(_09824_));
 sg13g2_nor2_1 _32956_ (.A(net9512),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][18] ),
    .Y(_09829_));
 sg13g2_o21ai_1 _32957_ (.B1(net9478),
    .Y(_09830_),
    .A1(net9119),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][18] ));
 sg13g2_a22oi_1 _32958_ (.Y(_09831_),
    .B1(net8871),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][18] ),
    .A2(net8755),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][18] ));
 sg13g2_o21ai_1 _32959_ (.B1(_09831_),
    .Y(_09832_),
    .A1(_09829_),
    .A2(_09830_));
 sg13g2_mux2_1 _32960_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][18] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][18] ),
    .S(net9512),
    .X(_09833_));
 sg13g2_nand2_1 _32961_ (.Y(_09834_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][18] ),
    .B(net8861));
 sg13g2_a22oi_1 _32962_ (.Y(_09835_),
    .B1(_09833_),
    .B2(net9478),
    .A2(net8755),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][18] ));
 sg13g2_a21oi_1 _32963_ (.A1(_09834_),
    .A2(_09835_),
    .Y(_09836_),
    .B1(net8908));
 sg13g2_a221oi_1 _32964_ (.B2(net8922),
    .C1(_09836_),
    .B1(_09832_),
    .A1(net9440),
    .Y(_09837_),
    .A2(_09828_));
 sg13g2_a21oi_1 _32965_ (.A1(net9123),
    .A2(_10764_),
    .Y(_09838_),
    .B1(net9159));
 sg13g2_o21ai_1 _32966_ (.B1(_09838_),
    .Y(_09839_),
    .A1(net9123),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][18] ));
 sg13g2_a221oi_1 _32967_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][18] ),
    .C1(net9455),
    .B1(net8866),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][18] ),
    .Y(_09840_),
    .A2(net8756));
 sg13g2_o21ai_1 _32968_ (.B1(net9483),
    .Y(_09841_),
    .A1(net9517),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][18] ));
 sg13g2_a21oi_1 _32969_ (.A1(net9517),
    .A2(_10765_),
    .Y(_09842_),
    .B1(_09841_));
 sg13g2_a221oi_1 _32970_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][18] ),
    .C1(_09842_),
    .B1(net8869),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][18] ),
    .Y(_09843_),
    .A2(net8759));
 sg13g2_a22oi_1 _32971_ (.Y(_09844_),
    .B1(_09843_),
    .B2(net9455),
    .A2(_09840_),
    .A1(_09839_));
 sg13g2_nor2_1 _32972_ (.A(net9517),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][18] ),
    .Y(_09845_));
 sg13g2_o21ai_1 _32973_ (.B1(net9484),
    .Y(_09846_),
    .A1(net9125),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][18] ));
 sg13g2_a22oi_1 _32974_ (.Y(_09847_),
    .B1(net8870),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][18] ),
    .A2(net8760),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][18] ));
 sg13g2_o21ai_1 _32975_ (.B1(_09847_),
    .Y(_09848_),
    .A1(_09845_),
    .A2(_09846_));
 sg13g2_mux2_1 _32976_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][18] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][18] ),
    .S(net9515),
    .X(_09849_));
 sg13g2_nand2_1 _32977_ (.Y(_09850_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][18] ),
    .B(net8866));
 sg13g2_a22oi_1 _32978_ (.Y(_09851_),
    .B1(_09849_),
    .B2(net9481),
    .A2(net8757),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][18] ));
 sg13g2_a21oi_1 _32979_ (.A1(_09850_),
    .A2(_09851_),
    .Y(_09852_),
    .B1(net8907));
 sg13g2_a221oi_1 _32980_ (.B2(net8923),
    .C1(_09852_),
    .B1(_09848_),
    .A1(net9441),
    .Y(_09853_),
    .A2(_09844_));
 sg13g2_nand2b_1 _32981_ (.Y(_09854_),
    .B(net9433),
    .A_N(_09853_));
 sg13g2_o21ai_1 _32982_ (.B1(_09854_),
    .Y(_02699_),
    .A1(net8745),
    .A2(_09837_));
 sg13g2_a21oi_1 _32983_ (.A1(net9127),
    .A2(_10767_),
    .Y(_09855_),
    .B1(net9160));
 sg13g2_o21ai_1 _32984_ (.B1(_09855_),
    .Y(_09856_),
    .A1(net9127),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][19] ));
 sg13g2_a221oi_1 _32985_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][19] ),
    .C1(net9457),
    .B1(net8872),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][19] ),
    .Y(_09857_),
    .A2(net8761));
 sg13g2_mux2_1 _32986_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][19] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][19] ),
    .S(net9520),
    .X(_09858_));
 sg13g2_a22oi_1 _32987_ (.Y(_09859_),
    .B1(net8872),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][19] ),
    .A2(net8761),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][19] ));
 sg13g2_nand2_1 _32988_ (.Y(_09860_),
    .A(net9457),
    .B(_09859_));
 sg13g2_a21oi_1 _32989_ (.A1(net9485),
    .A2(_09858_),
    .Y(_09861_),
    .B1(_09860_));
 sg13g2_a21oi_1 _32990_ (.A1(_09856_),
    .A2(_09857_),
    .Y(_09862_),
    .B1(_09861_));
 sg13g2_nor2_1 _32991_ (.A(net9517),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][19] ),
    .Y(_09863_));
 sg13g2_o21ai_1 _32992_ (.B1(net9483),
    .Y(_09864_),
    .A1(net9125),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][19] ));
 sg13g2_a22oi_1 _32993_ (.Y(_09865_),
    .B1(net8869),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][19] ),
    .A2(net8759),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][19] ));
 sg13g2_o21ai_1 _32994_ (.B1(_09865_),
    .Y(_09866_),
    .A1(_09863_),
    .A2(_09864_));
 sg13g2_mux2_1 _32995_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][19] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][19] ),
    .S(net9520),
    .X(_09867_));
 sg13g2_nand2_1 _32996_ (.Y(_09868_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][19] ),
    .B(net8872));
 sg13g2_a22oi_1 _32997_ (.Y(_09869_),
    .B1(_09867_),
    .B2(net9485),
    .A2(net8761),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][19] ));
 sg13g2_a21oi_1 _32998_ (.A1(_09868_),
    .A2(_09869_),
    .Y(_09870_),
    .B1(net8910));
 sg13g2_a221oi_1 _32999_ (.B2(net8922),
    .C1(_09870_),
    .B1(_09866_),
    .A1(net9441),
    .Y(_09871_),
    .A2(_09862_));
 sg13g2_a21oi_1 _33000_ (.A1(net9127),
    .A2(_10770_),
    .Y(_09872_),
    .B1(net9159));
 sg13g2_o21ai_1 _33001_ (.B1(_09872_),
    .Y(_09873_),
    .A1(net9127),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][19] ));
 sg13g2_a22oi_1 _33002_ (.Y(_09874_),
    .B1(net8872),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][19] ),
    .A2(net8761),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][19] ));
 sg13g2_nand3_1 _33003_ (.B(_09873_),
    .C(_09874_),
    .A(net9457),
    .Y(_09875_));
 sg13g2_nor2_1 _33004_ (.A(net9517),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][19] ),
    .Y(_09876_));
 sg13g2_o21ai_1 _33005_ (.B1(net9483),
    .Y(_09877_),
    .A1(net9126),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][19] ));
 sg13g2_a221oi_1 _33006_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][19] ),
    .C1(net9456),
    .B1(net8869),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][19] ),
    .Y(_09878_),
    .A2(net8759));
 sg13g2_o21ai_1 _33007_ (.B1(_09878_),
    .Y(_09879_),
    .A1(_09876_),
    .A2(_09877_));
 sg13g2_nand3_1 _33008_ (.B(_09875_),
    .C(_09879_),
    .A(net9441),
    .Y(_09880_));
 sg13g2_mux2_1 _33009_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][19] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][19] ),
    .S(net9517),
    .X(_09881_));
 sg13g2_nand2_1 _33010_ (.Y(_09882_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][19] ),
    .B(net8869));
 sg13g2_a22oi_1 _33011_ (.Y(_09883_),
    .B1(_09881_),
    .B2(net9483),
    .A2(net8759),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][19] ));
 sg13g2_a21oi_1 _33012_ (.A1(_09882_),
    .A2(_09883_),
    .Y(_09884_),
    .B1(net8917));
 sg13g2_o21ai_1 _33013_ (.B1(net9483),
    .Y(_09885_),
    .A1(net9125),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][19] ));
 sg13g2_a21oi_1 _33014_ (.A1(net9125),
    .A2(_10768_),
    .Y(_09886_),
    .B1(_09885_));
 sg13g2_a221oi_1 _33015_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][19] ),
    .C1(_09886_),
    .B1(net8869),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][19] ),
    .Y(_09887_),
    .A2(net8759));
 sg13g2_o21ai_1 _33016_ (.B1(_09880_),
    .Y(_09888_),
    .A1(net8910),
    .A2(_09887_));
 sg13g2_o21ai_1 _33017_ (.B1(net9433),
    .Y(_09889_),
    .A1(_09884_),
    .A2(_09888_));
 sg13g2_o21ai_1 _33018_ (.B1(_09889_),
    .Y(_02700_),
    .A1(net8745),
    .A2(_09871_));
 sg13g2_mux2_1 _33019_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][20] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][20] ),
    .S(net9533),
    .X(_09890_));
 sg13g2_a22oi_1 _33020_ (.Y(_09891_),
    .B1(net8889),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][20] ),
    .A2(net8780),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][20] ));
 sg13g2_nand2_1 _33021_ (.Y(_09892_),
    .A(net9467),
    .B(_09891_));
 sg13g2_a21oi_1 _33022_ (.A1(net9497),
    .A2(_09890_),
    .Y(_09893_),
    .B1(_09892_));
 sg13g2_mux2_1 _33023_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][20] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][20] ),
    .S(net9532),
    .X(_09894_));
 sg13g2_nand2_1 _33024_ (.Y(_09895_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][20] ),
    .B(net8889));
 sg13g2_a221oi_1 _33025_ (.B2(net9496),
    .C1(net9467),
    .B1(_09894_),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][20] ),
    .Y(_09896_),
    .A2(net8779));
 sg13g2_a21oi_2 _33026_ (.B1(_09893_),
    .Y(_09897_),
    .A2(_09896_),
    .A1(_09895_));
 sg13g2_nor2_1 _33027_ (.A(net9530),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][20] ),
    .Y(_09898_));
 sg13g2_o21ai_1 _33028_ (.B1(net9493),
    .Y(_09899_),
    .A1(net9138),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][20] ));
 sg13g2_a22oi_1 _33029_ (.Y(_09900_),
    .B1(net8884),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][20] ),
    .A2(net8775),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][20] ));
 sg13g2_o21ai_1 _33030_ (.B1(_09900_),
    .Y(_09901_),
    .A1(_09898_),
    .A2(_09899_));
 sg13g2_mux2_1 _33031_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][20] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][20] ),
    .S(net9530),
    .X(_09902_));
 sg13g2_nand2_1 _33032_ (.Y(_09903_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][20] ),
    .B(net8884));
 sg13g2_a22oi_1 _33033_ (.Y(_09904_),
    .B1(_09902_),
    .B2(net9493),
    .A2(net8775),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][20] ));
 sg13g2_a21oi_1 _33034_ (.A1(_09903_),
    .A2(_09904_),
    .Y(_09905_),
    .B1(net8912));
 sg13g2_a221oi_1 _33035_ (.B2(net8925),
    .C1(_09905_),
    .B1(_09901_),
    .A1(net9445),
    .Y(_09906_),
    .A2(_09897_));
 sg13g2_a21oi_1 _33036_ (.A1(net9141),
    .A2(_10774_),
    .Y(_09907_),
    .B1(net9164));
 sg13g2_o21ai_1 _33037_ (.B1(_09907_),
    .Y(_09908_),
    .A1(net9141),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][20] ));
 sg13g2_a22oi_1 _33038_ (.Y(_09909_),
    .B1(net8889),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][20] ),
    .A2(net8779),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][20] ));
 sg13g2_nand3_1 _33039_ (.B(_09908_),
    .C(_09909_),
    .A(net9467),
    .Y(_09910_));
 sg13g2_nor2_1 _33040_ (.A(net9532),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][20] ),
    .Y(_09911_));
 sg13g2_o21ai_1 _33041_ (.B1(net9496),
    .Y(_09912_),
    .A1(net9141),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][20] ));
 sg13g2_a221oi_1 _33042_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][20] ),
    .C1(net9467),
    .B1(net8889),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][20] ),
    .Y(_09913_),
    .A2(net8779));
 sg13g2_o21ai_1 _33043_ (.B1(_09913_),
    .Y(_09914_),
    .A1(_09911_),
    .A2(_09912_));
 sg13g2_nand3_1 _33044_ (.B(_09910_),
    .C(_09914_),
    .A(net9449),
    .Y(_09915_));
 sg13g2_mux2_1 _33045_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][20] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][20] ),
    .S(net9530),
    .X(_09916_));
 sg13g2_nand2_1 _33046_ (.Y(_09917_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][20] ),
    .B(net8884));
 sg13g2_a22oi_1 _33047_ (.Y(_09918_),
    .B1(_09916_),
    .B2(net9493),
    .A2(net8775),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][20] ));
 sg13g2_a21oi_1 _33048_ (.A1(_09917_),
    .A2(_09918_),
    .Y(_09919_),
    .B1(net8921));
 sg13g2_o21ai_1 _33049_ (.B1(net9494),
    .Y(_09920_),
    .A1(net9138),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][20] ));
 sg13g2_a21oi_1 _33050_ (.A1(net9138),
    .A2(_10772_),
    .Y(_09921_),
    .B1(_09920_));
 sg13g2_a221oi_1 _33051_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][20] ),
    .C1(_09921_),
    .B1(net8885),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][20] ),
    .Y(_09922_),
    .A2(net8776));
 sg13g2_o21ai_1 _33052_ (.B1(_09915_),
    .Y(_09923_),
    .A1(net8911),
    .A2(_09922_));
 sg13g2_o21ai_1 _33053_ (.B1(net9439),
    .Y(_09924_),
    .A1(_09919_),
    .A2(_09923_));
 sg13g2_o21ai_1 _33054_ (.B1(_09924_),
    .Y(_02701_),
    .A1(net8746),
    .A2(_09906_));
 sg13g2_mux2_1 _33055_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][21] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][21] ),
    .S(net9527),
    .X(_09925_));
 sg13g2_a22oi_1 _33056_ (.Y(_09926_),
    .B1(net8878),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][21] ),
    .A2(net8769),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][21] ));
 sg13g2_nand2_1 _33057_ (.Y(_09927_),
    .A(net9462),
    .B(_09926_));
 sg13g2_a21oi_1 _33058_ (.A1(net9491),
    .A2(_09925_),
    .Y(_09928_),
    .B1(_09927_));
 sg13g2_a21oi_1 _33059_ (.A1(net9135),
    .A2(_10775_),
    .Y(_09929_),
    .B1(net9163));
 sg13g2_o21ai_1 _33060_ (.B1(_09929_),
    .Y(_09930_),
    .A1(net9135),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][21] ));
 sg13g2_a221oi_1 _33061_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][21] ),
    .C1(net9462),
    .B1(net8879),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][21] ),
    .Y(_09931_),
    .A2(net8770));
 sg13g2_a21oi_1 _33062_ (.A1(_09930_),
    .A2(_09931_),
    .Y(_09932_),
    .B1(_09928_));
 sg13g2_nor2_1 _33063_ (.A(net9527),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][21] ),
    .Y(_09933_));
 sg13g2_o21ai_1 _33064_ (.B1(net9489),
    .Y(_09934_),
    .A1(net9135),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][21] ));
 sg13g2_a22oi_1 _33065_ (.Y(_09935_),
    .B1(net8878),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][21] ),
    .A2(net8770),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][21] ));
 sg13g2_o21ai_1 _33066_ (.B1(_09935_),
    .Y(_09936_),
    .A1(_09933_),
    .A2(_09934_));
 sg13g2_mux2_1 _33067_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][21] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][21] ),
    .S(net9527),
    .X(_09937_));
 sg13g2_nand2_1 _33068_ (.Y(_09938_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][21] ),
    .B(net8878));
 sg13g2_a22oi_1 _33069_ (.Y(_09939_),
    .B1(_09937_),
    .B2(net9489),
    .A2(net8769),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][21] ));
 sg13g2_a21oi_1 _33070_ (.A1(_09938_),
    .A2(_09939_),
    .Y(_09940_),
    .B1(net8911));
 sg13g2_a221oi_1 _33071_ (.B2(net8925),
    .C1(_09940_),
    .B1(_09936_),
    .A1(net9444),
    .Y(_09941_),
    .A2(_09932_));
 sg13g2_a21oi_1 _33072_ (.A1(net9131),
    .A2(_10778_),
    .Y(_09942_),
    .B1(net9161));
 sg13g2_o21ai_1 _33073_ (.B1(_09942_),
    .Y(_09943_),
    .A1(net9131),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][21] ));
 sg13g2_a22oi_1 _33074_ (.Y(_09944_),
    .B1(net8878),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][21] ),
    .A2(net8766),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][21] ));
 sg13g2_nand3_1 _33075_ (.B(_09943_),
    .C(_09944_),
    .A(net9459),
    .Y(_09945_));
 sg13g2_nor2_1 _33076_ (.A(net9527),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][21] ),
    .Y(_09946_));
 sg13g2_o21ai_1 _33077_ (.B1(net9489),
    .Y(_09947_),
    .A1(net9131),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][21] ));
 sg13g2_a221oi_1 _33078_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][21] ),
    .C1(net9462),
    .B1(net8878),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][21] ),
    .Y(_09948_),
    .A2(net8769));
 sg13g2_o21ai_1 _33079_ (.B1(_09948_),
    .Y(_09949_),
    .A1(_09946_),
    .A2(_09947_));
 sg13g2_nand3_1 _33080_ (.B(_09945_),
    .C(_09949_),
    .A(net9444),
    .Y(_09950_));
 sg13g2_mux2_1 _33081_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][21] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][21] ),
    .S(net9527),
    .X(_09951_));
 sg13g2_nand2_1 _33082_ (.Y(_09952_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][21] ),
    .B(net8878));
 sg13g2_a22oi_1 _33083_ (.Y(_09953_),
    .B1(_09951_),
    .B2(net9489),
    .A2(net8769),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][21] ));
 sg13g2_a21oi_1 _33084_ (.A1(_09952_),
    .A2(_09953_),
    .Y(_09954_),
    .B1(net8917));
 sg13g2_o21ai_1 _33085_ (.B1(net9487),
    .Y(_09955_),
    .A1(net9131),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][21] ));
 sg13g2_a21oi_1 _33086_ (.A1(net9130),
    .A2(_10776_),
    .Y(_09956_),
    .B1(_09955_));
 sg13g2_a221oi_1 _33087_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][21] ),
    .C1(_09956_),
    .B1(net8876),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][21] ),
    .Y(_09957_),
    .A2(net8765));
 sg13g2_o21ai_1 _33088_ (.B1(_09950_),
    .Y(_09958_),
    .A1(net8909),
    .A2(_09957_));
 sg13g2_o21ai_1 _33089_ (.B1(net9435),
    .Y(_09959_),
    .A1(_09954_),
    .A2(_09958_));
 sg13g2_o21ai_1 _33090_ (.B1(_09959_),
    .Y(_02702_),
    .A1(net8746),
    .A2(_09941_));
 sg13g2_nor2_1 _33091_ (.A(net9543),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][22] ),
    .Y(_09960_));
 sg13g2_o21ai_1 _33092_ (.B1(net9508),
    .Y(_09961_),
    .A1(net9155),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][22] ));
 sg13g2_a221oi_1 _33093_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][22] ),
    .C1(net9473),
    .B1(net8903),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][22] ),
    .Y(_09962_),
    .A2(net8792));
 sg13g2_o21ai_1 _33094_ (.B1(_09962_),
    .Y(_09963_),
    .A1(_09960_),
    .A2(_09961_));
 sg13g2_a21oi_1 _33095_ (.A1(net9155),
    .A2(_10781_),
    .Y(_09964_),
    .B1(net9166));
 sg13g2_o21ai_1 _33096_ (.B1(_09964_),
    .Y(_09965_),
    .A1(net9155),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][22] ));
 sg13g2_a22oi_1 _33097_ (.Y(_09966_),
    .B1(net8903),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][22] ),
    .A2(net8792),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][22] ));
 sg13g2_nand3_1 _33098_ (.B(_09965_),
    .C(_09966_),
    .A(net9473),
    .Y(_09967_));
 sg13g2_and3_1 _33099_ (.X(_09968_),
    .A(net9447),
    .B(_09963_),
    .C(_09967_));
 sg13g2_a21oi_1 _33100_ (.A1(net9155),
    .A2(_10780_),
    .Y(_09969_),
    .B1(net9165));
 sg13g2_o21ai_1 _33101_ (.B1(_09969_),
    .Y(_09970_),
    .A1(net9155),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][22] ));
 sg13g2_a22oi_1 _33102_ (.Y(_09971_),
    .B1(net8903),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][22] ),
    .A2(net8792),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][22] ));
 sg13g2_a21oi_1 _33103_ (.A1(_09970_),
    .A2(_09971_),
    .Y(_09972_),
    .B1(net8914));
 sg13g2_a21oi_1 _33104_ (.A1(net9156),
    .A2(_10779_),
    .Y(_09973_),
    .B1(net9165));
 sg13g2_o21ai_1 _33105_ (.B1(_09973_),
    .Y(_09974_),
    .A1(net9155),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][22] ));
 sg13g2_a22oi_1 _33106_ (.Y(_09975_),
    .B1(net8903),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][22] ),
    .A2(net8792),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][22] ));
 sg13g2_a21oi_1 _33107_ (.A1(_09974_),
    .A2(_09975_),
    .Y(_09976_),
    .B1(net8919));
 sg13g2_nor4_2 _33108_ (.A(net9436),
    .B(_09968_),
    .C(_09972_),
    .Y(_09977_),
    .D(_09976_));
 sg13g2_mux2_1 _33109_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][22] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][22] ),
    .S(net9542),
    .X(_09978_));
 sg13g2_a22oi_1 _33110_ (.Y(_09979_),
    .B1(net8904),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][22] ),
    .A2(net8793),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][22] ));
 sg13g2_nand2_1 _33111_ (.Y(_09980_),
    .A(net9472),
    .B(_09979_));
 sg13g2_a21oi_1 _33112_ (.A1(net9507),
    .A2(_09978_),
    .Y(_09981_),
    .B1(_09980_));
 sg13g2_a21oi_1 _33113_ (.A1(net9153),
    .A2(_10783_),
    .Y(_09982_),
    .B1(net9167));
 sg13g2_o21ai_1 _33114_ (.B1(_09982_),
    .Y(_09983_),
    .A1(net9149),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][22] ));
 sg13g2_a221oi_1 _33115_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][22] ),
    .C1(net9472),
    .B1(net8897),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][22] ),
    .Y(_09984_),
    .A2(net8787));
 sg13g2_a21oi_1 _33116_ (.A1(_09983_),
    .A2(_09984_),
    .Y(_09985_),
    .B1(_09981_));
 sg13g2_o21ai_1 _33117_ (.B1(net9502),
    .Y(_09986_),
    .A1(net9539),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][22] ));
 sg13g2_a21oi_1 _33118_ (.A1(net9538),
    .A2(_10782_),
    .Y(_09987_),
    .B1(_09986_));
 sg13g2_a221oi_1 _33119_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][22] ),
    .C1(_09987_),
    .B1(net8897),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][22] ),
    .Y(_09988_),
    .A2(net8787));
 sg13g2_nor2_1 _33120_ (.A(net9149),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][22] ),
    .Y(_09989_));
 sg13g2_o21ai_1 _33121_ (.B1(net9502),
    .Y(_09990_),
    .A1(net9538),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][22] ));
 sg13g2_a22oi_1 _33122_ (.Y(_09991_),
    .B1(net8898),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][22] ),
    .A2(net8788),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][22] ));
 sg13g2_o21ai_1 _33123_ (.B1(_09991_),
    .Y(_09992_),
    .A1(_09989_),
    .A2(_09990_));
 sg13g2_o21ai_1 _33124_ (.B1(net9436),
    .Y(_09993_),
    .A1(net8913),
    .A2(_09988_));
 sg13g2_a221oi_1 _33125_ (.B2(net8926),
    .C1(_09993_),
    .B1(_09992_),
    .A1(net9447),
    .Y(_09994_),
    .A2(_09985_));
 sg13g2_nor3_2 _33126_ (.A(_09316_),
    .B(_09977_),
    .C(_09994_),
    .Y(_02703_));
 sg13g2_mux2_1 _33127_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][23] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][23] ),
    .S(net9514),
    .X(_09995_));
 sg13g2_a22oi_1 _33128_ (.Y(_09996_),
    .B1(net8865),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][23] ),
    .A2(net8754),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][23] ));
 sg13g2_nand2_1 _33129_ (.Y(_09997_),
    .A(net9454),
    .B(_09996_));
 sg13g2_a21oi_1 _33130_ (.A1(net9480),
    .A2(_09995_),
    .Y(_09998_),
    .B1(_09997_));
 sg13g2_a21oi_1 _33131_ (.A1(net9118),
    .A2(_10784_),
    .Y(_09999_),
    .B1(net9158));
 sg13g2_o21ai_1 _33132_ (.B1(_09999_),
    .Y(_10000_),
    .A1(net9118),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][23] ));
 sg13g2_a221oi_1 _33133_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][23] ),
    .C1(net9451),
    .B1(net8863),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][23] ),
    .Y(_10001_),
    .A2(net8752));
 sg13g2_a21oi_1 _33134_ (.A1(_10000_),
    .A2(_10001_),
    .Y(_10002_),
    .B1(_09998_));
 sg13g2_nor2_1 _33135_ (.A(net9513),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][23] ),
    .Y(_10003_));
 sg13g2_o21ai_1 _33136_ (.B1(net9479),
    .Y(_10004_),
    .A1(net9120),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][23] ));
 sg13g2_a22oi_1 _33137_ (.Y(_10005_),
    .B1(net8863),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][23] ),
    .A2(net8752),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][23] ));
 sg13g2_o21ai_1 _33138_ (.B1(_10005_),
    .Y(_10006_),
    .A1(_10003_),
    .A2(_10004_));
 sg13g2_mux2_1 _33139_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][23] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][23] ),
    .S(net9514),
    .X(_10007_));
 sg13g2_nand2_1 _33140_ (.Y(_10008_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][23] ),
    .B(net8863));
 sg13g2_a22oi_1 _33141_ (.Y(_10009_),
    .B1(_10007_),
    .B2(net9480),
    .A2(net8754),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][23] ));
 sg13g2_a21oi_1 _33142_ (.A1(_10008_),
    .A2(_10009_),
    .Y(_10010_),
    .B1(net8908));
 sg13g2_a221oi_1 _33143_ (.B2(net8922),
    .C1(_10010_),
    .B1(_10006_),
    .A1(net9441),
    .Y(_10011_),
    .A2(_10002_));
 sg13g2_nor2_1 _33144_ (.A(net9514),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][23] ),
    .Y(_10012_));
 sg13g2_o21ai_1 _33145_ (.B1(net9480),
    .Y(_10013_),
    .A1(net9121),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][23] ));
 sg13g2_a221oi_1 _33146_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][23] ),
    .C1(net9454),
    .B1(net8865),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][23] ),
    .Y(_10014_),
    .A2(net8754));
 sg13g2_o21ai_1 _33147_ (.B1(_10014_),
    .Y(_10015_),
    .A1(_10012_),
    .A2(_10013_));
 sg13g2_a21oi_1 _33148_ (.A1(net9124),
    .A2(_10787_),
    .Y(_10016_),
    .B1(net9159));
 sg13g2_o21ai_1 _33149_ (.B1(_10016_),
    .Y(_10017_),
    .A1(net9124),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][23] ));
 sg13g2_a22oi_1 _33150_ (.Y(_10018_),
    .B1(net8868),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][23] ),
    .A2(net8758),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][23] ));
 sg13g2_nand3_1 _33151_ (.B(_10017_),
    .C(_10018_),
    .A(net9455),
    .Y(_10019_));
 sg13g2_nand3_1 _33152_ (.B(_10015_),
    .C(_10019_),
    .A(net9440),
    .Y(_10020_));
 sg13g2_mux2_1 _33153_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][23] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][23] ),
    .S(net9516),
    .X(_10021_));
 sg13g2_nand2_1 _33154_ (.Y(_10022_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][23] ),
    .B(net8868));
 sg13g2_a22oi_1 _33155_ (.Y(_10023_),
    .B1(_10021_),
    .B2(net9482),
    .A2(net8758),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][23] ));
 sg13g2_a21oi_1 _33156_ (.A1(_10022_),
    .A2(_10023_),
    .Y(_10024_),
    .B1(net8917));
 sg13g2_o21ai_1 _33157_ (.B1(net9481),
    .Y(_10025_),
    .A1(net9122),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][23] ));
 sg13g2_a21oi_1 _33158_ (.A1(net9122),
    .A2(_10786_),
    .Y(_10026_),
    .B1(_10025_));
 sg13g2_a221oi_1 _33159_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][23] ),
    .C1(_10026_),
    .B1(net8867),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][23] ),
    .Y(_10027_),
    .A2(net8756));
 sg13g2_o21ai_1 _33160_ (.B1(_10020_),
    .Y(_10028_),
    .A1(net8907),
    .A2(_10027_));
 sg13g2_o21ai_1 _33161_ (.B1(net9433),
    .Y(_10029_),
    .A1(_10024_),
    .A2(_10028_));
 sg13g2_o21ai_1 _33162_ (.B1(_10029_),
    .Y(_02704_),
    .A1(net8745),
    .A2(_10011_));
 sg13g2_a21oi_1 _33163_ (.A1(net9134),
    .A2(_10788_),
    .Y(_10030_),
    .B1(net9163));
 sg13g2_o21ai_1 _33164_ (.B1(_10030_),
    .Y(_10031_),
    .A1(net9134),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][24] ));
 sg13g2_a221oi_1 _33165_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][24] ),
    .C1(net9462),
    .B1(net8880),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][24] ),
    .Y(_10032_),
    .A2(net8771));
 sg13g2_mux2_1 _33166_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][24] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][24] ),
    .S(net9525),
    .X(_10033_));
 sg13g2_a22oi_1 _33167_ (.Y(_10034_),
    .B1(net8880),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][24] ),
    .A2(net8771),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][24] ));
 sg13g2_nand2_1 _33168_ (.Y(_10035_),
    .A(net9463),
    .B(_10034_));
 sg13g2_a21oi_1 _33169_ (.A1(net9490),
    .A2(_10033_),
    .Y(_10036_),
    .B1(_10035_));
 sg13g2_a21oi_1 _33170_ (.A1(_10031_),
    .A2(_10032_),
    .Y(_10037_),
    .B1(_10036_));
 sg13g2_nor2_1 _33171_ (.A(net9525),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][24] ),
    .Y(_10038_));
 sg13g2_o21ai_1 _33172_ (.B1(net9490),
    .Y(_10039_),
    .A1(net9134),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][24] ));
 sg13g2_a22oi_1 _33173_ (.Y(_10040_),
    .B1(net8880),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][24] ),
    .A2(net8771),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][24] ));
 sg13g2_o21ai_1 _33174_ (.B1(_10040_),
    .Y(_10041_),
    .A1(_10038_),
    .A2(_10039_));
 sg13g2_mux2_1 _33175_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][24] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][24] ),
    .S(net9526),
    .X(_10042_));
 sg13g2_nand2_1 _33176_ (.Y(_10043_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][24] ),
    .B(net8880));
 sg13g2_a22oi_1 _33177_ (.Y(_10044_),
    .B1(_10042_),
    .B2(net9490),
    .A2(net8771),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][24] ));
 sg13g2_a21oi_1 _33178_ (.A1(_10043_),
    .A2(_10044_),
    .Y(_10045_),
    .B1(net8911));
 sg13g2_a221oi_1 _33179_ (.B2(net8925),
    .C1(_10045_),
    .B1(_10041_),
    .A1(net9444),
    .Y(_10046_),
    .A2(_10037_));
 sg13g2_a21oi_1 _33180_ (.A1(net9135),
    .A2(_10789_),
    .Y(_10047_),
    .B1(net9163));
 sg13g2_o21ai_1 _33181_ (.B1(_10047_),
    .Y(_10048_),
    .A1(net9135),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][24] ));
 sg13g2_a221oi_1 _33182_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][24] ),
    .C1(net9462),
    .B1(net8879),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][24] ),
    .Y(_10049_),
    .A2(net8770));
 sg13g2_o21ai_1 _33183_ (.B1(net9489),
    .Y(_10050_),
    .A1(net9525),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][24] ));
 sg13g2_a21oi_1 _33184_ (.A1(net9525),
    .A2(_10790_),
    .Y(_10051_),
    .B1(_10050_));
 sg13g2_a221oi_1 _33185_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][24] ),
    .C1(_10051_),
    .B1(net8879),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][24] ),
    .Y(_10052_),
    .A2(net8770));
 sg13g2_a22oi_1 _33186_ (.Y(_10053_),
    .B1(_10052_),
    .B2(net9462),
    .A2(_10049_),
    .A1(_10048_));
 sg13g2_nor2_1 _33187_ (.A(net9527),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][24] ),
    .Y(_10054_));
 sg13g2_o21ai_1 _33188_ (.B1(net9489),
    .Y(_10055_),
    .A1(net9135),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][24] ));
 sg13g2_a22oi_1 _33189_ (.Y(_10056_),
    .B1(net8878),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][24] ),
    .A2(net8769),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][24] ));
 sg13g2_o21ai_1 _33190_ (.B1(_10056_),
    .Y(_10057_),
    .A1(_10054_),
    .A2(_10055_));
 sg13g2_mux2_1 _33191_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][24] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][24] ),
    .S(net9527),
    .X(_10058_));
 sg13g2_nand2_1 _33192_ (.Y(_10059_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][24] ),
    .B(net8879));
 sg13g2_a22oi_1 _33193_ (.Y(_10060_),
    .B1(_10058_),
    .B2(net9489),
    .A2(net8769),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][24] ));
 sg13g2_a21oi_1 _33194_ (.A1(_10059_),
    .A2(_10060_),
    .Y(_10061_),
    .B1(net8911));
 sg13g2_a221oi_1 _33195_ (.B2(net8925),
    .C1(_10061_),
    .B1(_10057_),
    .A1(net9444),
    .Y(_10062_),
    .A2(_10053_));
 sg13g2_nand2b_1 _33196_ (.Y(_10063_),
    .B(net9434),
    .A_N(_10062_));
 sg13g2_o21ai_1 _33197_ (.B1(_10063_),
    .Y(_02705_),
    .A1(net8746),
    .A2(_10046_));
 sg13g2_a21oi_1 _33198_ (.A1(net9142),
    .A2(_10793_),
    .Y(_10064_),
    .B1(net9164));
 sg13g2_o21ai_1 _33199_ (.B1(_10064_),
    .Y(_10065_),
    .A1(net9142),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][25] ));
 sg13g2_a221oi_1 _33200_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][25] ),
    .C1(net9467),
    .B1(net8894),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][25] ),
    .Y(_10066_),
    .A2(net8780));
 sg13g2_mux2_1 _33201_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][25] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][25] ),
    .S(net9534),
    .X(_10067_));
 sg13g2_a22oi_1 _33202_ (.Y(_10068_),
    .B1(net8894),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][25] ),
    .A2(net8780),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][25] ));
 sg13g2_nand2_1 _33203_ (.Y(_10069_),
    .A(net9469),
    .B(_10068_));
 sg13g2_a21oi_1 _33204_ (.A1(net9497),
    .A2(_10067_),
    .Y(_10070_),
    .B1(_10069_));
 sg13g2_a21oi_1 _33205_ (.A1(_10065_),
    .A2(_10066_),
    .Y(_10071_),
    .B1(_10070_));
 sg13g2_o21ai_1 _33206_ (.B1(net9496),
    .Y(_10072_),
    .A1(net9532),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][25] ));
 sg13g2_a21oi_1 _33207_ (.A1(net9532),
    .A2(_10792_),
    .Y(_10073_),
    .B1(_10072_));
 sg13g2_a221oi_1 _33208_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][25] ),
    .C1(_10073_),
    .B1(net8889),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][25] ),
    .Y(_10074_),
    .A2(net8775));
 sg13g2_nor2_1 _33209_ (.A(net9534),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][25] ),
    .Y(_10075_));
 sg13g2_o21ai_1 _33210_ (.B1(net9497),
    .Y(_10076_),
    .A1(net9139),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][25] ));
 sg13g2_a22oi_1 _33211_ (.Y(_10077_),
    .B1(net8886),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][25] ),
    .A2(net8777),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][25] ));
 sg13g2_o21ai_1 _33212_ (.B1(_10077_),
    .Y(_10078_),
    .A1(_10075_),
    .A2(_10076_));
 sg13g2_o21ai_1 _33213_ (.B1(net9439),
    .Y(_10079_),
    .A1(net8915),
    .A2(_10074_));
 sg13g2_a221oi_1 _33214_ (.B2(net8927),
    .C1(_10079_),
    .B1(_10078_),
    .A1(net9449),
    .Y(_10080_),
    .A2(_10071_));
 sg13g2_nor2_1 _33215_ (.A(net9530),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][25] ),
    .Y(_10081_));
 sg13g2_o21ai_1 _33216_ (.B1(net9494),
    .Y(_10082_),
    .A1(net9138),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][25] ));
 sg13g2_a221oi_1 _33217_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][25] ),
    .C1(net9465),
    .B1(net8884),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][25] ),
    .Y(_10083_),
    .A2(net8776));
 sg13g2_o21ai_1 _33218_ (.B1(_10083_),
    .Y(_10084_),
    .A1(_10081_),
    .A2(_10082_));
 sg13g2_a21oi_1 _33219_ (.A1(net9139),
    .A2(_10791_),
    .Y(_10085_),
    .B1(net9169));
 sg13g2_o21ai_1 _33220_ (.B1(_10085_),
    .Y(_10086_),
    .A1(net9139),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][25] ));
 sg13g2_a22oi_1 _33221_ (.Y(_10087_),
    .B1(net8886),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][25] ),
    .A2(net8777),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][25] ));
 sg13g2_nand3_1 _33222_ (.B(_10086_),
    .C(_10087_),
    .A(net9465),
    .Y(_10088_));
 sg13g2_nand3_1 _33223_ (.B(_10084_),
    .C(_10088_),
    .A(net9445),
    .Y(_10089_));
 sg13g2_mux2_1 _33224_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][25] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][25] ),
    .S(net9534),
    .X(_10090_));
 sg13g2_nand2_1 _33225_ (.Y(_10091_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][25] ),
    .B(net8888));
 sg13g2_a22oi_1 _33226_ (.Y(_10092_),
    .B1(_10090_),
    .B2(net9497),
    .A2(net8780),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][25] ));
 sg13g2_a21oi_1 _33227_ (.A1(_10091_),
    .A2(_10092_),
    .Y(_10093_),
    .B1(net8915));
 sg13g2_a21o_1 _33228_ (.A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][25] ),
    .A1(net9141),
    .B1(net9164),
    .X(_10094_));
 sg13g2_a21oi_1 _33229_ (.A1(net9532),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][25] ),
    .Y(_10095_),
    .B1(_10094_));
 sg13g2_nor2_1 _33230_ (.A(net9496),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][25] ),
    .Y(_10096_));
 sg13g2_nor4_1 _33231_ (.A(net8919),
    .B(net8888),
    .C(_10095_),
    .D(_10096_),
    .Y(_10097_));
 sg13g2_nor3_2 _33232_ (.A(net9438),
    .B(_10093_),
    .C(_10097_),
    .Y(_10098_));
 sg13g2_a21oi_2 _33233_ (.B1(_10080_),
    .Y(_02706_),
    .A2(_10098_),
    .A1(_10089_));
 sg13g2_a21oi_1 _33234_ (.A1(net9154),
    .A2(_10796_),
    .Y(_10099_),
    .B1(net9165));
 sg13g2_o21ai_1 _33235_ (.B1(_10099_),
    .Y(_10100_),
    .A1(net9154),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][26] ));
 sg13g2_a22oi_1 _33236_ (.Y(_10101_),
    .B1(net8904),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][26] ),
    .A2(net8792),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][26] ));
 sg13g2_nand3_1 _33237_ (.B(_10100_),
    .C(_10101_),
    .A(net9473),
    .Y(_10102_));
 sg13g2_nor2_1 _33238_ (.A(net9542),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][26] ),
    .Y(_10103_));
 sg13g2_o21ai_1 _33239_ (.B1(net9507),
    .Y(_10104_),
    .A1(net9154),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][26] ));
 sg13g2_a221oi_1 _33240_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][26] ),
    .C1(net9473),
    .B1(net8904),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][26] ),
    .Y(_10105_),
    .A2(net8792));
 sg13g2_o21ai_1 _33241_ (.B1(_10105_),
    .Y(_10106_),
    .A1(_10103_),
    .A2(_10104_));
 sg13g2_nand3_1 _33242_ (.B(_10102_),
    .C(_10106_),
    .A(net9447),
    .Y(_10107_));
 sg13g2_a21oi_1 _33243_ (.A1(net9156),
    .A2(_10794_),
    .Y(_10108_),
    .B1(net9165));
 sg13g2_o21ai_1 _33244_ (.B1(_10108_),
    .Y(_10109_),
    .A1(net9154),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][26] ));
 sg13g2_a22oi_1 _33245_ (.Y(_10110_),
    .B1(net8903),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][26] ),
    .A2(net8793),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][26] ));
 sg13g2_a21oi_1 _33246_ (.A1(_10109_),
    .A2(_10110_),
    .Y(_10111_),
    .B1(net8920));
 sg13g2_a21oi_1 _33247_ (.A1(net9154),
    .A2(_10795_),
    .Y(_10112_),
    .B1(net9165));
 sg13g2_o21ai_1 _33248_ (.B1(_10112_),
    .Y(_10113_),
    .A1(net9154),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][26] ));
 sg13g2_a22oi_1 _33249_ (.Y(_10114_),
    .B1(net8903),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][26] ),
    .A2(net8793),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][26] ));
 sg13g2_a21oi_1 _33250_ (.A1(_10113_),
    .A2(_10114_),
    .Y(_10115_),
    .B1(net8914));
 sg13g2_nor3_2 _33251_ (.A(net9436),
    .B(_10111_),
    .C(_10115_),
    .Y(_10116_));
 sg13g2_nor2_1 _33252_ (.A(net9542),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][26] ),
    .Y(_10117_));
 sg13g2_o21ai_1 _33253_ (.B1(net9507),
    .Y(_10118_),
    .A1(net9149),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][26] ));
 sg13g2_a221oi_1 _33254_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][26] ),
    .C1(net9472),
    .B1(net8897),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][26] ),
    .Y(_10119_),
    .A2(net8787));
 sg13g2_o21ai_1 _33255_ (.B1(_10119_),
    .Y(_10120_),
    .A1(_10117_),
    .A2(_10118_));
 sg13g2_a21oi_1 _33256_ (.A1(net9153),
    .A2(_10798_),
    .Y(_10121_),
    .B1(net9165));
 sg13g2_o21ai_1 _33257_ (.B1(_10121_),
    .Y(_10122_),
    .A1(net9153),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][26] ));
 sg13g2_a22oi_1 _33258_ (.Y(_10123_),
    .B1(net8904),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][26] ),
    .A2(net8793),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][26] ));
 sg13g2_nand3_1 _33259_ (.B(_10122_),
    .C(_10123_),
    .A(net9472),
    .Y(_10124_));
 sg13g2_nand3_1 _33260_ (.B(_10120_),
    .C(_10124_),
    .A(net9448),
    .Y(_10125_));
 sg13g2_nor2_1 _33261_ (.A(net9153),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][26] ),
    .Y(_10126_));
 sg13g2_o21ai_1 _33262_ (.B1(net9507),
    .Y(_10127_),
    .A1(net9542),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][26] ));
 sg13g2_a22oi_1 _33263_ (.Y(_10128_),
    .B1(net8904),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][26] ),
    .A2(net8793),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][26] ));
 sg13g2_o21ai_1 _33264_ (.B1(_10128_),
    .Y(_10129_),
    .A1(_10126_),
    .A2(_10127_));
 sg13g2_o21ai_1 _33265_ (.B1(net9503),
    .Y(_10130_),
    .A1(net9538),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][26] ));
 sg13g2_a21oi_1 _33266_ (.A1(net9538),
    .A2(_10797_),
    .Y(_10131_),
    .B1(_10130_));
 sg13g2_a221oi_1 _33267_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][26] ),
    .C1(_10131_),
    .B1(net8898),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][26] ),
    .Y(_10132_),
    .A2(net8788));
 sg13g2_o21ai_1 _33268_ (.B1(net9436),
    .Y(_10133_),
    .A1(net8913),
    .A2(_10132_));
 sg13g2_a21oi_1 _33269_ (.A1(net8926),
    .A2(_10129_),
    .Y(_10134_),
    .B1(_10133_));
 sg13g2_a221oi_1 _33270_ (.B2(_10134_),
    .C1(_09316_),
    .B1(_10125_),
    .A1(_10107_),
    .Y(_02707_),
    .A2(_10116_));
 sg13g2_a21oi_1 _33271_ (.A1(net9132),
    .A2(_10799_),
    .Y(_10135_),
    .B1(net9161));
 sg13g2_o21ai_1 _33272_ (.B1(_10135_),
    .Y(_10136_),
    .A1(net9129),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][27] ));
 sg13g2_a221oi_1 _33273_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][27] ),
    .C1(net9458),
    .B1(net8875),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][27] ),
    .Y(_10137_),
    .A2(net8764));
 sg13g2_mux2_1 _33274_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][27] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][27] ),
    .S(net9521),
    .X(_10138_));
 sg13g2_a22oi_1 _33275_ (.Y(_10139_),
    .B1(net8875),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][27] ),
    .A2(net8763),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][27] ));
 sg13g2_nand2_1 _33276_ (.Y(_10140_),
    .A(net9458),
    .B(_10139_));
 sg13g2_a21oi_1 _33277_ (.A1(net9486),
    .A2(_10138_),
    .Y(_10141_),
    .B1(_10140_));
 sg13g2_a21oi_1 _33278_ (.A1(_10136_),
    .A2(_10137_),
    .Y(_10142_),
    .B1(_10141_));
 sg13g2_nor2_1 _33279_ (.A(net9521),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][27] ),
    .Y(_10143_));
 sg13g2_o21ai_1 _33280_ (.B1(net9487),
    .Y(_10144_),
    .A1(net9129),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][27] ));
 sg13g2_a22oi_1 _33281_ (.Y(_10145_),
    .B1(net8874),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][27] ),
    .A2(net8764),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][27] ));
 sg13g2_o21ai_1 _33282_ (.B1(_10145_),
    .Y(_10146_),
    .A1(_10143_),
    .A2(_10144_));
 sg13g2_mux2_1 _33283_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][27] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][27] ),
    .S(net9521),
    .X(_10147_));
 sg13g2_nand2_1 _33284_ (.Y(_10148_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][27] ),
    .B(net8874));
 sg13g2_a22oi_1 _33285_ (.Y(_10149_),
    .B1(_10147_),
    .B2(net9486),
    .A2(net8763),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][27] ));
 sg13g2_a21oi_1 _33286_ (.A1(_10148_),
    .A2(_10149_),
    .Y(_10150_),
    .B1(net8910));
 sg13g2_a221oi_1 _33287_ (.B2(net8924),
    .C1(_10150_),
    .B1(_10146_),
    .A1(net9443),
    .Y(_10151_),
    .A2(_10142_));
 sg13g2_a21oi_1 _33288_ (.A1(net9129),
    .A2(_10801_),
    .Y(_10152_),
    .B1(net9161));
 sg13g2_o21ai_1 _33289_ (.B1(_10152_),
    .Y(_10153_),
    .A1(net9129),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][27] ));
 sg13g2_a22oi_1 _33290_ (.Y(_10154_),
    .B1(net8875),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][27] ),
    .A2(net8764),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][27] ));
 sg13g2_nand3_1 _33291_ (.B(_10153_),
    .C(_10154_),
    .A(net9458),
    .Y(_10155_));
 sg13g2_nor2_1 _33292_ (.A(net9521),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][27] ),
    .Y(_10156_));
 sg13g2_o21ai_1 _33293_ (.B1(net9486),
    .Y(_10157_),
    .A1(net9129),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][27] ));
 sg13g2_a221oi_1 _33294_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][27] ),
    .C1(net9458),
    .B1(net8874),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][27] ),
    .Y(_10158_),
    .A2(net8763));
 sg13g2_o21ai_1 _33295_ (.B1(_10158_),
    .Y(_10159_),
    .A1(_10156_),
    .A2(_10157_));
 sg13g2_nand3_1 _33296_ (.B(_10155_),
    .C(_10159_),
    .A(net9443),
    .Y(_10160_));
 sg13g2_mux2_1 _33297_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][27] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][27] ),
    .S(net9521),
    .X(_10161_));
 sg13g2_nand2_1 _33298_ (.Y(_10162_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][27] ),
    .B(net8874));
 sg13g2_a22oi_1 _33299_ (.Y(_10163_),
    .B1(_10161_),
    .B2(net9486),
    .A2(net8763),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][27] ));
 sg13g2_a21oi_1 _33300_ (.A1(_10162_),
    .A2(_10163_),
    .Y(_10164_),
    .B1(net8918));
 sg13g2_o21ai_1 _33301_ (.B1(net9486),
    .Y(_10165_),
    .A1(net9129),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][27] ));
 sg13g2_a21oi_1 _33302_ (.A1(net9129),
    .A2(_10800_),
    .Y(_10166_),
    .B1(_10165_));
 sg13g2_a221oi_1 _33303_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][27] ),
    .C1(_10166_),
    .B1(net8874),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][27] ),
    .Y(_10167_),
    .A2(net8763));
 sg13g2_o21ai_1 _33304_ (.B1(_10160_),
    .Y(_10168_),
    .A1(net8909),
    .A2(_10167_));
 sg13g2_o21ai_1 _33305_ (.B1(net9434),
    .Y(_10169_),
    .A1(_10164_),
    .A2(_10168_));
 sg13g2_o21ai_1 _33306_ (.B1(_10169_),
    .Y(_02708_),
    .A1(net8745),
    .A2(_10151_));
 sg13g2_mux2_1 _33307_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][28] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][28] ),
    .S(net9523),
    .X(_10170_));
 sg13g2_a22oi_1 _33308_ (.Y(_10171_),
    .B1(net8876),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][28] ),
    .A2(net8765),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][28] ));
 sg13g2_nand2_1 _33309_ (.Y(_10172_),
    .A(net9459),
    .B(_10171_));
 sg13g2_a21oi_1 _33310_ (.A1(net9488),
    .A2(_10170_),
    .Y(_10173_),
    .B1(_10172_));
 sg13g2_a21oi_1 _33311_ (.A1(net9131),
    .A2(_10803_),
    .Y(_10174_),
    .B1(net9160));
 sg13g2_o21ai_1 _33312_ (.B1(_10174_),
    .Y(_10175_),
    .A1(net9130),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][28] ));
 sg13g2_a221oi_1 _33313_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][28] ),
    .C1(net9459),
    .B1(net8876),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][28] ),
    .Y(_10176_),
    .A2(net8765));
 sg13g2_a21oi_1 _33314_ (.A1(_10175_),
    .A2(_10176_),
    .Y(_10177_),
    .B1(_10173_));
 sg13g2_nor2_1 _33315_ (.A(net9522),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][28] ),
    .Y(_10178_));
 sg13g2_o21ai_1 _33316_ (.B1(net9487),
    .Y(_10179_),
    .A1(net9130),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][28] ));
 sg13g2_a22oi_1 _33317_ (.Y(_10180_),
    .B1(net8876),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][28] ),
    .A2(net8765),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][28] ));
 sg13g2_o21ai_1 _33318_ (.B1(_10180_),
    .Y(_10181_),
    .A1(_10178_),
    .A2(_10179_));
 sg13g2_mux2_1 _33319_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][28] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][28] ),
    .S(net9522),
    .X(_10182_));
 sg13g2_nand2_1 _33320_ (.Y(_10183_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][28] ),
    .B(net8876));
 sg13g2_a22oi_1 _33321_ (.Y(_10184_),
    .B1(_10182_),
    .B2(net9487),
    .A2(net8765),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][28] ));
 sg13g2_a21oi_1 _33322_ (.A1(_10183_),
    .A2(_10184_),
    .Y(_10185_),
    .B1(net8909));
 sg13g2_a221oi_1 _33323_ (.B2(net8923),
    .C1(_10185_),
    .B1(_10181_),
    .A1(net9442),
    .Y(_10186_),
    .A2(_10177_));
 sg13g2_a21oi_1 _33324_ (.A1(net9130),
    .A2(_10806_),
    .Y(_10187_),
    .B1(net9161));
 sg13g2_o21ai_1 _33325_ (.B1(_10187_),
    .Y(_10188_),
    .A1(net9130),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][28] ));
 sg13g2_a22oi_1 _33326_ (.Y(_10189_),
    .B1(net8876),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][28] ),
    .A2(net8765),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][28] ));
 sg13g2_nand3_1 _33327_ (.B(_10188_),
    .C(_10189_),
    .A(net9459),
    .Y(_10190_));
 sg13g2_nor2_1 _33328_ (.A(net9523),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][28] ),
    .Y(_10191_));
 sg13g2_o21ai_1 _33329_ (.B1(net9488),
    .Y(_10192_),
    .A1(net9130),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][28] ));
 sg13g2_a221oi_1 _33330_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][28] ),
    .C1(net9458),
    .B1(net8876),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][28] ),
    .Y(_10193_),
    .A2(net8765));
 sg13g2_o21ai_1 _33331_ (.B1(_10193_),
    .Y(_10194_),
    .A1(_10191_),
    .A2(_10192_));
 sg13g2_nand3_1 _33332_ (.B(_10190_),
    .C(_10194_),
    .A(net9442),
    .Y(_10195_));
 sg13g2_mux2_1 _33333_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][28] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][28] ),
    .S(net9522),
    .X(_10196_));
 sg13g2_nand2_1 _33334_ (.Y(_10197_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][28] ),
    .B(net8876));
 sg13g2_a22oi_1 _33335_ (.Y(_10198_),
    .B1(_10196_),
    .B2(net9488),
    .A2(net8765),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][28] ));
 sg13g2_a21oi_1 _33336_ (.A1(_10197_),
    .A2(_10198_),
    .Y(_10199_),
    .B1(net8918));
 sg13g2_o21ai_1 _33337_ (.B1(net9487),
    .Y(_10200_),
    .A1(net9130),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][28] ));
 sg13g2_a21oi_1 _33338_ (.A1(net9130),
    .A2(_10804_),
    .Y(_10201_),
    .B1(_10200_));
 sg13g2_a221oi_1 _33339_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][28] ),
    .C1(_10201_),
    .B1(net8877),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][28] ),
    .Y(_10202_),
    .A2(net8766));
 sg13g2_o21ai_1 _33340_ (.B1(_10195_),
    .Y(_10203_),
    .A1(net8909),
    .A2(_10202_));
 sg13g2_o21ai_1 _33341_ (.B1(net9434),
    .Y(_10204_),
    .A1(_10199_),
    .A2(_10203_));
 sg13g2_o21ai_1 _33342_ (.B1(_10204_),
    .Y(_02709_),
    .A1(net8748),
    .A2(_10186_));
 sg13g2_mux2_1 _33343_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][29] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][29] ),
    .S(net9528),
    .X(_10205_));
 sg13g2_a22oi_1 _33344_ (.Y(_10206_),
    .B1(net8882),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][29] ),
    .A2(net8774),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][29] ));
 sg13g2_nand2_1 _33345_ (.Y(_10207_),
    .A(net9464),
    .B(_10206_));
 sg13g2_a21oi_1 _33346_ (.A1(net9492),
    .A2(_10205_),
    .Y(_10208_),
    .B1(_10207_));
 sg13g2_a21oi_1 _33347_ (.A1(net9136),
    .A2(_10808_),
    .Y(_10209_),
    .B1(net9163));
 sg13g2_o21ai_1 _33348_ (.B1(_10209_),
    .Y(_10210_),
    .A1(net9136),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][29] ));
 sg13g2_a221oi_1 _33349_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][29] ),
    .C1(net9464),
    .B1(net8882),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][29] ),
    .Y(_10211_),
    .A2(net8773));
 sg13g2_a21oi_1 _33350_ (.A1(_10210_),
    .A2(_10211_),
    .Y(_10212_),
    .B1(_10208_));
 sg13g2_nor2_1 _33351_ (.A(net9528),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][29] ),
    .Y(_10213_));
 sg13g2_o21ai_1 _33352_ (.B1(net9492),
    .Y(_10214_),
    .A1(net9136),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][29] ));
 sg13g2_a22oi_1 _33353_ (.Y(_10215_),
    .B1(net8882),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][29] ),
    .A2(net8773),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][29] ));
 sg13g2_o21ai_1 _33354_ (.B1(_10215_),
    .Y(_10216_),
    .A1(_10213_),
    .A2(_10214_));
 sg13g2_mux2_1 _33355_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][29] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][29] ),
    .S(net9528),
    .X(_10217_));
 sg13g2_nand2_1 _33356_ (.Y(_10218_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][29] ),
    .B(net8882));
 sg13g2_a22oi_1 _33357_ (.Y(_10219_),
    .B1(_10217_),
    .B2(net9492),
    .A2(net8773),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][29] ));
 sg13g2_a21oi_1 _33358_ (.A1(_10218_),
    .A2(_10219_),
    .Y(_10220_),
    .B1(net8911));
 sg13g2_a221oi_1 _33359_ (.B2(net8925),
    .C1(_10220_),
    .B1(_10216_),
    .A1(net9445),
    .Y(_10221_),
    .A2(_10212_));
 sg13g2_a21oi_1 _33360_ (.A1(net9137),
    .A2(_10810_),
    .Y(_10222_),
    .B1(net9163));
 sg13g2_o21ai_1 _33361_ (.B1(_10222_),
    .Y(_10223_),
    .A1(net9137),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][29] ));
 sg13g2_a22oi_1 _33362_ (.Y(_10224_),
    .B1(net8883),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][29] ),
    .A2(net8774),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][29] ));
 sg13g2_nand3_1 _33363_ (.B(_10223_),
    .C(_10224_),
    .A(net9464),
    .Y(_10225_));
 sg13g2_nor2_1 _33364_ (.A(net9528),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][29] ),
    .Y(_10226_));
 sg13g2_o21ai_1 _33365_ (.B1(net9492),
    .Y(_10227_),
    .A1(net9137),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][29] ));
 sg13g2_a221oi_1 _33366_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][29] ),
    .C1(net9464),
    .B1(net8883),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][29] ),
    .Y(_10228_),
    .A2(net8774));
 sg13g2_o21ai_1 _33367_ (.B1(_10228_),
    .Y(_10229_),
    .A1(_10226_),
    .A2(_10227_));
 sg13g2_nand3_1 _33368_ (.B(_10225_),
    .C(_10229_),
    .A(net9445),
    .Y(_10230_));
 sg13g2_mux2_1 _33369_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][29] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][29] ),
    .S(net9528),
    .X(_10231_));
 sg13g2_nand2_1 _33370_ (.Y(_10232_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][29] ),
    .B(net8882));
 sg13g2_a22oi_1 _33371_ (.Y(_10233_),
    .B1(_10231_),
    .B2(net9492),
    .A2(net8773),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][29] ));
 sg13g2_a21oi_1 _33372_ (.A1(_10232_),
    .A2(_10233_),
    .Y(_10234_),
    .B1(net8921));
 sg13g2_o21ai_1 _33373_ (.B1(net9493),
    .Y(_10235_),
    .A1(net9137),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][29] ));
 sg13g2_a21oi_1 _33374_ (.A1(net9137),
    .A2(_10809_),
    .Y(_10236_),
    .B1(_10235_));
 sg13g2_a221oi_1 _33375_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][29] ),
    .C1(_10236_),
    .B1(net8883),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][29] ),
    .Y(_10237_),
    .A2(net8774));
 sg13g2_o21ai_1 _33376_ (.B1(_10230_),
    .Y(_10238_),
    .A1(net8912),
    .A2(_10237_));
 sg13g2_o21ai_1 _33377_ (.B1(net9439),
    .Y(_10239_),
    .A1(_10234_),
    .A2(_10238_));
 sg13g2_o21ai_1 _33378_ (.B1(_10239_),
    .Y(_02710_),
    .A1(net8746),
    .A2(_10221_));
 sg13g2_mux2_1 _33379_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][30] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][30] ),
    .S(net9521),
    .X(_10240_));
 sg13g2_a22oi_1 _33380_ (.Y(_10241_),
    .B1(net8877),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][30] ),
    .A2(net8767),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][30] ));
 sg13g2_nand2_1 _33381_ (.Y(_10242_),
    .A(net9460),
    .B(_10241_));
 sg13g2_a21oi_1 _33382_ (.A1(net9486),
    .A2(_10240_),
    .Y(_10243_),
    .B1(_10242_));
 sg13g2_a21oi_1 _33383_ (.A1(net9128),
    .A2(_10811_),
    .Y(_10244_),
    .B1(net9160));
 sg13g2_o21ai_1 _33384_ (.B1(_10244_),
    .Y(_10245_),
    .A1(net9128),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][30] ));
 sg13g2_a221oi_1 _33385_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][30] ),
    .C1(net9458),
    .B1(net8874),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][30] ),
    .Y(_10246_),
    .A2(net8763));
 sg13g2_a21oi_1 _33386_ (.A1(_10245_),
    .A2(_10246_),
    .Y(_10247_),
    .B1(_10243_));
 sg13g2_nor2_1 _33387_ (.A(net9519),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][30] ),
    .Y(_10248_));
 sg13g2_o21ai_1 _33388_ (.B1(net9485),
    .Y(_10249_),
    .A1(net9128),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][30] ));
 sg13g2_a22oi_1 _33389_ (.Y(_10250_),
    .B1(net8873),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][30] ),
    .A2(net8762),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][30] ));
 sg13g2_o21ai_1 _33390_ (.B1(_10250_),
    .Y(_10251_),
    .A1(_10248_),
    .A2(_10249_));
 sg13g2_mux2_1 _33391_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][30] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][30] ),
    .S(net9519),
    .X(_10252_));
 sg13g2_nand2_1 _33392_ (.Y(_10253_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][30] ),
    .B(net8873));
 sg13g2_a22oi_1 _33393_ (.Y(_10254_),
    .B1(_10252_),
    .B2(net9485),
    .A2(net8762),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][30] ));
 sg13g2_a21oi_1 _33394_ (.A1(_10253_),
    .A2(_10254_),
    .Y(_10255_),
    .B1(net8909));
 sg13g2_a221oi_1 _33395_ (.B2(net8923),
    .C1(_10255_),
    .B1(_10251_),
    .A1(net9442),
    .Y(_10256_),
    .A2(_10247_));
 sg13g2_a21oi_1 _33396_ (.A1(net9133),
    .A2(_10812_),
    .Y(_10257_),
    .B1(net9160));
 sg13g2_o21ai_1 _33397_ (.B1(_10257_),
    .Y(_10258_),
    .A1(net9128),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][30] ));
 sg13g2_a221oi_1 _33398_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][30] ),
    .C1(net9460),
    .B1(net8873),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][30] ),
    .Y(_10259_),
    .A2(net8762));
 sg13g2_o21ai_1 _33399_ (.B1(net9488),
    .Y(_10260_),
    .A1(net9520),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][30] ));
 sg13g2_a21oi_1 _33400_ (.A1(net9519),
    .A2(_10813_),
    .Y(_10261_),
    .B1(_10260_));
 sg13g2_a221oi_1 _33401_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][30] ),
    .C1(_10261_),
    .B1(net8873),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][30] ),
    .Y(_10262_),
    .A2(net8762));
 sg13g2_a22oi_1 _33402_ (.Y(_10263_),
    .B1(_10262_),
    .B2(net9457),
    .A2(_10259_),
    .A1(_10258_));
 sg13g2_nor2_1 _33403_ (.A(net9519),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][30] ),
    .Y(_10264_));
 sg13g2_o21ai_1 _33404_ (.B1(net9485),
    .Y(_10265_),
    .A1(net9128),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][30] ));
 sg13g2_a22oi_1 _33405_ (.Y(_10266_),
    .B1(net8873),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][30] ),
    .A2(net8762),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][30] ));
 sg13g2_o21ai_1 _33406_ (.B1(_10266_),
    .Y(_10267_),
    .A1(_10264_),
    .A2(_10265_));
 sg13g2_mux2_1 _33407_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][30] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][30] ),
    .S(net9519),
    .X(_10268_));
 sg13g2_nand2_1 _33408_ (.Y(_10269_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][30] ),
    .B(net8873));
 sg13g2_a22oi_1 _33409_ (.Y(_10270_),
    .B1(_10268_),
    .B2(net9485),
    .A2(net8762),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][30] ));
 sg13g2_a21oi_1 _33410_ (.A1(_10269_),
    .A2(_10270_),
    .Y(_10271_),
    .B1(net8909));
 sg13g2_a221oi_1 _33411_ (.B2(net8924),
    .C1(_10271_),
    .B1(_10267_),
    .A1(net9442),
    .Y(_10272_),
    .A2(_10263_));
 sg13g2_nand2b_1 _33412_ (.Y(_10273_),
    .B(net9435),
    .A_N(_10272_));
 sg13g2_o21ai_1 _33413_ (.B1(_10273_),
    .Y(_02711_),
    .A1(net8748),
    .A2(_10256_));
 sg13g2_nor2_1 _33414_ (.A(net9515),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][31] ),
    .Y(_10274_));
 sg13g2_o21ai_1 _33415_ (.B1(net9482),
    .Y(_10275_),
    .A1(net9121),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][31] ));
 sg13g2_a221oi_1 _33416_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][31] ),
    .C1(net9453),
    .B1(net8868),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][31] ),
    .Y(_10276_),
    .A2(net8758));
 sg13g2_o21ai_1 _33417_ (.B1(_10276_),
    .Y(_10277_),
    .A1(_10274_),
    .A2(_10275_));
 sg13g2_a21oi_1 _33418_ (.A1(net9125),
    .A2(_10817_),
    .Y(_10278_),
    .B1(net9159));
 sg13g2_o21ai_1 _33419_ (.B1(_10278_),
    .Y(_10279_),
    .A1(net9125),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][31] ));
 sg13g2_a22oi_1 _33420_ (.Y(_10280_),
    .B1(net8870),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][31] ),
    .A2(net8760),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][31] ));
 sg13g2_nand3_1 _33421_ (.B(_10279_),
    .C(_10280_),
    .A(net9456),
    .Y(_10281_));
 sg13g2_nand3_1 _33422_ (.B(_10277_),
    .C(_10281_),
    .A(net9443),
    .Y(_10282_));
 sg13g2_o21ai_1 _33423_ (.B1(net9481),
    .Y(_10283_),
    .A1(net9515),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][31] ));
 sg13g2_a21oi_1 _33424_ (.A1(net9515),
    .A2(_10816_),
    .Y(_10284_),
    .B1(_10283_));
 sg13g2_a221oi_1 _33425_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][31] ),
    .C1(_10284_),
    .B1(net8866),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][31] ),
    .Y(_10285_),
    .A2(net8757));
 sg13g2_nor2_1 _33426_ (.A(net9122),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][31] ),
    .Y(_10286_));
 sg13g2_o21ai_1 _33427_ (.B1(net9481),
    .Y(_10287_),
    .A1(net9515),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][31] ));
 sg13g2_a22oi_1 _33428_ (.Y(_10288_),
    .B1(net8866),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][31] ),
    .A2(net8756),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][31] ));
 sg13g2_o21ai_1 _33429_ (.B1(_10288_),
    .Y(_10289_),
    .A1(_10286_),
    .A2(_10287_));
 sg13g2_o21ai_1 _33430_ (.B1(net9432),
    .Y(_10290_),
    .A1(net8907),
    .A2(_10285_));
 sg13g2_a21oi_1 _33431_ (.A1(net8922),
    .A2(_10289_),
    .Y(_10291_),
    .B1(_10290_));
 sg13g2_nor2_1 _33432_ (.A(net9517),
    .B(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][31] ),
    .Y(_10292_));
 sg13g2_o21ai_1 _33433_ (.B1(net9483),
    .Y(_10293_),
    .A1(net9125),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][31] ));
 sg13g2_a221oi_1 _33434_ (.B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][31] ),
    .C1(net9456),
    .B1(net8869),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][31] ),
    .Y(_10294_),
    .A2(net8759));
 sg13g2_o21ai_1 _33435_ (.B1(_10294_),
    .Y(_10295_),
    .A1(_10292_),
    .A2(_10293_));
 sg13g2_a21oi_1 _33436_ (.A1(net9126),
    .A2(_10815_),
    .Y(_10296_),
    .B1(net9159));
 sg13g2_o21ai_1 _33437_ (.B1(_10296_),
    .Y(_10297_),
    .A1(net9125),
    .A2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][31] ));
 sg13g2_a22oi_1 _33438_ (.Y(_10298_),
    .B1(net8870),
    .B2(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][31] ),
    .A2(net8760),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][31] ));
 sg13g2_nand3_1 _33439_ (.B(_10297_),
    .C(_10298_),
    .A(net9456),
    .Y(_10299_));
 sg13g2_nand3_1 _33440_ (.B(_10295_),
    .C(_10299_),
    .A(net9443),
    .Y(_10300_));
 sg13g2_mux2_1 _33441_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][31] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][31] ),
    .S(net9515),
    .X(_10301_));
 sg13g2_nand2_1 _33442_ (.Y(_10302_),
    .A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][31] ),
    .B(net8867));
 sg13g2_a22oi_1 _33443_ (.Y(_10303_),
    .B1(_10301_),
    .B2(net9481),
    .A2(net8756),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][31] ));
 sg13g2_a21oi_1 _33444_ (.A1(_10302_),
    .A2(_10303_),
    .Y(_10304_),
    .B1(net8907));
 sg13g2_mux2_1 _33445_ (.A0(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][31] ),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][31] ),
    .S(net9517),
    .X(_10305_));
 sg13g2_a22oi_1 _33446_ (.Y(_10306_),
    .B1(_10305_),
    .B2(net9481),
    .A2(net8756),
    .A1(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][31] ));
 sg13g2_nor3_1 _33447_ (.A(net8917),
    .B(net8866),
    .C(_10306_),
    .Y(_10307_));
 sg13g2_nor3_1 _33448_ (.A(net9432),
    .B(_10304_),
    .C(_10307_),
    .Y(_10308_));
 sg13g2_a22oi_1 _33449_ (.Y(_02712_),
    .B1(_10300_),
    .B2(_10308_),
    .A2(_10291_),
    .A1(_10282_));
 sg13g2_nand2_1 _33450_ (.Y(_10309_),
    .A(net8961),
    .B(_08924_));
 sg13g2_nand2_1 _33451_ (.Y(_10310_),
    .A(net2934),
    .B(net7953));
 sg13g2_o21ai_1 _33452_ (.B1(_10310_),
    .Y(_02713_),
    .A1(net7485),
    .A2(net7953));
 sg13g2_nand2_1 _33453_ (.Y(_10311_),
    .A(net3672),
    .B(net7956));
 sg13g2_o21ai_1 _33454_ (.B1(_10311_),
    .Y(_02714_),
    .A1(net7664),
    .A2(net7954));
 sg13g2_nand2_1 _33455_ (.Y(_10312_),
    .A(net2923),
    .B(net7954));
 sg13g2_o21ai_1 _33456_ (.B1(_10312_),
    .Y(_02715_),
    .A1(net7615),
    .A2(net7954));
 sg13g2_nand2_1 _33457_ (.Y(_10313_),
    .A(net4108),
    .B(net7955));
 sg13g2_o21ai_1 _33458_ (.B1(_10313_),
    .Y(_02716_),
    .A1(net7608),
    .A2(net7955));
 sg13g2_nand2_1 _33459_ (.Y(_10314_),
    .A(net3750),
    .B(net7953));
 sg13g2_o21ai_1 _33460_ (.B1(_10314_),
    .Y(_02717_),
    .A1(net7590),
    .A2(net7953));
 sg13g2_nand2_1 _33461_ (.Y(_10315_),
    .A(net3407),
    .B(net7957));
 sg13g2_o21ai_1 _33462_ (.B1(_10315_),
    .Y(_02718_),
    .A1(net7599),
    .A2(net7957));
 sg13g2_nand2_1 _33463_ (.Y(_10316_),
    .A(net2911),
    .B(net7955));
 sg13g2_o21ai_1 _33464_ (.B1(_10316_),
    .Y(_02719_),
    .A1(net7592),
    .A2(net7955));
 sg13g2_nand2_1 _33465_ (.Y(_10317_),
    .A(net3417),
    .B(net7951));
 sg13g2_o21ai_1 _33466_ (.B1(_10317_),
    .Y(_02720_),
    .A1(net7606),
    .A2(net7950));
 sg13g2_nand2_1 _33467_ (.Y(_10318_),
    .A(net3877),
    .B(net7957));
 sg13g2_o21ai_1 _33468_ (.B1(_10318_),
    .Y(_02721_),
    .A1(net7561),
    .A2(net7957));
 sg13g2_nand2_1 _33469_ (.Y(_10319_),
    .A(net2833),
    .B(net7954));
 sg13g2_o21ai_1 _33470_ (.B1(_10319_),
    .Y(_02722_),
    .A1(net7578),
    .A2(net7954));
 sg13g2_nand2_1 _33471_ (.Y(_10320_),
    .A(net2931),
    .B(net7956));
 sg13g2_o21ai_1 _33472_ (.B1(_10320_),
    .Y(_02723_),
    .A1(net7549),
    .A2(net7956));
 sg13g2_nand2_1 _33473_ (.Y(_10321_),
    .A(net3121),
    .B(net7949));
 sg13g2_o21ai_1 _33474_ (.B1(_10321_),
    .Y(_02724_),
    .A1(net7571),
    .A2(net7949));
 sg13g2_nand2_1 _33475_ (.Y(_10322_),
    .A(net3658),
    .B(net7954));
 sg13g2_o21ai_1 _33476_ (.B1(_10322_),
    .Y(_02725_),
    .A1(net7540),
    .A2(net7958));
 sg13g2_nand2_1 _33477_ (.Y(_10323_),
    .A(net3276),
    .B(net7954));
 sg13g2_o21ai_1 _33478_ (.B1(_10323_),
    .Y(_02726_),
    .A1(net7554),
    .A2(net7954));
 sg13g2_nand2_1 _33479_ (.Y(_10324_),
    .A(net3519),
    .B(net7951));
 sg13g2_o21ai_1 _33480_ (.B1(_10324_),
    .Y(_02727_),
    .A1(net7581),
    .A2(net7951));
 sg13g2_nand2_1 _33481_ (.Y(_10325_),
    .A(net3436),
    .B(net7949));
 sg13g2_o21ai_1 _33482_ (.B1(_10325_),
    .Y(_02728_),
    .A1(net7565),
    .A2(net7950));
 sg13g2_nand2_1 _33483_ (.Y(_10326_),
    .A(net3032),
    .B(net7949));
 sg13g2_o21ai_1 _33484_ (.B1(_10326_),
    .Y(_02729_),
    .A1(net7524),
    .A2(net7949));
 sg13g2_nand2_1 _33485_ (.Y(_10327_),
    .A(net2897),
    .B(net7949));
 sg13g2_o21ai_1 _33486_ (.B1(_10327_),
    .Y(_02730_),
    .A1(net7539),
    .A2(net7949));
 sg13g2_nand2_1 _33487_ (.Y(_10328_),
    .A(net3952),
    .B(net7950));
 sg13g2_o21ai_1 _33488_ (.B1(_10328_),
    .Y(_02731_),
    .A1(net7530),
    .A2(net7950));
 sg13g2_nand2_1 _33489_ (.Y(_10329_),
    .A(net3383),
    .B(net7951));
 sg13g2_o21ai_1 _33490_ (.B1(_10329_),
    .Y(_02732_),
    .A1(net7521),
    .A2(net7951));
 sg13g2_nand2_1 _33491_ (.Y(_10330_),
    .A(net3265),
    .B(net7953));
 sg13g2_o21ai_1 _33492_ (.B1(_10330_),
    .Y(_02733_),
    .A1(net7508),
    .A2(net7953));
 sg13g2_nand2_1 _33493_ (.Y(_10331_),
    .A(net3845),
    .B(net7952));
 sg13g2_o21ai_1 _33494_ (.B1(_10331_),
    .Y(_02734_),
    .A1(net7511),
    .A2(net7952));
 sg13g2_nand2_1 _33495_ (.Y(_10332_),
    .A(net2926),
    .B(net7955));
 sg13g2_o21ai_1 _33496_ (.B1(_10332_),
    .Y(_02735_),
    .A1(net7497),
    .A2(net7955));
 sg13g2_nand2_1 _33497_ (.Y(_10333_),
    .A(net3024),
    .B(net7950));
 sg13g2_o21ai_1 _33498_ (.B1(_10333_),
    .Y(_02736_),
    .A1(net7499),
    .A2(net7949));
 sg13g2_nand2_1 _33499_ (.Y(_10334_),
    .A(net3805),
    .B(net7957));
 sg13g2_o21ai_1 _33500_ (.B1(_10334_),
    .Y(_02737_),
    .A1(net7642),
    .A2(net7957));
 sg13g2_nand2_1 _33501_ (.Y(_10335_),
    .A(net3084),
    .B(net7953));
 sg13g2_o21ai_1 _33502_ (.B1(_10335_),
    .Y(_02738_),
    .A1(net7650),
    .A2(net7953));
 sg13g2_nand2_1 _33503_ (.Y(_10336_),
    .A(net3793),
    .B(net7955));
 sg13g2_o21ai_1 _33504_ (.B1(_10336_),
    .Y(_02739_),
    .A1(net7653),
    .A2(net7955));
 sg13g2_nand2_1 _33505_ (.Y(_10337_),
    .A(net3838),
    .B(net7952));
 sg13g2_o21ai_1 _33506_ (.B1(_10337_),
    .Y(_02740_),
    .A1(net7659),
    .A2(net7952));
 sg13g2_nand2_1 _33507_ (.Y(_10338_),
    .A(net3342),
    .B(net7952));
 sg13g2_o21ai_1 _33508_ (.B1(_10338_),
    .Y(_02741_),
    .A1(net7637),
    .A2(net7952));
 sg13g2_nand2_1 _33509_ (.Y(_10339_),
    .A(net3019),
    .B(net7957));
 sg13g2_o21ai_1 _33510_ (.B1(_10339_),
    .Y(_02742_),
    .A1(net7627),
    .A2(net7957));
 sg13g2_nand2_1 _33511_ (.Y(_10340_),
    .A(net4175),
    .B(net7958));
 sg13g2_o21ai_1 _33512_ (.B1(_10340_),
    .Y(_02743_),
    .A1(net7622),
    .A2(net7952));
 sg13g2_nand2_1 _33513_ (.Y(_10341_),
    .A(net3221),
    .B(net7950));
 sg13g2_o21ai_1 _33514_ (.B1(_10341_),
    .Y(_02744_),
    .A1(net7631),
    .A2(net7950));
 sg13g2_nand2_1 _33515_ (.Y(_10342_),
    .A(_14126_),
    .B(_08924_));
 sg13g2_nand2_1 _33516_ (.Y(_10343_),
    .A(net3061),
    .B(net7947));
 sg13g2_o21ai_1 _33517_ (.B1(_10343_),
    .Y(_02745_),
    .A1(net7485),
    .A2(net7947));
 sg13g2_nand2_1 _33518_ (.Y(_10344_),
    .A(net2637),
    .B(net7944));
 sg13g2_o21ai_1 _33519_ (.B1(_10344_),
    .Y(_02746_),
    .A1(net7666),
    .A2(net7945));
 sg13g2_nand2_1 _33520_ (.Y(_10345_),
    .A(net2673),
    .B(net7945));
 sg13g2_o21ai_1 _33521_ (.B1(_10345_),
    .Y(_02747_),
    .A1(net7615),
    .A2(net7945));
 sg13g2_nand2_1 _33522_ (.Y(_10346_),
    .A(net3470),
    .B(net7945));
 sg13g2_o21ai_1 _33523_ (.B1(_10346_),
    .Y(_02748_),
    .A1(net7608),
    .A2(net7944));
 sg13g2_nand2_1 _33524_ (.Y(_10347_),
    .A(net3633),
    .B(net7947));
 sg13g2_o21ai_1 _33525_ (.B1(_10347_),
    .Y(_02749_),
    .A1(net7590),
    .A2(net7947));
 sg13g2_nand2_1 _33526_ (.Y(_10348_),
    .A(net3162),
    .B(net7943));
 sg13g2_o21ai_1 _33527_ (.B1(_10348_),
    .Y(_02750_),
    .A1(net7599),
    .A2(net7943));
 sg13g2_nand2_1 _33528_ (.Y(_10349_),
    .A(net3283),
    .B(net7948));
 sg13g2_o21ai_1 _33529_ (.B1(_10349_),
    .Y(_02751_),
    .A1(net7592),
    .A2(net7948));
 sg13g2_nand2_1 _33530_ (.Y(_10350_),
    .A(net3294),
    .B(net7941));
 sg13g2_o21ai_1 _33531_ (.B1(_10350_),
    .Y(_02752_),
    .A1(net7605),
    .A2(net7941));
 sg13g2_nand2_1 _33532_ (.Y(_10351_),
    .A(net3214),
    .B(net7948));
 sg13g2_o21ai_1 _33533_ (.B1(_10351_),
    .Y(_02753_),
    .A1(net7561),
    .A2(net7948));
 sg13g2_nand2_1 _33534_ (.Y(_10352_),
    .A(net3243),
    .B(net7944));
 sg13g2_o21ai_1 _33535_ (.B1(_10352_),
    .Y(_02754_),
    .A1(net7578),
    .A2(net7944));
 sg13g2_nand2_1 _33536_ (.Y(_10353_),
    .A(net2905),
    .B(net7946));
 sg13g2_o21ai_1 _33537_ (.B1(_10353_),
    .Y(_02755_),
    .A1(net7549),
    .A2(net7946));
 sg13g2_nand2_1 _33538_ (.Y(_10354_),
    .A(net4425),
    .B(net7939));
 sg13g2_o21ai_1 _33539_ (.B1(_10354_),
    .Y(_02756_),
    .A1(net7570),
    .A2(net7939));
 sg13g2_nand2_1 _33540_ (.Y(_10355_),
    .A(net2735),
    .B(net7944));
 sg13g2_o21ai_1 _33541_ (.B1(_10355_),
    .Y(_02757_),
    .A1(net7545),
    .A2(net7944));
 sg13g2_nand2_1 _33542_ (.Y(_10356_),
    .A(net2629),
    .B(net7944));
 sg13g2_o21ai_1 _33543_ (.B1(_10356_),
    .Y(_02758_),
    .A1(net7554),
    .A2(net7944));
 sg13g2_nand2_1 _33544_ (.Y(_10357_),
    .A(net3955),
    .B(net7940));
 sg13g2_o21ai_1 _33545_ (.B1(_10357_),
    .Y(_02759_),
    .A1(net7581),
    .A2(net7940));
 sg13g2_nand2_1 _33546_ (.Y(_10358_),
    .A(net3376),
    .B(net7941));
 sg13g2_o21ai_1 _33547_ (.B1(_10358_),
    .Y(_02760_),
    .A1(net7564),
    .A2(net7941));
 sg13g2_nand2_1 _33548_ (.Y(_10359_),
    .A(net2675),
    .B(net7939));
 sg13g2_o21ai_1 _33549_ (.B1(_10359_),
    .Y(_02761_),
    .A1(net7524),
    .A2(net7939));
 sg13g2_nand2_1 _33550_ (.Y(_10360_),
    .A(net2889),
    .B(net7939));
 sg13g2_o21ai_1 _33551_ (.B1(_10360_),
    .Y(_02762_),
    .A1(net7536),
    .A2(net7939));
 sg13g2_nand2_1 _33552_ (.Y(_10361_),
    .A(net3133),
    .B(net7940));
 sg13g2_o21ai_1 _33553_ (.B1(_10361_),
    .Y(_02763_),
    .A1(net7531),
    .A2(net7940));
 sg13g2_nand2_1 _33554_ (.Y(_10362_),
    .A(net2672),
    .B(net7940));
 sg13g2_o21ai_1 _33555_ (.B1(_10362_),
    .Y(_02764_),
    .A1(net7519),
    .A2(net7940));
 sg13g2_nand2_1 _33556_ (.Y(_10363_),
    .A(net2734),
    .B(net7947));
 sg13g2_o21ai_1 _33557_ (.B1(_10363_),
    .Y(_02765_),
    .A1(net7506),
    .A2(net7947));
 sg13g2_nand2_1 _33558_ (.Y(_10364_),
    .A(net2717),
    .B(net7943));
 sg13g2_o21ai_1 _33559_ (.B1(_10364_),
    .Y(_02766_),
    .A1(net7511),
    .A2(net7943));
 sg13g2_nand2_1 _33560_ (.Y(_10365_),
    .A(net2702),
    .B(net7946));
 sg13g2_o21ai_1 _33561_ (.B1(_10365_),
    .Y(_02767_),
    .A1(net7497),
    .A2(net7946));
 sg13g2_nand2_1 _33562_ (.Y(_10366_),
    .A(net3188),
    .B(net7939));
 sg13g2_o21ai_1 _33563_ (.B1(_10366_),
    .Y(_02768_),
    .A1(net7500),
    .A2(net7939));
 sg13g2_nand2_1 _33564_ (.Y(_10367_),
    .A(net3794),
    .B(net7943));
 sg13g2_o21ai_1 _33565_ (.B1(_10367_),
    .Y(_02769_),
    .A1(net7642),
    .A2(net7943));
 sg13g2_nand2_1 _33566_ (.Y(_10368_),
    .A(net2712),
    .B(net7947));
 sg13g2_o21ai_1 _33567_ (.B1(_10368_),
    .Y(_02770_),
    .A1(net7651),
    .A2(net7947));
 sg13g2_nand2_1 _33568_ (.Y(_10369_),
    .A(net3023),
    .B(net7946));
 sg13g2_o21ai_1 _33569_ (.B1(_10369_),
    .Y(_02771_),
    .A1(net7653),
    .A2(net7946));
 sg13g2_nand2_1 _33570_ (.Y(_10370_),
    .A(net3515),
    .B(net7942));
 sg13g2_o21ai_1 _33571_ (.B1(_10370_),
    .Y(_02772_),
    .A1(net7658),
    .A2(net7942));
 sg13g2_nand2_1 _33572_ (.Y(_10371_),
    .A(net2646),
    .B(net7942));
 sg13g2_o21ai_1 _33573_ (.B1(_10371_),
    .Y(_02773_),
    .A1(net7637),
    .A2(net7942));
 sg13g2_nand2_1 _33574_ (.Y(_10372_),
    .A(net3451),
    .B(net7943));
 sg13g2_o21ai_1 _33575_ (.B1(_10372_),
    .Y(_02774_),
    .A1(net7627),
    .A2(net7943));
 sg13g2_nand2_1 _33576_ (.Y(_10373_),
    .A(net3218),
    .B(net7942));
 sg13g2_o21ai_1 _33577_ (.B1(_10373_),
    .Y(_02775_),
    .A1(net7621),
    .A2(net7942));
 sg13g2_nand2_1 _33578_ (.Y(_10374_),
    .A(net2795),
    .B(net7940));
 sg13g2_o21ai_1 _33579_ (.B1(_10374_),
    .Y(_02776_),
    .A1(net7634),
    .A2(net7940));
 sg13g2_a21oi_1 _33580_ (.A1(net3926),
    .A2(_06645_),
    .Y(_02777_),
    .B1(_06953_));
 sg13g2_buf_1 _33581_ (.A(net2947),
    .X(_02617_));
 sg13g2_buf_1 _33582_ (.A(net2636),
    .X(_02618_));
 sg13g2_buf_1 _33583_ (.A(net2704),
    .X(_02619_));
 sg13g2_buf_1 _33584_ (.A(net2623),
    .X(_02620_));
 sg13g2_buf_1 _33585_ (.A(net2756),
    .X(_02621_));
 sg13g2_buf_1 _33586_ (.A(net2628),
    .X(_02622_));
 sg13g2_buf_1 _33587_ (.A(net2614),
    .X(_02623_));
 sg13g2_buf_1 _33588_ (.A(net3357),
    .X(_02624_));
 sg13g2_buf_1 _33589_ (.A(net3057),
    .X(_02625_));
 sg13g2_buf_1 _33590_ (.A(net2612),
    .X(_02626_));
 sg13g2_buf_1 _33591_ (.A(net2757),
    .X(_02627_));
 sg13g2_buf_1 _33592_ (.A(net2666),
    .X(_02628_));
 sg13g2_buf_1 _33593_ (.A(net2835),
    .X(_02629_));
 sg13g2_buf_1 _33594_ (.A(net2764),
    .X(_02630_));
 sg13g2_buf_1 _33595_ (.A(net2876),
    .X(_02631_));
 sg13g2_buf_1 _33596_ (.A(net2615),
    .X(_02632_));
 sg13g2_buf_1 _33597_ (.A(net2619),
    .X(_02633_));
 sg13g2_buf_1 _33598_ (.A(net2714),
    .X(_02634_));
 sg13g2_buf_1 _33599_ (.A(net2707),
    .X(_02635_));
 sg13g2_buf_1 _33600_ (.A(net2618),
    .X(_02636_));
 sg13g2_buf_1 _33601_ (.A(net2684),
    .X(_02637_));
 sg13g2_buf_1 _33602_ (.A(net2688),
    .X(_02638_));
 sg13g2_buf_1 _33603_ (.A(net2727),
    .X(_02639_));
 sg13g2_buf_1 _33604_ (.A(net2724),
    .X(_02640_));
 sg13g2_buf_1 _33605_ (.A(net2674),
    .X(_02641_));
 sg13g2_buf_1 _33606_ (.A(net2613),
    .X(_02642_));
 sg13g2_buf_1 _33607_ (.A(net2659),
    .X(_02643_));
 sg13g2_buf_1 _33608_ (.A(net2809),
    .X(_02644_));
 sg13g2_buf_1 _33609_ (.A(net2653),
    .X(_02645_));
 sg13g2_buf_1 _33610_ (.A(net2692),
    .X(_02646_));
 sg13g2_buf_1 _33611_ (.A(net2700),
    .X(_02647_));
 sg13g2_buf_1 _33612_ (.A(net2610),
    .X(_02648_));
 sg13g2_nor2_1 _33613_ (.A(net3908),
    .B(_06956_),
    .Y(_02778_));
 sg13g2_and3_1 _33614_ (.X(_02779_),
    .A(net9298),
    .B(_06957_),
    .C(net3577));
 sg13g2_a21oi_1 _33615_ (.A1(_10389_),
    .A2(_06958_),
    .Y(_02780_),
    .B1(_06959_));
 sg13g2_dfrbp_1 _33616_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1308),
    .D(_00306_),
    .Q_N(_00076_),
    .Q(\soc_I.clint_I.mtimecmp[40] ));
 sg13g2_dfrbp_1 _33617_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2320),
    .D(_00307_),
    .Q_N(_00080_),
    .Q(\soc_I.clint_I.mtimecmp[41] ));
 sg13g2_dfrbp_1 _33618_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2318),
    .D(_00308_),
    .Q_N(_00084_),
    .Q(\soc_I.clint_I.mtimecmp[42] ));
 sg13g2_dfrbp_1 _33619_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2316),
    .D(_00309_),
    .Q_N(_00088_),
    .Q(\soc_I.clint_I.mtimecmp[43] ));
 sg13g2_dfrbp_1 _33620_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2314),
    .D(_00310_),
    .Q_N(_00092_),
    .Q(\soc_I.clint_I.mtimecmp[44] ));
 sg13g2_dfrbp_1 _33621_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2312),
    .D(_00311_),
    .Q_N(_00096_),
    .Q(\soc_I.clint_I.mtimecmp[45] ));
 sg13g2_dfrbp_1 _33622_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2310),
    .D(_00312_),
    .Q_N(_00100_),
    .Q(\soc_I.clint_I.mtimecmp[46] ));
 sg13g2_dfrbp_1 _33623_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2308),
    .D(_00313_),
    .Q_N(_00104_),
    .Q(\soc_I.clint_I.mtimecmp[47] ));
 sg13g2_dfrbp_1 _33624_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net2306),
    .D(_00314_),
    .Q_N(_00014_),
    .Q(\soc_I.clint_I.mtimecmp[48] ));
 sg13g2_dfrbp_1 _33625_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net2304),
    .D(_00315_),
    .Q_N(_00021_),
    .Q(\soc_I.clint_I.mtimecmp[49] ));
 sg13g2_dfrbp_1 _33626_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2302),
    .D(_00316_),
    .Q_N(_00029_),
    .Q(\soc_I.clint_I.mtimecmp[50] ));
 sg13g2_dfrbp_1 _33627_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net2300),
    .D(_00317_),
    .Q_N(_00037_),
    .Q(\soc_I.clint_I.mtimecmp[51] ));
 sg13g2_dfrbp_1 _33628_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2298),
    .D(_00318_),
    .Q_N(_00044_),
    .Q(\soc_I.clint_I.mtimecmp[52] ));
 sg13g2_dfrbp_1 _33629_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2296),
    .D(_00319_),
    .Q_N(_00051_),
    .Q(\soc_I.clint_I.mtimecmp[53] ));
 sg13g2_dfrbp_1 _33630_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2294),
    .D(_00320_),
    .Q_N(_00059_),
    .Q(\soc_I.clint_I.mtimecmp[54] ));
 sg13g2_dfrbp_1 _33631_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2292),
    .D(_00321_),
    .Q_N(_00067_),
    .Q(\soc_I.clint_I.mtimecmp[55] ));
 sg13g2_dfrbp_1 _33632_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2290),
    .D(_00322_),
    .Q_N(_00017_),
    .Q(\soc_I.clint_I.mtimecmp[56] ));
 sg13g2_dfrbp_1 _33633_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2288),
    .D(_00323_),
    .Q_N(_00025_),
    .Q(\soc_I.clint_I.mtimecmp[57] ));
 sg13g2_dfrbp_1 _33634_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net2286),
    .D(_00324_),
    .Q_N(_00033_),
    .Q(\soc_I.clint_I.mtimecmp[58] ));
 sg13g2_dfrbp_1 _33635_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2284),
    .D(_00325_),
    .Q_N(_00041_),
    .Q(\soc_I.clint_I.mtimecmp[59] ));
 sg13g2_dfrbp_1 _33636_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net2282),
    .D(_00326_),
    .Q_N(_00047_),
    .Q(\soc_I.clint_I.mtimecmp[60] ));
 sg13g2_dfrbp_1 _33637_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2280),
    .D(_00327_),
    .Q_N(_00055_),
    .Q(\soc_I.clint_I.mtimecmp[61] ));
 sg13g2_dfrbp_1 _33638_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2278),
    .D(_00328_),
    .Q_N(_00063_),
    .Q(\soc_I.clint_I.mtimecmp[62] ));
 sg13g2_dfrbp_1 _33639_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net2276),
    .D(_00329_),
    .Q_N(_00072_),
    .Q(\soc_I.clint_I.mtimecmp[63] ));
 sg13g2_dfrbp_1 _33640_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net2274),
    .D(_00330_),
    .Q_N(_16654_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[4][0] ));
 sg13g2_dfrbp_1 _33641_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net2273),
    .D(net4137),
    .Q_N(_16653_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[4][1] ));
 sg13g2_dfrbp_1 _33642_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net2272),
    .D(net3942),
    .Q_N(_16652_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[4][2] ));
 sg13g2_dfrbp_1 _33643_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net2271),
    .D(net4075),
    .Q_N(_16651_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[4][3] ));
 sg13g2_dfrbp_1 _33644_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net2270),
    .D(net4083),
    .Q_N(_16650_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[4][4] ));
 sg13g2_dfrbp_1 _33645_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net2269),
    .D(net3922),
    .Q_N(_16649_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[4][5] ));
 sg13g2_dfrbp_1 _33646_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net2268),
    .D(_00336_),
    .Q_N(_16648_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[4][6] ));
 sg13g2_dfrbp_1 _33647_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net2267),
    .D(net4183),
    .Q_N(_16647_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[4][7] ));
 sg13g2_dfrbp_1 _33648_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2266),
    .D(_00338_),
    .Q_N(_16646_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][0] ));
 sg13g2_dfrbp_1 _33649_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2265),
    .D(_00339_),
    .Q_N(_16645_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][1] ));
 sg13g2_dfrbp_1 _33650_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2264),
    .D(_00340_),
    .Q_N(_16644_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][2] ));
 sg13g2_dfrbp_1 _33651_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2263),
    .D(_00341_),
    .Q_N(_16643_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][3] ));
 sg13g2_dfrbp_1 _33652_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2262),
    .D(_00342_),
    .Q_N(_16642_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][4] ));
 sg13g2_dfrbp_1 _33653_ (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2261),
    .D(_00343_),
    .Q_N(_16641_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][5] ));
 sg13g2_dfrbp_1 _33654_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2260),
    .D(_00344_),
    .Q_N(_16640_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][6] ));
 sg13g2_dfrbp_1 _33655_ (.CLK(clknet_leaf_322_clk),
    .RESET_B(net2259),
    .D(_00345_),
    .Q_N(_16639_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][7] ));
 sg13g2_dfrbp_1 _33656_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2258),
    .D(_00346_),
    .Q_N(_16638_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][8] ));
 sg13g2_dfrbp_1 _33657_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2257),
    .D(_00347_),
    .Q_N(_16637_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][9] ));
 sg13g2_dfrbp_1 _33658_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2256),
    .D(_00348_),
    .Q_N(_16636_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][10] ));
 sg13g2_dfrbp_1 _33659_ (.CLK(clknet_leaf_319_clk),
    .RESET_B(net2255),
    .D(_00349_),
    .Q_N(_16635_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][11] ));
 sg13g2_dfrbp_1 _33660_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2254),
    .D(_00350_),
    .Q_N(_16634_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][12] ));
 sg13g2_dfrbp_1 _33661_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2253),
    .D(_00351_),
    .Q_N(_16633_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][13] ));
 sg13g2_dfrbp_1 _33662_ (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2252),
    .D(_00352_),
    .Q_N(_16632_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][14] ));
 sg13g2_dfrbp_1 _33663_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2251),
    .D(_00353_),
    .Q_N(_16631_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][15] ));
 sg13g2_dfrbp_1 _33664_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net2250),
    .D(_00354_),
    .Q_N(_16630_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][16] ));
 sg13g2_dfrbp_1 _33665_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net2249),
    .D(_00355_),
    .Q_N(_16629_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][17] ));
 sg13g2_dfrbp_1 _33666_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net2248),
    .D(_00356_),
    .Q_N(_16628_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][18] ));
 sg13g2_dfrbp_1 _33667_ (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2247),
    .D(_00357_),
    .Q_N(_16627_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][19] ));
 sg13g2_dfrbp_1 _33668_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2246),
    .D(_00358_),
    .Q_N(_16626_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][20] ));
 sg13g2_dfrbp_1 _33669_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2245),
    .D(_00359_),
    .Q_N(_16625_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][21] ));
 sg13g2_dfrbp_1 _33670_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2244),
    .D(_00360_),
    .Q_N(_16624_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][22] ));
 sg13g2_dfrbp_1 _33671_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2243),
    .D(_00361_),
    .Q_N(_16623_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][23] ));
 sg13g2_dfrbp_1 _33672_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2242),
    .D(_00362_),
    .Q_N(_16622_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][24] ));
 sg13g2_dfrbp_1 _33673_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2241),
    .D(_00363_),
    .Q_N(_16621_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][25] ));
 sg13g2_dfrbp_1 _33674_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2240),
    .D(_00364_),
    .Q_N(_16620_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][26] ));
 sg13g2_dfrbp_1 _33675_ (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2239),
    .D(_00365_),
    .Q_N(_16619_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][27] ));
 sg13g2_dfrbp_1 _33676_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2238),
    .D(_00366_),
    .Q_N(_16618_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][28] ));
 sg13g2_dfrbp_1 _33677_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2237),
    .D(_00367_),
    .Q_N(_16617_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][29] ));
 sg13g2_dfrbp_1 _33678_ (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2236),
    .D(_00368_),
    .Q_N(_16616_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][30] ));
 sg13g2_dfrbp_1 _33679_ (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2235),
    .D(_00369_),
    .Q_N(_16615_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][31] ));
 sg13g2_dfrbp_1 _33680_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2234),
    .D(_00370_),
    .Q_N(_16614_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][0] ));
 sg13g2_dfrbp_1 _33681_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2233),
    .D(_00371_),
    .Q_N(_16613_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][1] ));
 sg13g2_dfrbp_1 _33682_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2232),
    .D(_00372_),
    .Q_N(_16612_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][2] ));
 sg13g2_dfrbp_1 _33683_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2231),
    .D(_00373_),
    .Q_N(_16611_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][3] ));
 sg13g2_dfrbp_1 _33684_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2230),
    .D(_00374_),
    .Q_N(_16610_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][4] ));
 sg13g2_dfrbp_1 _33685_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2229),
    .D(_00375_),
    .Q_N(_16609_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][5] ));
 sg13g2_dfrbp_1 _33686_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2228),
    .D(_00376_),
    .Q_N(_16608_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][6] ));
 sg13g2_dfrbp_1 _33687_ (.CLK(clknet_leaf_318_clk),
    .RESET_B(net2227),
    .D(_00377_),
    .Q_N(_16607_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][7] ));
 sg13g2_dfrbp_1 _33688_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2226),
    .D(_00378_),
    .Q_N(_16606_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][8] ));
 sg13g2_dfrbp_1 _33689_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2225),
    .D(_00379_),
    .Q_N(_16605_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][9] ));
 sg13g2_dfrbp_1 _33690_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2224),
    .D(_00380_),
    .Q_N(_16604_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][10] ));
 sg13g2_dfrbp_1 _33691_ (.CLK(clknet_leaf_318_clk),
    .RESET_B(net2223),
    .D(_00381_),
    .Q_N(_16603_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][11] ));
 sg13g2_dfrbp_1 _33692_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2222),
    .D(_00382_),
    .Q_N(_16602_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][12] ));
 sg13g2_dfrbp_1 _33693_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2221),
    .D(_00383_),
    .Q_N(_16601_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][13] ));
 sg13g2_dfrbp_1 _33694_ (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2220),
    .D(_00384_),
    .Q_N(_16600_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][14] ));
 sg13g2_dfrbp_1 _33695_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net2219),
    .D(_00385_),
    .Q_N(_16599_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][15] ));
 sg13g2_dfrbp_1 _33696_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net2218),
    .D(_00386_),
    .Q_N(_16598_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][16] ));
 sg13g2_dfrbp_1 _33697_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net2217),
    .D(_00387_),
    .Q_N(_16597_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][17] ));
 sg13g2_dfrbp_1 _33698_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net2216),
    .D(_00388_),
    .Q_N(_16596_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][18] ));
 sg13g2_dfrbp_1 _33699_ (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2215),
    .D(_00389_),
    .Q_N(_16595_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][19] ));
 sg13g2_dfrbp_1 _33700_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2214),
    .D(_00390_),
    .Q_N(_16594_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][20] ));
 sg13g2_dfrbp_1 _33701_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2213),
    .D(_00391_),
    .Q_N(_16593_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][21] ));
 sg13g2_dfrbp_1 _33702_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2212),
    .D(_00392_),
    .Q_N(_16592_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][22] ));
 sg13g2_dfrbp_1 _33703_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net2211),
    .D(_00393_),
    .Q_N(_16591_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][23] ));
 sg13g2_dfrbp_1 _33704_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2210),
    .D(_00394_),
    .Q_N(_16590_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][24] ));
 sg13g2_dfrbp_1 _33705_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2209),
    .D(_00395_),
    .Q_N(_16589_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][25] ));
 sg13g2_dfrbp_1 _33706_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2208),
    .D(_00396_),
    .Q_N(_16588_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][26] ));
 sg13g2_dfrbp_1 _33707_ (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2207),
    .D(_00397_),
    .Q_N(_16587_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][27] ));
 sg13g2_dfrbp_1 _33708_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2206),
    .D(_00398_),
    .Q_N(_16586_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][28] ));
 sg13g2_dfrbp_1 _33709_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2205),
    .D(_00399_),
    .Q_N(_16585_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][29] ));
 sg13g2_dfrbp_1 _33710_ (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2204),
    .D(_00400_),
    .Q_N(_16584_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][30] ));
 sg13g2_dfrbp_1 _33711_ (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2203),
    .D(_00401_),
    .Q_N(_16583_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][31] ));
 sg13g2_dfrbp_1 _33712_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2202),
    .D(_00402_),
    .Q_N(_16582_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][0] ));
 sg13g2_dfrbp_1 _33713_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2201),
    .D(_00403_),
    .Q_N(_16581_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][1] ));
 sg13g2_dfrbp_1 _33714_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2200),
    .D(_00404_),
    .Q_N(_16580_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][2] ));
 sg13g2_dfrbp_1 _33715_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2199),
    .D(_00405_),
    .Q_N(_16579_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][3] ));
 sg13g2_dfrbp_1 _33716_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2198),
    .D(_00406_),
    .Q_N(_16578_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][4] ));
 sg13g2_dfrbp_1 _33717_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2197),
    .D(_00407_),
    .Q_N(_16577_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][5] ));
 sg13g2_dfrbp_1 _33718_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2196),
    .D(_00408_),
    .Q_N(_16576_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][6] ));
 sg13g2_dfrbp_1 _33719_ (.CLK(clknet_leaf_319_clk),
    .RESET_B(net2195),
    .D(_00409_),
    .Q_N(_16575_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][7] ));
 sg13g2_dfrbp_1 _33720_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2194),
    .D(_00410_),
    .Q_N(_16574_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][8] ));
 sg13g2_dfrbp_1 _33721_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2193),
    .D(_00411_),
    .Q_N(_16573_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][9] ));
 sg13g2_dfrbp_1 _33722_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2192),
    .D(_00412_),
    .Q_N(_16572_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][10] ));
 sg13g2_dfrbp_1 _33723_ (.CLK(clknet_leaf_319_clk),
    .RESET_B(net2191),
    .D(_00413_),
    .Q_N(_16571_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][11] ));
 sg13g2_dfrbp_1 _33724_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2190),
    .D(_00414_),
    .Q_N(_16570_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][12] ));
 sg13g2_dfrbp_1 _33725_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2189),
    .D(_00415_),
    .Q_N(_16569_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][13] ));
 sg13g2_dfrbp_1 _33726_ (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2188),
    .D(_00416_),
    .Q_N(_16568_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][14] ));
 sg13g2_dfrbp_1 _33727_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net2187),
    .D(_00417_),
    .Q_N(_16567_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][15] ));
 sg13g2_dfrbp_1 _33728_ (.CLK(clknet_leaf_313_clk),
    .RESET_B(net2186),
    .D(_00418_),
    .Q_N(_16566_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][16] ));
 sg13g2_dfrbp_1 _33729_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net2185),
    .D(_00419_),
    .Q_N(_16565_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][17] ));
 sg13g2_dfrbp_1 _33730_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net2184),
    .D(_00420_),
    .Q_N(_16564_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][18] ));
 sg13g2_dfrbp_1 _33731_ (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2183),
    .D(_00421_),
    .Q_N(_16563_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][19] ));
 sg13g2_dfrbp_1 _33732_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2182),
    .D(_00422_),
    .Q_N(_16562_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][20] ));
 sg13g2_dfrbp_1 _33733_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net2181),
    .D(_00423_),
    .Q_N(_16561_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][21] ));
 sg13g2_dfrbp_1 _33734_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2180),
    .D(_00424_),
    .Q_N(_16560_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][22] ));
 sg13g2_dfrbp_1 _33735_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net2179),
    .D(_00425_),
    .Q_N(_16559_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][23] ));
 sg13g2_dfrbp_1 _33736_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2178),
    .D(_00426_),
    .Q_N(_16558_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][24] ));
 sg13g2_dfrbp_1 _33737_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2177),
    .D(_00427_),
    .Q_N(_16557_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][25] ));
 sg13g2_dfrbp_1 _33738_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2176),
    .D(_00428_),
    .Q_N(_16556_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][26] ));
 sg13g2_dfrbp_1 _33739_ (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2175),
    .D(_00429_),
    .Q_N(_16555_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][27] ));
 sg13g2_dfrbp_1 _33740_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net2174),
    .D(_00430_),
    .Q_N(_16554_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][28] ));
 sg13g2_dfrbp_1 _33741_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2173),
    .D(_00431_),
    .Q_N(_16553_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][29] ));
 sg13g2_dfrbp_1 _33742_ (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2172),
    .D(_00432_),
    .Q_N(_16552_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][30] ));
 sg13g2_dfrbp_1 _33743_ (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2171),
    .D(_00433_),
    .Q_N(_16551_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][31] ));
 sg13g2_dfrbp_1 _33744_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2170),
    .D(_00434_),
    .Q_N(_16550_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][0] ));
 sg13g2_dfrbp_1 _33745_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2169),
    .D(_00435_),
    .Q_N(_16549_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][1] ));
 sg13g2_dfrbp_1 _33746_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2168),
    .D(_00436_),
    .Q_N(_16548_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][2] ));
 sg13g2_dfrbp_1 _33747_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2167),
    .D(_00437_),
    .Q_N(_16547_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][3] ));
 sg13g2_dfrbp_1 _33748_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2166),
    .D(_00438_),
    .Q_N(_16546_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][4] ));
 sg13g2_dfrbp_1 _33749_ (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2165),
    .D(_00439_),
    .Q_N(_16545_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][5] ));
 sg13g2_dfrbp_1 _33750_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2164),
    .D(_00440_),
    .Q_N(_16544_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][6] ));
 sg13g2_dfrbp_1 _33751_ (.CLK(clknet_leaf_320_clk),
    .RESET_B(net2163),
    .D(_00441_),
    .Q_N(_16543_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][7] ));
 sg13g2_dfrbp_1 _33752_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2162),
    .D(_00442_),
    .Q_N(_16542_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][8] ));
 sg13g2_dfrbp_1 _33753_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2161),
    .D(_00443_),
    .Q_N(_16541_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][9] ));
 sg13g2_dfrbp_1 _33754_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2160),
    .D(_00444_),
    .Q_N(_16540_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][10] ));
 sg13g2_dfrbp_1 _33755_ (.CLK(clknet_leaf_320_clk),
    .RESET_B(net2159),
    .D(_00445_),
    .Q_N(_16539_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][11] ));
 sg13g2_dfrbp_1 _33756_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2158),
    .D(_00446_),
    .Q_N(_16538_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][12] ));
 sg13g2_dfrbp_1 _33757_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2157),
    .D(_00447_),
    .Q_N(_16537_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][13] ));
 sg13g2_dfrbp_1 _33758_ (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2156),
    .D(_00448_),
    .Q_N(_16536_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][14] ));
 sg13g2_dfrbp_1 _33759_ (.CLK(clknet_leaf_311_clk),
    .RESET_B(net2155),
    .D(_00449_),
    .Q_N(_16535_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][15] ));
 sg13g2_dfrbp_1 _33760_ (.CLK(clknet_leaf_320_clk),
    .RESET_B(net2154),
    .D(_00450_),
    .Q_N(_16534_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][16] ));
 sg13g2_dfrbp_1 _33761_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net2153),
    .D(_00451_),
    .Q_N(_16533_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][17] ));
 sg13g2_dfrbp_1 _33762_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net2152),
    .D(_00452_),
    .Q_N(_16532_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][18] ));
 sg13g2_dfrbp_1 _33763_ (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2151),
    .D(_00453_),
    .Q_N(_16531_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][19] ));
 sg13g2_dfrbp_1 _33764_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2150),
    .D(_00454_),
    .Q_N(_16530_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][20] ));
 sg13g2_dfrbp_1 _33765_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2149),
    .D(_00455_),
    .Q_N(_16529_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][21] ));
 sg13g2_dfrbp_1 _33766_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2148),
    .D(_00456_),
    .Q_N(_16528_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][22] ));
 sg13g2_dfrbp_1 _33767_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2147),
    .D(_00457_),
    .Q_N(_16527_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][23] ));
 sg13g2_dfrbp_1 _33768_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2146),
    .D(_00458_),
    .Q_N(_16526_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][24] ));
 sg13g2_dfrbp_1 _33769_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2145),
    .D(_00459_),
    .Q_N(_16525_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][25] ));
 sg13g2_dfrbp_1 _33770_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2144),
    .D(_00460_),
    .Q_N(_16524_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][26] ));
 sg13g2_dfrbp_1 _33771_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net2143),
    .D(_00461_),
    .Q_N(_16523_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][27] ));
 sg13g2_dfrbp_1 _33772_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net2142),
    .D(_00462_),
    .Q_N(_16522_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][28] ));
 sg13g2_dfrbp_1 _33773_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net2141),
    .D(_00463_),
    .Q_N(_16521_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][29] ));
 sg13g2_dfrbp_1 _33774_ (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2140),
    .D(_00464_),
    .Q_N(_16520_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][30] ));
 sg13g2_dfrbp_1 _33775_ (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2139),
    .D(_00465_),
    .Q_N(_16519_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][31] ));
 sg13g2_dfrbp_1 _33776_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net2138),
    .D(net4857),
    .Q_N(_00151_),
    .Q(\soc_I.qqspi_I.xfer_cycles[2] ));
 sg13g2_dfrbp_1 _33777_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net2136),
    .D(_00467_),
    .Q_N(_16518_),
    .Q(\soc_I.qqspi_I.xfer_cycles[3] ));
 sg13g2_dfrbp_1 _33778_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net2134),
    .D(net5051),
    .Q_N(_16517_),
    .Q(\soc_I.qqspi_I.xfer_cycles[4] ));
 sg13g2_dfrbp_1 _33779_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net2132),
    .D(net5105),
    .Q_N(_16516_),
    .Q(\soc_I.qqspi_I.xfer_cycles[5] ));
 sg13g2_dfrbp_1 _33780_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2130),
    .D(_00470_),
    .Q_N(_16515_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][0] ));
 sg13g2_dfrbp_1 _33781_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2129),
    .D(_00471_),
    .Q_N(_16514_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][1] ));
 sg13g2_dfrbp_1 _33782_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2128),
    .D(_00472_),
    .Q_N(_16513_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][2] ));
 sg13g2_dfrbp_1 _33783_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2127),
    .D(_00473_),
    .Q_N(_16512_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][3] ));
 sg13g2_dfrbp_1 _33784_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2126),
    .D(_00474_),
    .Q_N(_16511_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][4] ));
 sg13g2_dfrbp_1 _33785_ (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2125),
    .D(_00475_),
    .Q_N(_16510_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][5] ));
 sg13g2_dfrbp_1 _33786_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2124),
    .D(_00476_),
    .Q_N(_16509_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][6] ));
 sg13g2_dfrbp_1 _33787_ (.CLK(clknet_leaf_312_clk),
    .RESET_B(net2123),
    .D(_00477_),
    .Q_N(_16508_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][7] ));
 sg13g2_dfrbp_1 _33788_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2122),
    .D(_00478_),
    .Q_N(_16507_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][8] ));
 sg13g2_dfrbp_1 _33789_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2121),
    .D(_00479_),
    .Q_N(_16506_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][9] ));
 sg13g2_dfrbp_1 _33790_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2120),
    .D(_00480_),
    .Q_N(_16505_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][10] ));
 sg13g2_dfrbp_1 _33791_ (.CLK(clknet_leaf_313_clk),
    .RESET_B(net2119),
    .D(_00481_),
    .Q_N(_16504_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][11] ));
 sg13g2_dfrbp_1 _33792_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2118),
    .D(_00482_),
    .Q_N(_16503_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][12] ));
 sg13g2_dfrbp_1 _33793_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2117),
    .D(_00483_),
    .Q_N(_16502_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][13] ));
 sg13g2_dfrbp_1 _33794_ (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2116),
    .D(_00484_),
    .Q_N(_16501_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][14] ));
 sg13g2_dfrbp_1 _33795_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net2115),
    .D(_00485_),
    .Q_N(_16500_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][15] ));
 sg13g2_dfrbp_1 _33796_ (.CLK(clknet_leaf_313_clk),
    .RESET_B(net2114),
    .D(_00486_),
    .Q_N(_16499_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][16] ));
 sg13g2_dfrbp_1 _33797_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net2113),
    .D(_00487_),
    .Q_N(_16498_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][17] ));
 sg13g2_dfrbp_1 _33798_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net2112),
    .D(_00488_),
    .Q_N(_16497_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][18] ));
 sg13g2_dfrbp_1 _33799_ (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2111),
    .D(_00489_),
    .Q_N(_16496_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][19] ));
 sg13g2_dfrbp_1 _33800_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2110),
    .D(_00490_),
    .Q_N(_16495_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][20] ));
 sg13g2_dfrbp_1 _33801_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2109),
    .D(_00491_),
    .Q_N(_16494_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][21] ));
 sg13g2_dfrbp_1 _33802_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2108),
    .D(_00492_),
    .Q_N(_16493_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][22] ));
 sg13g2_dfrbp_1 _33803_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2107),
    .D(_00493_),
    .Q_N(_16492_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][23] ));
 sg13g2_dfrbp_1 _33804_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2106),
    .D(_00494_),
    .Q_N(_16491_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][24] ));
 sg13g2_dfrbp_1 _33805_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2105),
    .D(_00495_),
    .Q_N(_16490_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][25] ));
 sg13g2_dfrbp_1 _33806_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2104),
    .D(_00496_),
    .Q_N(_16489_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][26] ));
 sg13g2_dfrbp_1 _33807_ (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2103),
    .D(_00497_),
    .Q_N(_16488_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][27] ));
 sg13g2_dfrbp_1 _33808_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2102),
    .D(_00498_),
    .Q_N(_16487_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][28] ));
 sg13g2_dfrbp_1 _33809_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net2101),
    .D(_00499_),
    .Q_N(_16486_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][29] ));
 sg13g2_dfrbp_1 _33810_ (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2100),
    .D(_00500_),
    .Q_N(_16485_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][30] ));
 sg13g2_dfrbp_1 _33811_ (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2099),
    .D(_00501_),
    .Q_N(_16484_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][31] ));
 sg13g2_dfrbp_1 _33812_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2098),
    .D(_00502_),
    .Q_N(_16483_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][0] ));
 sg13g2_dfrbp_1 _33813_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2097),
    .D(_00503_),
    .Q_N(_16482_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][1] ));
 sg13g2_dfrbp_1 _33814_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2096),
    .D(_00504_),
    .Q_N(_16481_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][2] ));
 sg13g2_dfrbp_1 _33815_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2095),
    .D(_00505_),
    .Q_N(_16480_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][3] ));
 sg13g2_dfrbp_1 _33816_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2094),
    .D(_00506_),
    .Q_N(_16479_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][4] ));
 sg13g2_dfrbp_1 _33817_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2093),
    .D(_00507_),
    .Q_N(_16478_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][5] ));
 sg13g2_dfrbp_1 _33818_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2092),
    .D(_00508_),
    .Q_N(_16477_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][6] ));
 sg13g2_dfrbp_1 _33819_ (.CLK(clknet_leaf_320_clk),
    .RESET_B(net2091),
    .D(_00509_),
    .Q_N(_16476_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][7] ));
 sg13g2_dfrbp_1 _33820_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2090),
    .D(_00510_),
    .Q_N(_16475_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][8] ));
 sg13g2_dfrbp_1 _33821_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2089),
    .D(_00511_),
    .Q_N(_16474_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][9] ));
 sg13g2_dfrbp_1 _33822_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2088),
    .D(_00512_),
    .Q_N(_16473_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][10] ));
 sg13g2_dfrbp_1 _33823_ (.CLK(clknet_leaf_313_clk),
    .RESET_B(net2087),
    .D(_00513_),
    .Q_N(_16472_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][11] ));
 sg13g2_dfrbp_1 _33824_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2086),
    .D(_00514_),
    .Q_N(_16471_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][12] ));
 sg13g2_dfrbp_1 _33825_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2085),
    .D(_00515_),
    .Q_N(_16470_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][13] ));
 sg13g2_dfrbp_1 _33826_ (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2084),
    .D(_00516_),
    .Q_N(_16469_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][14] ));
 sg13g2_dfrbp_1 _33827_ (.CLK(clknet_leaf_311_clk),
    .RESET_B(net2083),
    .D(_00517_),
    .Q_N(_16468_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][15] ));
 sg13g2_dfrbp_1 _33828_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net2082),
    .D(_00518_),
    .Q_N(_16467_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][16] ));
 sg13g2_dfrbp_1 _33829_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net2081),
    .D(_00519_),
    .Q_N(_16466_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][17] ));
 sg13g2_dfrbp_1 _33830_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net2080),
    .D(_00520_),
    .Q_N(_16465_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][18] ));
 sg13g2_dfrbp_1 _33831_ (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2079),
    .D(_00521_),
    .Q_N(_16464_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][19] ));
 sg13g2_dfrbp_1 _33832_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2078),
    .D(_00522_),
    .Q_N(_16463_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][20] ));
 sg13g2_dfrbp_1 _33833_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2077),
    .D(_00523_),
    .Q_N(_16462_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][21] ));
 sg13g2_dfrbp_1 _33834_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2076),
    .D(_00524_),
    .Q_N(_16461_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][22] ));
 sg13g2_dfrbp_1 _33835_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2075),
    .D(_00525_),
    .Q_N(_16460_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][23] ));
 sg13g2_dfrbp_1 _33836_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2074),
    .D(_00526_),
    .Q_N(_16459_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][24] ));
 sg13g2_dfrbp_1 _33837_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2073),
    .D(_00527_),
    .Q_N(_16458_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][25] ));
 sg13g2_dfrbp_1 _33838_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2072),
    .D(_00528_),
    .Q_N(_16457_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][26] ));
 sg13g2_dfrbp_1 _33839_ (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2071),
    .D(_00529_),
    .Q_N(_16456_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][27] ));
 sg13g2_dfrbp_1 _33840_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2070),
    .D(_00530_),
    .Q_N(_16455_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][28] ));
 sg13g2_dfrbp_1 _33841_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2069),
    .D(_00531_),
    .Q_N(_16454_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][29] ));
 sg13g2_dfrbp_1 _33842_ (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2068),
    .D(_00532_),
    .Q_N(_16453_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][30] ));
 sg13g2_dfrbp_1 _33843_ (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2067),
    .D(_00533_),
    .Q_N(_16452_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][31] ));
 sg13g2_dfrbp_1 _33844_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2066),
    .D(_00534_),
    .Q_N(_16451_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][0] ));
 sg13g2_dfrbp_1 _33845_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2065),
    .D(_00535_),
    .Q_N(_16450_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][1] ));
 sg13g2_dfrbp_1 _33846_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2064),
    .D(_00536_),
    .Q_N(_16449_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][2] ));
 sg13g2_dfrbp_1 _33847_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2063),
    .D(_00537_),
    .Q_N(_16448_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][3] ));
 sg13g2_dfrbp_1 _33848_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2062),
    .D(_00538_),
    .Q_N(_16447_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][4] ));
 sg13g2_dfrbp_1 _33849_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2061),
    .D(_00539_),
    .Q_N(_16446_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][5] ));
 sg13g2_dfrbp_1 _33850_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2060),
    .D(_00540_),
    .Q_N(_16445_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][6] ));
 sg13g2_dfrbp_1 _33851_ (.CLK(clknet_leaf_307_clk),
    .RESET_B(net2059),
    .D(_00541_),
    .Q_N(_16444_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][7] ));
 sg13g2_dfrbp_1 _33852_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2058),
    .D(_00542_),
    .Q_N(_16443_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][8] ));
 sg13g2_dfrbp_1 _33853_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2057),
    .D(_00543_),
    .Q_N(_16442_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][9] ));
 sg13g2_dfrbp_1 _33854_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2056),
    .D(_00544_),
    .Q_N(_16441_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][10] ));
 sg13g2_dfrbp_1 _33855_ (.CLK(clknet_leaf_315_clk),
    .RESET_B(net2055),
    .D(_00545_),
    .Q_N(_16440_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][11] ));
 sg13g2_dfrbp_1 _33856_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2054),
    .D(_00546_),
    .Q_N(_16439_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][12] ));
 sg13g2_dfrbp_1 _33857_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2053),
    .D(_00547_),
    .Q_N(_16438_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][13] ));
 sg13g2_dfrbp_1 _33858_ (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2052),
    .D(_00548_),
    .Q_N(_16437_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][14] ));
 sg13g2_dfrbp_1 _33859_ (.CLK(clknet_leaf_310_clk),
    .RESET_B(net2051),
    .D(_00549_),
    .Q_N(_16436_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][15] ));
 sg13g2_dfrbp_1 _33860_ (.CLK(clknet_leaf_315_clk),
    .RESET_B(net2050),
    .D(_00550_),
    .Q_N(_16435_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][16] ));
 sg13g2_dfrbp_1 _33861_ (.CLK(clknet_leaf_312_clk),
    .RESET_B(net2049),
    .D(_00551_),
    .Q_N(_16434_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][17] ));
 sg13g2_dfrbp_1 _33862_ (.CLK(clknet_leaf_302_clk),
    .RESET_B(net2048),
    .D(_00552_),
    .Q_N(_16433_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][18] ));
 sg13g2_dfrbp_1 _33863_ (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2047),
    .D(_00553_),
    .Q_N(_16432_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][19] ));
 sg13g2_dfrbp_1 _33864_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2046),
    .D(_00554_),
    .Q_N(_16431_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][20] ));
 sg13g2_dfrbp_1 _33865_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2045),
    .D(_00555_),
    .Q_N(_16430_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][21] ));
 sg13g2_dfrbp_1 _33866_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2044),
    .D(_00556_),
    .Q_N(_16429_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][22] ));
 sg13g2_dfrbp_1 _33867_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2043),
    .D(_00557_),
    .Q_N(_16428_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][23] ));
 sg13g2_dfrbp_1 _33868_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2042),
    .D(_00558_),
    .Q_N(_16427_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][24] ));
 sg13g2_dfrbp_1 _33869_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2041),
    .D(_00559_),
    .Q_N(_16426_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][25] ));
 sg13g2_dfrbp_1 _33870_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2040),
    .D(_00560_),
    .Q_N(_16425_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][26] ));
 sg13g2_dfrbp_1 _33871_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2039),
    .D(_00561_),
    .Q_N(_16424_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][27] ));
 sg13g2_dfrbp_1 _33872_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2038),
    .D(_00562_),
    .Q_N(_16423_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][28] ));
 sg13g2_dfrbp_1 _33873_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2037),
    .D(_00563_),
    .Q_N(_16422_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][29] ));
 sg13g2_dfrbp_1 _33874_ (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2036),
    .D(_00564_),
    .Q_N(_16421_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][30] ));
 sg13g2_dfrbp_1 _33875_ (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2035),
    .D(_00565_),
    .Q_N(_16420_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][31] ));
 sg13g2_dfrbp_1 _33876_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2034),
    .D(_00566_),
    .Q_N(_16419_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][0] ));
 sg13g2_dfrbp_1 _33877_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2033),
    .D(_00567_),
    .Q_N(_16418_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][1] ));
 sg13g2_dfrbp_1 _33878_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2032),
    .D(_00568_),
    .Q_N(_16417_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][2] ));
 sg13g2_dfrbp_1 _33879_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2031),
    .D(_00569_),
    .Q_N(_16416_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][3] ));
 sg13g2_dfrbp_1 _33880_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2030),
    .D(_00570_),
    .Q_N(_16415_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][4] ));
 sg13g2_dfrbp_1 _33881_ (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2029),
    .D(_00571_),
    .Q_N(_16414_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][5] ));
 sg13g2_dfrbp_1 _33882_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2028),
    .D(_00572_),
    .Q_N(_16413_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][6] ));
 sg13g2_dfrbp_1 _33883_ (.CLK(clknet_leaf_322_clk),
    .RESET_B(net2027),
    .D(_00573_),
    .Q_N(_16412_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][7] ));
 sg13g2_dfrbp_1 _33884_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2026),
    .D(_00574_),
    .Q_N(_16411_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][8] ));
 sg13g2_dfrbp_1 _33885_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2025),
    .D(_00575_),
    .Q_N(_16410_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][9] ));
 sg13g2_dfrbp_1 _33886_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2024),
    .D(_00576_),
    .Q_N(_16409_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][10] ));
 sg13g2_dfrbp_1 _33887_ (.CLK(clknet_leaf_323_clk),
    .RESET_B(net2023),
    .D(_00577_),
    .Q_N(_16408_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][11] ));
 sg13g2_dfrbp_1 _33888_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2022),
    .D(_00578_),
    .Q_N(_16407_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][12] ));
 sg13g2_dfrbp_1 _33889_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2021),
    .D(_00579_),
    .Q_N(_16406_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][13] ));
 sg13g2_dfrbp_1 _33890_ (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2020),
    .D(_00580_),
    .Q_N(_16405_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][14] ));
 sg13g2_dfrbp_1 _33891_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2019),
    .D(_00581_),
    .Q_N(_16404_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][15] ));
 sg13g2_dfrbp_1 _33892_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net2018),
    .D(_00582_),
    .Q_N(_16403_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][16] ));
 sg13g2_dfrbp_1 _33893_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net2017),
    .D(_00583_),
    .Q_N(_16402_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][17] ));
 sg13g2_dfrbp_1 _33894_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net2016),
    .D(_00584_),
    .Q_N(_16401_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][18] ));
 sg13g2_dfrbp_1 _33895_ (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2015),
    .D(_00585_),
    .Q_N(_16400_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][19] ));
 sg13g2_dfrbp_1 _33896_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2014),
    .D(_00586_),
    .Q_N(_16399_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][20] ));
 sg13g2_dfrbp_1 _33897_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2013),
    .D(_00587_),
    .Q_N(_16398_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][21] ));
 sg13g2_dfrbp_1 _33898_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2012),
    .D(_00588_),
    .Q_N(_16397_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][22] ));
 sg13g2_dfrbp_1 _33899_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2011),
    .D(_00589_),
    .Q_N(_16396_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][23] ));
 sg13g2_dfrbp_1 _33900_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2010),
    .D(_00590_),
    .Q_N(_16395_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][24] ));
 sg13g2_dfrbp_1 _33901_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2009),
    .D(_00591_),
    .Q_N(_16394_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][25] ));
 sg13g2_dfrbp_1 _33902_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2008),
    .D(_00592_),
    .Q_N(_16393_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][26] ));
 sg13g2_dfrbp_1 _33903_ (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2007),
    .D(_00593_),
    .Q_N(_16392_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][27] ));
 sg13g2_dfrbp_1 _33904_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2006),
    .D(_00594_),
    .Q_N(_16391_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][28] ));
 sg13g2_dfrbp_1 _33905_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2005),
    .D(_00595_),
    .Q_N(_16390_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][29] ));
 sg13g2_dfrbp_1 _33906_ (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2004),
    .D(_00596_),
    .Q_N(_16389_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][30] ));
 sg13g2_dfrbp_1 _33907_ (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2003),
    .D(_00597_),
    .Q_N(_16388_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][31] ));
 sg13g2_dfrbp_1 _33908_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2002),
    .D(_00598_),
    .Q_N(_00110_),
    .Q(\soc_I.clint_I.mtimecmp[0] ));
 sg13g2_dfrbp_1 _33909_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net2000),
    .D(_00599_),
    .Q_N(_00115_),
    .Q(\soc_I.clint_I.mtimecmp[1] ));
 sg13g2_dfrbp_1 _33910_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1998),
    .D(_00600_),
    .Q_N(_00120_),
    .Q(\soc_I.clint_I.mtimecmp[2] ));
 sg13g2_dfrbp_1 _33911_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1996),
    .D(_00601_),
    .Q_N(_00125_),
    .Q(\soc_I.clint_I.mtimecmp[3] ));
 sg13g2_dfrbp_1 _33912_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1994),
    .D(_00602_),
    .Q_N(_00130_),
    .Q(\soc_I.clint_I.mtimecmp[4] ));
 sg13g2_dfrbp_1 _33913_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1992),
    .D(_00603_),
    .Q_N(_00135_),
    .Q(\soc_I.clint_I.mtimecmp[5] ));
 sg13g2_dfrbp_1 _33914_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1990),
    .D(_00604_),
    .Q_N(_00140_),
    .Q(\soc_I.clint_I.mtimecmp[6] ));
 sg13g2_dfrbp_1 _33915_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1988),
    .D(_00605_),
    .Q_N(_00145_),
    .Q(\soc_I.clint_I.mtimecmp[7] ));
 sg13g2_dfrbp_1 _33916_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1986),
    .D(_00606_),
    .Q_N(_00075_),
    .Q(\soc_I.clint_I.mtimecmp[8] ));
 sg13g2_dfrbp_1 _33917_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1984),
    .D(_00607_),
    .Q_N(_00079_),
    .Q(\soc_I.clint_I.mtimecmp[9] ));
 sg13g2_dfrbp_1 _33918_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1982),
    .D(_00608_),
    .Q_N(_00083_),
    .Q(\soc_I.clint_I.mtimecmp[10] ));
 sg13g2_dfrbp_1 _33919_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1980),
    .D(_00609_),
    .Q_N(_00087_),
    .Q(\soc_I.clint_I.mtimecmp[11] ));
 sg13g2_dfrbp_1 _33920_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1978),
    .D(_00610_),
    .Q_N(_00091_),
    .Q(\soc_I.clint_I.mtimecmp[12] ));
 sg13g2_dfrbp_1 _33921_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1976),
    .D(_00611_),
    .Q_N(_00095_),
    .Q(\soc_I.clint_I.mtimecmp[13] ));
 sg13g2_dfrbp_1 _33922_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1974),
    .D(_00612_),
    .Q_N(_00099_),
    .Q(\soc_I.clint_I.mtimecmp[14] ));
 sg13g2_dfrbp_1 _33923_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1972),
    .D(_00613_),
    .Q_N(_00103_),
    .Q(\soc_I.clint_I.mtimecmp[15] ));
 sg13g2_dfrbp_1 _33924_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1970),
    .D(_00614_),
    .Q_N(_00013_),
    .Q(\soc_I.clint_I.mtimecmp[16] ));
 sg13g2_dfrbp_1 _33925_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1968),
    .D(_00615_),
    .Q_N(_00020_),
    .Q(\soc_I.clint_I.mtimecmp[17] ));
 sg13g2_dfrbp_1 _33926_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1966),
    .D(_00616_),
    .Q_N(_00028_),
    .Q(\soc_I.clint_I.mtimecmp[18] ));
 sg13g2_dfrbp_1 _33927_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1964),
    .D(_00617_),
    .Q_N(_00036_),
    .Q(\soc_I.clint_I.mtimecmp[19] ));
 sg13g2_dfrbp_1 _33928_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1962),
    .D(_00618_),
    .Q_N(_00043_),
    .Q(\soc_I.clint_I.mtimecmp[20] ));
 sg13g2_dfrbp_1 _33929_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1960),
    .D(_00619_),
    .Q_N(_00050_),
    .Q(\soc_I.clint_I.mtimecmp[21] ));
 sg13g2_dfrbp_1 _33930_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1958),
    .D(_00620_),
    .Q_N(_00058_),
    .Q(\soc_I.clint_I.mtimecmp[22] ));
 sg13g2_dfrbp_1 _33931_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1956),
    .D(_00621_),
    .Q_N(_00066_),
    .Q(\soc_I.clint_I.mtimecmp[23] ));
 sg13g2_dfrbp_1 _33932_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1954),
    .D(_00622_),
    .Q_N(_00016_),
    .Q(\soc_I.clint_I.mtimecmp[24] ));
 sg13g2_dfrbp_1 _33933_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1952),
    .D(_00623_),
    .Q_N(_00024_),
    .Q(\soc_I.clint_I.mtimecmp[25] ));
 sg13g2_dfrbp_1 _33934_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1950),
    .D(_00624_),
    .Q_N(_00032_),
    .Q(\soc_I.clint_I.mtimecmp[26] ));
 sg13g2_dfrbp_1 _33935_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1948),
    .D(_00625_),
    .Q_N(_00040_),
    .Q(\soc_I.clint_I.mtimecmp[27] ));
 sg13g2_dfrbp_1 _33936_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1946),
    .D(_00626_),
    .Q_N(_00046_),
    .Q(\soc_I.clint_I.mtimecmp[28] ));
 sg13g2_dfrbp_1 _33937_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1944),
    .D(_00627_),
    .Q_N(_00054_),
    .Q(\soc_I.clint_I.mtimecmp[29] ));
 sg13g2_dfrbp_1 _33938_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1942),
    .D(_00628_),
    .Q_N(_00062_),
    .Q(\soc_I.clint_I.mtimecmp[30] ));
 sg13g2_dfrbp_1 _33939_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1940),
    .D(_00629_),
    .Q_N(_00071_),
    .Q(\soc_I.clint_I.mtimecmp[31] ));
 sg13g2_dfrbp_1 _33940_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1938),
    .D(_00630_),
    .Q_N(_16387_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[0][0] ));
 sg13g2_dfrbp_1 _33941_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1937),
    .D(net4329),
    .Q_N(_16386_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[0][1] ));
 sg13g2_dfrbp_1 _33942_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1936),
    .D(net3982),
    .Q_N(_16385_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[0][2] ));
 sg13g2_dfrbp_1 _33943_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1935),
    .D(net4143),
    .Q_N(_16384_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[0][3] ));
 sg13g2_dfrbp_1 _33944_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1934),
    .D(net4215),
    .Q_N(_16383_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[0][4] ));
 sg13g2_dfrbp_1 _33945_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1933),
    .D(_00635_),
    .Q_N(_16382_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[0][5] ));
 sg13g2_dfrbp_1 _33946_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1932),
    .D(net4128),
    .Q_N(_16381_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[0][6] ));
 sg13g2_dfrbp_1 _33947_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1931),
    .D(_00637_),
    .Q_N(_16380_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[0][7] ));
 sg13g2_dfrbp_1 _33948_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1930),
    .D(net2745),
    .Q_N(_16379_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[10][0] ));
 sg13g2_dfrbp_1 _33949_ (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1929),
    .D(net3640),
    .Q_N(_16378_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[10][1] ));
 sg13g2_dfrbp_1 _33950_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1928),
    .D(_00640_),
    .Q_N(_16377_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[10][2] ));
 sg13g2_dfrbp_1 _33951_ (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1927),
    .D(net4162),
    .Q_N(_16376_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[10][3] ));
 sg13g2_dfrbp_1 _33952_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1926),
    .D(net3753),
    .Q_N(_16375_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[10][4] ));
 sg13g2_dfrbp_1 _33953_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1925),
    .D(net3610),
    .Q_N(_16374_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[10][5] ));
 sg13g2_dfrbp_1 _33954_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1924),
    .D(net4105),
    .Q_N(_16373_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[10][6] ));
 sg13g2_dfrbp_1 _33955_ (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1923),
    .D(net4078),
    .Q_N(_16372_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[10][7] ));
 sg13g2_dfrbp_1 _33956_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1922),
    .D(net2711),
    .Q_N(_16371_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[11][0] ));
 sg13g2_dfrbp_1 _33957_ (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1921),
    .D(net4213),
    .Q_N(_16370_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[11][1] ));
 sg13g2_dfrbp_1 _33958_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1920),
    .D(_00648_),
    .Q_N(_16369_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[11][2] ));
 sg13g2_dfrbp_1 _33959_ (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1919),
    .D(net3913),
    .Q_N(_16368_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[11][3] ));
 sg13g2_dfrbp_1 _33960_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1918),
    .D(net4220),
    .Q_N(_16367_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[11][4] ));
 sg13g2_dfrbp_1 _33961_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1917),
    .D(net4100),
    .Q_N(_16366_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[11][5] ));
 sg13g2_dfrbp_1 _33962_ (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1916),
    .D(net4238),
    .Q_N(_16365_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[11][6] ));
 sg13g2_dfrbp_1 _33963_ (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1915),
    .D(_00653_),
    .Q_N(_16364_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[11][7] ));
 sg13g2_dfrbp_1 _33964_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1914),
    .D(net2649),
    .Q_N(_16363_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[12][0] ));
 sg13g2_dfrbp_1 _33965_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1913),
    .D(_00655_),
    .Q_N(_16362_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[12][1] ));
 sg13g2_dfrbp_1 _33966_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1912),
    .D(_00656_),
    .Q_N(_16361_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[12][2] ));
 sg13g2_dfrbp_1 _33967_ (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1911),
    .D(net4193),
    .Q_N(_16360_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[12][3] ));
 sg13g2_dfrbp_1 _33968_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1910),
    .D(net4110),
    .Q_N(_16359_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[12][4] ));
 sg13g2_dfrbp_1 _33969_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1909),
    .D(_00659_),
    .Q_N(_16358_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[12][5] ));
 sg13g2_dfrbp_1 _33970_ (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1908),
    .D(_00660_),
    .Q_N(_16357_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[12][6] ));
 sg13g2_dfrbp_1 _33971_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1907),
    .D(_00661_),
    .Q_N(_16356_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[12][7] ));
 sg13g2_dfrbp_1 _33972_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1906),
    .D(net3385),
    .Q_N(_16355_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[13][0] ));
 sg13g2_dfrbp_1 _33973_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1905),
    .D(_00663_),
    .Q_N(_16354_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[13][1] ));
 sg13g2_dfrbp_1 _33974_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1904),
    .D(_00664_),
    .Q_N(_16353_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[13][2] ));
 sg13g2_dfrbp_1 _33975_ (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1903),
    .D(net3432),
    .Q_N(_16352_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[13][3] ));
 sg13g2_dfrbp_1 _33976_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1902),
    .D(net3131),
    .Q_N(_16351_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[13][4] ));
 sg13g2_dfrbp_1 _33977_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1901),
    .D(_00667_),
    .Q_N(_16350_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[13][5] ));
 sg13g2_dfrbp_1 _33978_ (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1900),
    .D(_00668_),
    .Q_N(_16349_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[13][6] ));
 sg13g2_dfrbp_1 _33979_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1899),
    .D(_00669_),
    .Q_N(_16348_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[13][7] ));
 sg13g2_dfrbp_1 _33980_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1898),
    .D(net3986),
    .Q_N(_16347_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[14][0] ));
 sg13g2_dfrbp_1 _33981_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1897),
    .D(_00671_),
    .Q_N(_16346_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[14][1] ));
 sg13g2_dfrbp_1 _33982_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1896),
    .D(net2732),
    .Q_N(_16345_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[14][2] ));
 sg13g2_dfrbp_1 _33983_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1895),
    .D(net3260),
    .Q_N(_16344_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[14][3] ));
 sg13g2_dfrbp_1 _33984_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1894),
    .D(net3394),
    .Q_N(_16343_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[14][4] ));
 sg13g2_dfrbp_1 _33985_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1893),
    .D(_00675_),
    .Q_N(_16342_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[14][5] ));
 sg13g2_dfrbp_1 _33986_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1892),
    .D(_00676_),
    .Q_N(_16341_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[14][6] ));
 sg13g2_dfrbp_1 _33987_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1891),
    .D(_00677_),
    .Q_N(_16340_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[14][7] ));
 sg13g2_dfrbp_1 _33988_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1890),
    .D(_00678_),
    .Q_N(_16339_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][0] ));
 sg13g2_dfrbp_1 _33989_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1889),
    .D(_00679_),
    .Q_N(_16338_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][1] ));
 sg13g2_dfrbp_1 _33990_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1888),
    .D(_00680_),
    .Q_N(_16337_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][2] ));
 sg13g2_dfrbp_1 _33991_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1887),
    .D(_00681_),
    .Q_N(_16336_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][3] ));
 sg13g2_dfrbp_1 _33992_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1886),
    .D(_00682_),
    .Q_N(_16335_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][4] ));
 sg13g2_dfrbp_1 _33993_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1885),
    .D(_00683_),
    .Q_N(_16334_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][5] ));
 sg13g2_dfrbp_1 _33994_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1884),
    .D(_00684_),
    .Q_N(_16333_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][6] ));
 sg13g2_dfrbp_1 _33995_ (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1883),
    .D(_00685_),
    .Q_N(_16332_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][7] ));
 sg13g2_dfrbp_1 _33996_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1882),
    .D(_00686_),
    .Q_N(_16331_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][8] ));
 sg13g2_dfrbp_1 _33997_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1881),
    .D(_00687_),
    .Q_N(_16330_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][9] ));
 sg13g2_dfrbp_1 _33998_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1880),
    .D(_00688_),
    .Q_N(_16329_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][10] ));
 sg13g2_dfrbp_1 _33999_ (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1879),
    .D(_00689_),
    .Q_N(_16328_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][11] ));
 sg13g2_dfrbp_1 _34000_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1878),
    .D(_00690_),
    .Q_N(_16327_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][12] ));
 sg13g2_dfrbp_1 _34001_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1877),
    .D(_00691_),
    .Q_N(_16326_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][13] ));
 sg13g2_dfrbp_1 _34002_ (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1876),
    .D(_00692_),
    .Q_N(_16325_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][14] ));
 sg13g2_dfrbp_1 _34003_ (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1875),
    .D(_00693_),
    .Q_N(_16324_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][15] ));
 sg13g2_dfrbp_1 _34004_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1874),
    .D(_00694_),
    .Q_N(_16323_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][16] ));
 sg13g2_dfrbp_1 _34005_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1873),
    .D(_00695_),
    .Q_N(_16322_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][17] ));
 sg13g2_dfrbp_1 _34006_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1872),
    .D(_00696_),
    .Q_N(_16321_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][18] ));
 sg13g2_dfrbp_1 _34007_ (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1871),
    .D(_00697_),
    .Q_N(_16320_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][19] ));
 sg13g2_dfrbp_1 _34008_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1870),
    .D(_00698_),
    .Q_N(_16319_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][20] ));
 sg13g2_dfrbp_1 _34009_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1869),
    .D(_00699_),
    .Q_N(_16318_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][21] ));
 sg13g2_dfrbp_1 _34010_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1868),
    .D(_00700_),
    .Q_N(_16317_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][22] ));
 sg13g2_dfrbp_1 _34011_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1867),
    .D(_00701_),
    .Q_N(_16316_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][23] ));
 sg13g2_dfrbp_1 _34012_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1866),
    .D(_00702_),
    .Q_N(_16315_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][24] ));
 sg13g2_dfrbp_1 _34013_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1865),
    .D(_00703_),
    .Q_N(_16314_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][25] ));
 sg13g2_dfrbp_1 _34014_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1864),
    .D(_00704_),
    .Q_N(_16313_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][26] ));
 sg13g2_dfrbp_1 _34015_ (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1863),
    .D(_00705_),
    .Q_N(_16312_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][27] ));
 sg13g2_dfrbp_1 _34016_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1862),
    .D(_00706_),
    .Q_N(_16311_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][28] ));
 sg13g2_dfrbp_1 _34017_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1861),
    .D(_00707_),
    .Q_N(_16310_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][29] ));
 sg13g2_dfrbp_1 _34018_ (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1860),
    .D(_00708_),
    .Q_N(_16309_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][30] ));
 sg13g2_dfrbp_1 _34019_ (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1859),
    .D(_00709_),
    .Q_N(_16308_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][31] ));
 sg13g2_dfrbp_1 _34020_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1858),
    .D(_00710_),
    .Q_N(_16307_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][0] ));
 sg13g2_dfrbp_1 _34021_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1857),
    .D(_00711_),
    .Q_N(_16306_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][1] ));
 sg13g2_dfrbp_1 _34022_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1856),
    .D(_00712_),
    .Q_N(_16305_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][2] ));
 sg13g2_dfrbp_1 _34023_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1855),
    .D(_00713_),
    .Q_N(_16304_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][3] ));
 sg13g2_dfrbp_1 _34024_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1854),
    .D(_00714_),
    .Q_N(_16303_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][4] ));
 sg13g2_dfrbp_1 _34025_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1853),
    .D(_00715_),
    .Q_N(_16302_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][5] ));
 sg13g2_dfrbp_1 _34026_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1852),
    .D(_00716_),
    .Q_N(_16301_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][6] ));
 sg13g2_dfrbp_1 _34027_ (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1851),
    .D(_00717_),
    .Q_N(_16300_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][7] ));
 sg13g2_dfrbp_1 _34028_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1850),
    .D(_00718_),
    .Q_N(_16299_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][8] ));
 sg13g2_dfrbp_1 _34029_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1849),
    .D(_00719_),
    .Q_N(_16298_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][9] ));
 sg13g2_dfrbp_1 _34030_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1848),
    .D(_00720_),
    .Q_N(_16297_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][10] ));
 sg13g2_dfrbp_1 _34031_ (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1847),
    .D(_00721_),
    .Q_N(_16296_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][11] ));
 sg13g2_dfrbp_1 _34032_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1846),
    .D(_00722_),
    .Q_N(_16295_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][12] ));
 sg13g2_dfrbp_1 _34033_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1845),
    .D(_00723_),
    .Q_N(_16294_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][13] ));
 sg13g2_dfrbp_1 _34034_ (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1844),
    .D(_00724_),
    .Q_N(_16293_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][14] ));
 sg13g2_dfrbp_1 _34035_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1843),
    .D(net3904),
    .Q_N(_16292_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][15] ));
 sg13g2_dfrbp_1 _34036_ (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1842),
    .D(_00726_),
    .Q_N(_16291_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][16] ));
 sg13g2_dfrbp_1 _34037_ (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1841),
    .D(net2827),
    .Q_N(_16290_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][17] ));
 sg13g2_dfrbp_1 _34038_ (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1840),
    .D(_00728_),
    .Q_N(_16289_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][18] ));
 sg13g2_dfrbp_1 _34039_ (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1839),
    .D(_00729_),
    .Q_N(_16288_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][19] ));
 sg13g2_dfrbp_1 _34040_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1838),
    .D(_00730_),
    .Q_N(_16287_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][20] ));
 sg13g2_dfrbp_1 _34041_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1837),
    .D(_00731_),
    .Q_N(_16286_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][21] ));
 sg13g2_dfrbp_1 _34042_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1836),
    .D(_00732_),
    .Q_N(_16285_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][22] ));
 sg13g2_dfrbp_1 _34043_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1835),
    .D(_00733_),
    .Q_N(_16284_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][23] ));
 sg13g2_dfrbp_1 _34044_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1834),
    .D(_00734_),
    .Q_N(_16283_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][24] ));
 sg13g2_dfrbp_1 _34045_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1833),
    .D(_00735_),
    .Q_N(_16282_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][25] ));
 sg13g2_dfrbp_1 _34046_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1832),
    .D(_00736_),
    .Q_N(_16281_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][26] ));
 sg13g2_dfrbp_1 _34047_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1831),
    .D(_00737_),
    .Q_N(_16280_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][27] ));
 sg13g2_dfrbp_1 _34048_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1830),
    .D(_00738_),
    .Q_N(_16279_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][28] ));
 sg13g2_dfrbp_1 _34049_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1829),
    .D(_00739_),
    .Q_N(_16278_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][29] ));
 sg13g2_dfrbp_1 _34050_ (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1828),
    .D(_00740_),
    .Q_N(_16277_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][30] ));
 sg13g2_dfrbp_1 _34051_ (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1827),
    .D(_00741_),
    .Q_N(_16276_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][31] ));
 sg13g2_dfrbp_1 _34052_ (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1826),
    .D(_00742_),
    .Q_N(_16275_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[0] ));
 sg13g2_dfrbp_1 _34053_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1825),
    .D(_00743_),
    .Q_N(_16274_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[1] ));
 sg13g2_dfrbp_1 _34054_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1824),
    .D(_00744_),
    .Q_N(_16273_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[2] ));
 sg13g2_dfrbp_1 _34055_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1823),
    .D(_00745_),
    .Q_N(_16272_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[3] ));
 sg13g2_dfrbp_1 _34056_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1822),
    .D(_00746_),
    .Q_N(_16271_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[4] ));
 sg13g2_dfrbp_1 _34057_ (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1821),
    .D(_00747_),
    .Q_N(_16270_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[5] ));
 sg13g2_dfrbp_1 _34058_ (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1820),
    .D(_00748_),
    .Q_N(_16269_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[6] ));
 sg13g2_dfrbp_1 _34059_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1819),
    .D(_00749_),
    .Q_N(_16268_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[7] ));
 sg13g2_dfrbp_1 _34060_ (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1818),
    .D(_00750_),
    .Q_N(_16267_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[8] ));
 sg13g2_dfrbp_1 _34061_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1817),
    .D(_00751_),
    .Q_N(_16266_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[9] ));
 sg13g2_dfrbp_1 _34062_ (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1816),
    .D(_00752_),
    .Q_N(_16265_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[10] ));
 sg13g2_dfrbp_1 _34063_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1815),
    .D(_00753_),
    .Q_N(_16264_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[11] ));
 sg13g2_dfrbp_1 _34064_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1814),
    .D(_00754_),
    .Q_N(_16263_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[12] ));
 sg13g2_dfrbp_1 _34065_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1813),
    .D(_00755_),
    .Q_N(_16262_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[13] ));
 sg13g2_dfrbp_1 _34066_ (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1812),
    .D(_00756_),
    .Q_N(_16261_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[14] ));
 sg13g2_dfrbp_1 _34067_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1811),
    .D(_00757_),
    .Q_N(_16260_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[15] ));
 sg13g2_dfrbp_1 _34068_ (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1810),
    .D(_00758_),
    .Q_N(_16259_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[16] ));
 sg13g2_dfrbp_1 _34069_ (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1809),
    .D(_00759_),
    .Q_N(_16258_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[17] ));
 sg13g2_dfrbp_1 _34070_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1808),
    .D(_00760_),
    .Q_N(_16257_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[18] ));
 sg13g2_dfrbp_1 _34071_ (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1807),
    .D(_00761_),
    .Q_N(_16256_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[19] ));
 sg13g2_dfrbp_1 _34072_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1806),
    .D(_00762_),
    .Q_N(_16255_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[20] ));
 sg13g2_dfrbp_1 _34073_ (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1805),
    .D(_00763_),
    .Q_N(_16254_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[21] ));
 sg13g2_dfrbp_1 _34074_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1804),
    .D(_00764_),
    .Q_N(_16253_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[22] ));
 sg13g2_dfrbp_1 _34075_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1803),
    .D(_00765_),
    .Q_N(_16252_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[23] ));
 sg13g2_dfrbp_1 _34076_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1802),
    .D(_00766_),
    .Q_N(_16251_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[24] ));
 sg13g2_dfrbp_1 _34077_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1801),
    .D(_00767_),
    .Q_N(_16250_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[25] ));
 sg13g2_dfrbp_1 _34078_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1800),
    .D(_00768_),
    .Q_N(_16249_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[26] ));
 sg13g2_dfrbp_1 _34079_ (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1799),
    .D(_00769_),
    .Q_N(_16248_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[27] ));
 sg13g2_dfrbp_1 _34080_ (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1798),
    .D(_00770_),
    .Q_N(_16247_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[28] ));
 sg13g2_dfrbp_1 _34081_ (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1797),
    .D(_00771_),
    .Q_N(_16246_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[29] ));
 sg13g2_dfrbp_1 _34082_ (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1796),
    .D(_00772_),
    .Q_N(_16245_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[30] ));
 sg13g2_dfrbp_1 _34083_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1795),
    .D(_00773_),
    .Q_N(_16244_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A1[31] ));
 sg13g2_dfrbp_1 _34084_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1794),
    .D(net4705),
    .Q_N(_16243_),
    .Q(\soc_I.qqspi_I.xfer_cycles[0] ));
 sg13g2_dfrbp_1 _34085_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1792),
    .D(net4478),
    .Q_N(_16242_),
    .Q(\soc_I.qqspi_I.xfer_cycles[1] ));
 sg13g2_dfrbp_1 _34086_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1790),
    .D(_00776_),
    .Q_N(_16241_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][0] ));
 sg13g2_dfrbp_1 _34087_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1789),
    .D(_00777_),
    .Q_N(_16240_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][1] ));
 sg13g2_dfrbp_1 _34088_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1788),
    .D(_00778_),
    .Q_N(_16239_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][2] ));
 sg13g2_dfrbp_1 _34089_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1787),
    .D(_00779_),
    .Q_N(_16238_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][3] ));
 sg13g2_dfrbp_1 _34090_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1786),
    .D(_00780_),
    .Q_N(_16237_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][4] ));
 sg13g2_dfrbp_1 _34091_ (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1785),
    .D(_00781_),
    .Q_N(_16236_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][5] ));
 sg13g2_dfrbp_1 _34092_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1784),
    .D(_00782_),
    .Q_N(_16235_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][6] ));
 sg13g2_dfrbp_1 _34093_ (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1783),
    .D(_00783_),
    .Q_N(_16234_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][7] ));
 sg13g2_dfrbp_1 _34094_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1782),
    .D(_00784_),
    .Q_N(_16233_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][8] ));
 sg13g2_dfrbp_1 _34095_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1781),
    .D(_00785_),
    .Q_N(_16232_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][9] ));
 sg13g2_dfrbp_1 _34096_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1780),
    .D(_00786_),
    .Q_N(_16231_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][10] ));
 sg13g2_dfrbp_1 _34097_ (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1779),
    .D(_00787_),
    .Q_N(_16230_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][11] ));
 sg13g2_dfrbp_1 _34098_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net1778),
    .D(_00788_),
    .Q_N(_16229_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][12] ));
 sg13g2_dfrbp_1 _34099_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1777),
    .D(_00789_),
    .Q_N(_16228_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][13] ));
 sg13g2_dfrbp_1 _34100_ (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1776),
    .D(_00790_),
    .Q_N(_16227_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][14] ));
 sg13g2_dfrbp_1 _34101_ (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1775),
    .D(_00791_),
    .Q_N(_16226_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][15] ));
 sg13g2_dfrbp_1 _34102_ (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1774),
    .D(_00792_),
    .Q_N(_16225_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][16] ));
 sg13g2_dfrbp_1 _34103_ (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1773),
    .D(_00793_),
    .Q_N(_16224_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][17] ));
 sg13g2_dfrbp_1 _34104_ (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1772),
    .D(_00794_),
    .Q_N(_16223_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][18] ));
 sg13g2_dfrbp_1 _34105_ (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1771),
    .D(_00795_),
    .Q_N(_16222_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][19] ));
 sg13g2_dfrbp_1 _34106_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1770),
    .D(_00796_),
    .Q_N(_16221_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][20] ));
 sg13g2_dfrbp_1 _34107_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1769),
    .D(_00797_),
    .Q_N(_16220_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][21] ));
 sg13g2_dfrbp_1 _34108_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1768),
    .D(_00798_),
    .Q_N(_16219_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][22] ));
 sg13g2_dfrbp_1 _34109_ (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1767),
    .D(_00799_),
    .Q_N(_16218_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][23] ));
 sg13g2_dfrbp_1 _34110_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1766),
    .D(_00800_),
    .Q_N(_16217_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][24] ));
 sg13g2_dfrbp_1 _34111_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1765),
    .D(_00801_),
    .Q_N(_16216_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][25] ));
 sg13g2_dfrbp_1 _34112_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1764),
    .D(_00802_),
    .Q_N(_16215_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][26] ));
 sg13g2_dfrbp_1 _34113_ (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1763),
    .D(_00803_),
    .Q_N(_16214_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][27] ));
 sg13g2_dfrbp_1 _34114_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1762),
    .D(_00804_),
    .Q_N(_16213_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][28] ));
 sg13g2_dfrbp_1 _34115_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1761),
    .D(_00805_),
    .Q_N(_16212_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][29] ));
 sg13g2_dfrbp_1 _34116_ (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1760),
    .D(_00806_),
    .Q_N(_16211_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][30] ));
 sg13g2_dfrbp_1 _34117_ (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1759),
    .D(_00807_),
    .Q_N(_16210_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][31] ));
 sg13g2_dfrbp_1 _34118_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1758),
    .D(_00808_),
    .Q_N(_16209_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][0] ));
 sg13g2_dfrbp_1 _34119_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1757),
    .D(_00809_),
    .Q_N(_16208_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][1] ));
 sg13g2_dfrbp_1 _34120_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1756),
    .D(_00810_),
    .Q_N(_16207_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][2] ));
 sg13g2_dfrbp_1 _34121_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1755),
    .D(_00811_),
    .Q_N(_16206_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][3] ));
 sg13g2_dfrbp_1 _34122_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1754),
    .D(_00812_),
    .Q_N(_16205_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][4] ));
 sg13g2_dfrbp_1 _34123_ (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1753),
    .D(_00813_),
    .Q_N(_16204_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][5] ));
 sg13g2_dfrbp_1 _34124_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1752),
    .D(_00814_),
    .Q_N(_16203_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][6] ));
 sg13g2_dfrbp_1 _34125_ (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1751),
    .D(_00815_),
    .Q_N(_16202_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][7] ));
 sg13g2_dfrbp_1 _34126_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1750),
    .D(_00816_),
    .Q_N(_16201_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][8] ));
 sg13g2_dfrbp_1 _34127_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1749),
    .D(_00817_),
    .Q_N(_16200_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][9] ));
 sg13g2_dfrbp_1 _34128_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1748),
    .D(_00818_),
    .Q_N(_16199_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][10] ));
 sg13g2_dfrbp_1 _34129_ (.CLK(clknet_leaf_319_clk),
    .RESET_B(net1747),
    .D(_00819_),
    .Q_N(_16198_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][11] ));
 sg13g2_dfrbp_1 _34130_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1746),
    .D(_00820_),
    .Q_N(_16197_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][12] ));
 sg13g2_dfrbp_1 _34131_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1745),
    .D(_00821_),
    .Q_N(_16196_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][13] ));
 sg13g2_dfrbp_1 _34132_ (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1744),
    .D(_00822_),
    .Q_N(_16195_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][14] ));
 sg13g2_dfrbp_1 _34133_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1743),
    .D(_00823_),
    .Q_N(_16194_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][15] ));
 sg13g2_dfrbp_1 _34134_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1742),
    .D(_00824_),
    .Q_N(_16193_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][16] ));
 sg13g2_dfrbp_1 _34135_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1741),
    .D(_00825_),
    .Q_N(_16192_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][17] ));
 sg13g2_dfrbp_1 _34136_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1740),
    .D(_00826_),
    .Q_N(_16191_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][18] ));
 sg13g2_dfrbp_1 _34137_ (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1739),
    .D(_00827_),
    .Q_N(_16190_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][19] ));
 sg13g2_dfrbp_1 _34138_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1738),
    .D(_00828_),
    .Q_N(_16189_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][20] ));
 sg13g2_dfrbp_1 _34139_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1737),
    .D(_00829_),
    .Q_N(_16188_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][21] ));
 sg13g2_dfrbp_1 _34140_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1736),
    .D(_00830_),
    .Q_N(_16187_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][22] ));
 sg13g2_dfrbp_1 _34141_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1735),
    .D(_00831_),
    .Q_N(_16186_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][23] ));
 sg13g2_dfrbp_1 _34142_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1734),
    .D(_00832_),
    .Q_N(_16185_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][24] ));
 sg13g2_dfrbp_1 _34143_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1733),
    .D(_00833_),
    .Q_N(_16184_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][25] ));
 sg13g2_dfrbp_1 _34144_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1732),
    .D(_00834_),
    .Q_N(_16183_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][26] ));
 sg13g2_dfrbp_1 _34145_ (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1731),
    .D(_00835_),
    .Q_N(_16182_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][27] ));
 sg13g2_dfrbp_1 _34146_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1730),
    .D(_00836_),
    .Q_N(_16181_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][28] ));
 sg13g2_dfrbp_1 _34147_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1729),
    .D(_00837_),
    .Q_N(_16180_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][29] ));
 sg13g2_dfrbp_1 _34148_ (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1728),
    .D(_00838_),
    .Q_N(_16179_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][30] ));
 sg13g2_dfrbp_1 _34149_ (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1727),
    .D(_00839_),
    .Q_N(_16178_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][31] ));
 sg13g2_dfrbp_1 _34150_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1726),
    .D(_00840_),
    .Q_N(_16177_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[0] ));
 sg13g2_dfrbp_1 _34151_ (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1724),
    .D(_00841_),
    .Q_N(_16176_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[1] ));
 sg13g2_dfrbp_1 _34152_ (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1722),
    .D(_00842_),
    .Q_N(_16175_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[2] ));
 sg13g2_dfrbp_1 _34153_ (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1720),
    .D(_00843_),
    .Q_N(_16174_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[3] ));
 sg13g2_dfrbp_1 _34154_ (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1718),
    .D(_00844_),
    .Q_N(_16173_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[4] ));
 sg13g2_dfrbp_1 _34155_ (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1716),
    .D(_00845_),
    .Q_N(_16172_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[5] ));
 sg13g2_dfrbp_1 _34156_ (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1714),
    .D(_00846_),
    .Q_N(_16171_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[6] ));
 sg13g2_dfrbp_1 _34157_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1712),
    .D(_00847_),
    .Q_N(_16170_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[7] ));
 sg13g2_dfrbp_1 _34158_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1710),
    .D(_00848_),
    .Q_N(_16169_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[8] ));
 sg13g2_dfrbp_1 _34159_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1708),
    .D(_00849_),
    .Q_N(_16168_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[9] ));
 sg13g2_dfrbp_1 _34160_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1706),
    .D(net4258),
    .Q_N(_16167_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[10] ));
 sg13g2_dfrbp_1 _34161_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1704),
    .D(_00851_),
    .Q_N(_16166_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[11] ));
 sg13g2_dfrbp_1 _34162_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1702),
    .D(_00852_),
    .Q_N(_16165_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[12] ));
 sg13g2_dfrbp_1 _34163_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1700),
    .D(_00853_),
    .Q_N(_16164_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[13] ));
 sg13g2_dfrbp_1 _34164_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1698),
    .D(net4624),
    .Q_N(_16163_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[14] ));
 sg13g2_dfrbp_1 _34165_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1696),
    .D(_00855_),
    .Q_N(_16162_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[15] ));
 sg13g2_dfrbp_1 _34166_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1694),
    .D(net4460),
    .Q_N(_16161_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[16] ));
 sg13g2_dfrbp_1 _34167_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1692),
    .D(net4358),
    .Q_N(_16160_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[17] ));
 sg13g2_dfrbp_1 _34168_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1690),
    .D(net4869),
    .Q_N(_16159_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[18] ));
 sg13g2_dfrbp_1 _34169_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1688),
    .D(net4789),
    .Q_N(_16158_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[19] ));
 sg13g2_dfrbp_1 _34170_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1686),
    .D(net4679),
    .Q_N(_16157_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[20] ));
 sg13g2_dfrbp_1 _34171_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1684),
    .D(net4728),
    .Q_N(_16156_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[21] ));
 sg13g2_dfrbp_1 _34172_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1682),
    .D(net4742),
    .Q_N(_16155_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[22] ));
 sg13g2_dfrbp_1 _34173_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1680),
    .D(_00863_),
    .Q_N(_16154_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[23] ));
 sg13g2_dfrbp_1 _34174_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1678),
    .D(net4578),
    .Q_N(_16153_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[24] ));
 sg13g2_dfrbp_1 _34175_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1676),
    .D(net4653),
    .Q_N(_16152_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[25] ));
 sg13g2_dfrbp_1 _34176_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1674),
    .D(net4731),
    .Q_N(_16151_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[26] ));
 sg13g2_dfrbp_1 _34177_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1672),
    .D(net4457),
    .Q_N(_16150_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[27] ));
 sg13g2_dfrbp_1 _34178_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1670),
    .D(net4573),
    .Q_N(_16149_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[28] ));
 sg13g2_dfrbp_1 _34179_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1668),
    .D(net4462),
    .Q_N(_16148_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[29] ));
 sg13g2_dfrbp_1 _34180_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1666),
    .D(net4506),
    .Q_N(_16147_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[30] ));
 sg13g2_dfrbp_1 _34181_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1664),
    .D(net4651),
    .Q_N(_16146_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[31] ));
 sg13g2_dfrbp_1 _34182_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1662),
    .D(_00872_),
    .Q_N(_16145_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[0] ));
 sg13g2_dfrbp_1 _34183_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1660),
    .D(_00873_),
    .Q_N(_16144_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[1] ));
 sg13g2_dfrbp_1 _34184_ (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1658),
    .D(_00874_),
    .Q_N(_16143_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[2] ));
 sg13g2_dfrbp_1 _34185_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1656),
    .D(_00875_),
    .Q_N(_16142_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[3] ));
 sg13g2_dfrbp_1 _34186_ (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1654),
    .D(_00876_),
    .Q_N(_16141_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[4] ));
 sg13g2_dfrbp_1 _34187_ (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1652),
    .D(_00877_),
    .Q_N(_16140_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[5] ));
 sg13g2_dfrbp_1 _34188_ (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1650),
    .D(_00878_),
    .Q_N(_16139_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[6] ));
 sg13g2_dfrbp_1 _34189_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1648),
    .D(_00879_),
    .Q_N(_16138_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[7] ));
 sg13g2_dfrbp_1 _34190_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1646),
    .D(_00880_),
    .Q_N(_16137_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[8] ));
 sg13g2_dfrbp_1 _34191_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1644),
    .D(_00881_),
    .Q_N(_16136_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[9] ));
 sg13g2_dfrbp_1 _34192_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1642),
    .D(_00882_),
    .Q_N(_16135_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[10] ));
 sg13g2_dfrbp_1 _34193_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1640),
    .D(_00883_),
    .Q_N(_16134_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[11] ));
 sg13g2_dfrbp_1 _34194_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1638),
    .D(_00884_),
    .Q_N(_16133_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[12] ));
 sg13g2_dfrbp_1 _34195_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1636),
    .D(_00885_),
    .Q_N(_16132_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[13] ));
 sg13g2_dfrbp_1 _34196_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1634),
    .D(_00886_),
    .Q_N(_16131_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[14] ));
 sg13g2_dfrbp_1 _34197_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1632),
    .D(_00887_),
    .Q_N(_16130_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[15] ));
 sg13g2_dfrbp_1 _34198_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1630),
    .D(_00888_),
    .Q_N(_16129_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[16] ));
 sg13g2_dfrbp_1 _34199_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1628),
    .D(_00889_),
    .Q_N(_16128_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[17] ));
 sg13g2_dfrbp_1 _34200_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1626),
    .D(_00890_),
    .Q_N(_16127_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[18] ));
 sg13g2_dfrbp_1 _34201_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1624),
    .D(_00891_),
    .Q_N(_16126_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[19] ));
 sg13g2_dfrbp_1 _34202_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1622),
    .D(_00892_),
    .Q_N(_16125_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[20] ));
 sg13g2_dfrbp_1 _34203_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1620),
    .D(_00893_),
    .Q_N(_16124_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[21] ));
 sg13g2_dfrbp_1 _34204_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1618),
    .D(_00894_),
    .Q_N(_16123_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[22] ));
 sg13g2_dfrbp_1 _34205_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1616),
    .D(_00895_),
    .Q_N(_16122_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[23] ));
 sg13g2_dfrbp_1 _34206_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1614),
    .D(_00896_),
    .Q_N(_16121_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[24] ));
 sg13g2_dfrbp_1 _34207_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1612),
    .D(_00897_),
    .Q_N(_16120_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[25] ));
 sg13g2_dfrbp_1 _34208_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1610),
    .D(_00898_),
    .Q_N(_16119_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[26] ));
 sg13g2_dfrbp_1 _34209_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1608),
    .D(_00899_),
    .Q_N(_16118_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[27] ));
 sg13g2_dfrbp_1 _34210_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1606),
    .D(_00900_),
    .Q_N(_16117_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[28] ));
 sg13g2_dfrbp_1 _34211_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1604),
    .D(_00901_),
    .Q_N(_16116_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[29] ));
 sg13g2_dfrbp_1 _34212_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1602),
    .D(_00902_),
    .Q_N(_16115_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[30] ));
 sg13g2_dfrbp_1 _34213_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1600),
    .D(_00903_),
    .Q_N(_16114_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[31] ));
 sg13g2_dfrbp_1 _34214_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1598),
    .D(_00904_),
    .Q_N(_16113_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[0] ));
 sg13g2_dfrbp_1 _34215_ (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1596),
    .D(_00905_),
    .Q_N(_16112_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[1] ));
 sg13g2_dfrbp_1 _34216_ (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1594),
    .D(_00906_),
    .Q_N(_16111_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[2] ));
 sg13g2_dfrbp_1 _34217_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1592),
    .D(_00907_),
    .Q_N(_16110_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[3] ));
 sg13g2_dfrbp_1 _34218_ (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1590),
    .D(net4854),
    .Q_N(_16109_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[4] ));
 sg13g2_dfrbp_1 _34219_ (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1588),
    .D(net4696),
    .Q_N(_16108_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[5] ));
 sg13g2_dfrbp_1 _34220_ (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1586),
    .D(net4733),
    .Q_N(_16107_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[6] ));
 sg13g2_dfrbp_1 _34221_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1584),
    .D(_00911_),
    .Q_N(_16106_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[7] ));
 sg13g2_dfrbp_1 _34222_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1582),
    .D(_00912_),
    .Q_N(_16105_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[8] ));
 sg13g2_dfrbp_1 _34223_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1580),
    .D(_00913_),
    .Q_N(_16104_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[9] ));
 sg13g2_dfrbp_1 _34224_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1578),
    .D(_00914_),
    .Q_N(_16103_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[10] ));
 sg13g2_dfrbp_1 _34225_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1576),
    .D(_00915_),
    .Q_N(_16102_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[11] ));
 sg13g2_dfrbp_1 _34226_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1574),
    .D(_00916_),
    .Q_N(_16101_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[12] ));
 sg13g2_dfrbp_1 _34227_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1572),
    .D(_00917_),
    .Q_N(_16100_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[13] ));
 sg13g2_dfrbp_1 _34228_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1570),
    .D(net4882),
    .Q_N(_16099_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[14] ));
 sg13g2_dfrbp_1 _34229_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1568),
    .D(_00919_),
    .Q_N(_16098_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[15] ));
 sg13g2_dfrbp_1 _34230_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1566),
    .D(net4993),
    .Q_N(_16097_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[16] ));
 sg13g2_dfrbp_1 _34231_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1564),
    .D(net4884),
    .Q_N(_16096_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[17] ));
 sg13g2_dfrbp_1 _34232_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1562),
    .D(_00922_),
    .Q_N(_16095_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[18] ));
 sg13g2_dfrbp_1 _34233_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1560),
    .D(net4906),
    .Q_N(_16094_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[19] ));
 sg13g2_dfrbp_1 _34234_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1558),
    .D(_00924_),
    .Q_N(_16093_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[20] ));
 sg13g2_dfrbp_1 _34235_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1556),
    .D(_00925_),
    .Q_N(_16092_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[21] ));
 sg13g2_dfrbp_1 _34236_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1554),
    .D(_00926_),
    .Q_N(_16091_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[22] ));
 sg13g2_dfrbp_1 _34237_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1552),
    .D(_00927_),
    .Q_N(_16090_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[23] ));
 sg13g2_dfrbp_1 _34238_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1550),
    .D(_00928_),
    .Q_N(_16089_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[24] ));
 sg13g2_dfrbp_1 _34239_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1548),
    .D(_00929_),
    .Q_N(_16088_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[25] ));
 sg13g2_dfrbp_1 _34240_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1546),
    .D(net4877),
    .Q_N(_16087_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[26] ));
 sg13g2_dfrbp_1 _34241_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1544),
    .D(_00931_),
    .Q_N(_16086_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[27] ));
 sg13g2_dfrbp_1 _34242_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1542),
    .D(_00932_),
    .Q_N(_16085_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[28] ));
 sg13g2_dfrbp_1 _34243_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1540),
    .D(_00933_),
    .Q_N(_16084_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[29] ));
 sg13g2_dfrbp_1 _34244_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1538),
    .D(_00934_),
    .Q_N(_16083_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[30] ));
 sg13g2_dfrbp_1 _34245_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1536),
    .D(_00935_),
    .Q_N(_16082_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[31] ));
 sg13g2_dfrbp_1 _34246_ (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1534),
    .D(_00936_),
    .Q_N(_16081_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[0] ));
 sg13g2_dfrbp_1 _34247_ (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1532),
    .D(_00937_),
    .Q_N(_16080_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[1] ));
 sg13g2_dfrbp_1 _34248_ (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1530),
    .D(_00938_),
    .Q_N(_16079_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[2] ));
 sg13g2_dfrbp_1 _34249_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1528),
    .D(_00939_),
    .Q_N(_16078_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[3] ));
 sg13g2_dfrbp_1 _34250_ (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1526),
    .D(_00940_),
    .Q_N(_16077_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[4] ));
 sg13g2_dfrbp_1 _34251_ (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1524),
    .D(_00941_),
    .Q_N(_16076_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[5] ));
 sg13g2_dfrbp_1 _34252_ (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1522),
    .D(_00942_),
    .Q_N(_16075_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[6] ));
 sg13g2_dfrbp_1 _34253_ (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1520),
    .D(_00943_),
    .Q_N(_16074_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[7] ));
 sg13g2_dfrbp_1 _34254_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1518),
    .D(_00944_),
    .Q_N(_16073_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[8] ));
 sg13g2_dfrbp_1 _34255_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1516),
    .D(_00945_),
    .Q_N(_16072_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[9] ));
 sg13g2_dfrbp_1 _34256_ (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1514),
    .D(_00946_),
    .Q_N(_16071_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[10] ));
 sg13g2_dfrbp_1 _34257_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1512),
    .D(_00947_),
    .Q_N(_16070_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[11] ));
 sg13g2_dfrbp_1 _34258_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1510),
    .D(_00948_),
    .Q_N(_16069_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[12] ));
 sg13g2_dfrbp_1 _34259_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1508),
    .D(_00949_),
    .Q_N(_16068_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[13] ));
 sg13g2_dfrbp_1 _34260_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1506),
    .D(_00950_),
    .Q_N(_16067_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[14] ));
 sg13g2_dfrbp_1 _34261_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1504),
    .D(_00951_),
    .Q_N(_16066_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[15] ));
 sg13g2_dfrbp_1 _34262_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1502),
    .D(_00952_),
    .Q_N(_16065_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[16] ));
 sg13g2_dfrbp_1 _34263_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1500),
    .D(_00953_),
    .Q_N(_16064_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[17] ));
 sg13g2_dfrbp_1 _34264_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1498),
    .D(_00954_),
    .Q_N(_16063_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[18] ));
 sg13g2_dfrbp_1 _34265_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1496),
    .D(_00955_),
    .Q_N(_16062_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[19] ));
 sg13g2_dfrbp_1 _34266_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1494),
    .D(_00956_),
    .Q_N(_16061_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[20] ));
 sg13g2_dfrbp_1 _34267_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1492),
    .D(_00957_),
    .Q_N(_16060_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[21] ));
 sg13g2_dfrbp_1 _34268_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1490),
    .D(_00958_),
    .Q_N(_16059_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[22] ));
 sg13g2_dfrbp_1 _34269_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1488),
    .D(_00959_),
    .Q_N(_16058_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[23] ));
 sg13g2_dfrbp_1 _34270_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1486),
    .D(_00960_),
    .Q_N(_16057_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[24] ));
 sg13g2_dfrbp_1 _34271_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1484),
    .D(_00961_),
    .Q_N(_16056_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[25] ));
 sg13g2_dfrbp_1 _34272_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1482),
    .D(_00962_),
    .Q_N(_16055_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[26] ));
 sg13g2_dfrbp_1 _34273_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1480),
    .D(_00963_),
    .Q_N(_16054_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[27] ));
 sg13g2_dfrbp_1 _34274_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1478),
    .D(_00964_),
    .Q_N(_16053_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[28] ));
 sg13g2_dfrbp_1 _34275_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1476),
    .D(_00965_),
    .Q_N(_16052_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[29] ));
 sg13g2_dfrbp_1 _34276_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1474),
    .D(_00966_),
    .Q_N(_16051_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[30] ));
 sg13g2_dfrbp_1 _34277_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1472),
    .D(_00967_),
    .Q_N(_16050_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[31] ));
 sg13g2_dfrbp_1 _34278_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1470),
    .D(_00968_),
    .Q_N(_16049_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[0] ));
 sg13g2_dfrbp_1 _34279_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1468),
    .D(_00969_),
    .Q_N(_16048_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[1] ));
 sg13g2_dfrbp_1 _34280_ (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1466),
    .D(_00970_),
    .Q_N(_16047_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[2] ));
 sg13g2_dfrbp_1 _34281_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1464),
    .D(_00971_),
    .Q_N(_16046_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[3] ));
 sg13g2_dfrbp_1 _34282_ (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1462),
    .D(_00972_),
    .Q_N(_16045_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[4] ));
 sg13g2_dfrbp_1 _34283_ (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1460),
    .D(_00973_),
    .Q_N(_16044_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[5] ));
 sg13g2_dfrbp_1 _34284_ (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1458),
    .D(_00974_),
    .Q_N(_16043_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[6] ));
 sg13g2_dfrbp_1 _34285_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1456),
    .D(_00975_),
    .Q_N(_16042_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[7] ));
 sg13g2_dfrbp_1 _34286_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1454),
    .D(_00976_),
    .Q_N(_16041_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[8] ));
 sg13g2_dfrbp_1 _34287_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1452),
    .D(_00977_),
    .Q_N(_16040_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[9] ));
 sg13g2_dfrbp_1 _34288_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1450),
    .D(_00978_),
    .Q_N(_16039_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[10] ));
 sg13g2_dfrbp_1 _34289_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1448),
    .D(_00979_),
    .Q_N(_16038_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[11] ));
 sg13g2_dfrbp_1 _34290_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1446),
    .D(_00980_),
    .Q_N(_16037_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[12] ));
 sg13g2_dfrbp_1 _34291_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1444),
    .D(_00981_),
    .Q_N(_16036_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[13] ));
 sg13g2_dfrbp_1 _34292_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1442),
    .D(_00982_),
    .Q_N(_16035_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[14] ));
 sg13g2_dfrbp_1 _34293_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1440),
    .D(_00983_),
    .Q_N(_16034_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[15] ));
 sg13g2_dfrbp_1 _34294_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1438),
    .D(_00984_),
    .Q_N(_16033_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[16] ));
 sg13g2_dfrbp_1 _34295_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1436),
    .D(_00985_),
    .Q_N(_16032_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[17] ));
 sg13g2_dfrbp_1 _34296_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1434),
    .D(_00986_),
    .Q_N(_16031_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[18] ));
 sg13g2_dfrbp_1 _34297_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1432),
    .D(_00987_),
    .Q_N(_16030_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[19] ));
 sg13g2_dfrbp_1 _34298_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1430),
    .D(_00988_),
    .Q_N(_16029_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[20] ));
 sg13g2_dfrbp_1 _34299_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1428),
    .D(_00989_),
    .Q_N(_16028_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[21] ));
 sg13g2_dfrbp_1 _34300_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1426),
    .D(_00990_),
    .Q_N(_16027_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[22] ));
 sg13g2_dfrbp_1 _34301_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1424),
    .D(_00991_),
    .Q_N(_16026_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[23] ));
 sg13g2_dfrbp_1 _34302_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1422),
    .D(_00992_),
    .Q_N(_16025_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[24] ));
 sg13g2_dfrbp_1 _34303_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1420),
    .D(_00993_),
    .Q_N(_16024_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[25] ));
 sg13g2_dfrbp_1 _34304_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1418),
    .D(_00994_),
    .Q_N(_16023_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[26] ));
 sg13g2_dfrbp_1 _34305_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1416),
    .D(_00995_),
    .Q_N(_16022_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[27] ));
 sg13g2_dfrbp_1 _34306_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1414),
    .D(_00996_),
    .Q_N(_16021_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[28] ));
 sg13g2_dfrbp_1 _34307_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1412),
    .D(_00997_),
    .Q_N(_16020_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[29] ));
 sg13g2_dfrbp_1 _34308_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1410),
    .D(_00998_),
    .Q_N(_16019_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[30] ));
 sg13g2_dfrbp_1 _34309_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1408),
    .D(_00999_),
    .Q_N(_16018_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[31] ));
 sg13g2_dfrbp_1 _34310_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1404),
    .D(_01000_),
    .Q_N(_16017_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_select ));
 sg13g2_dfrbp_1 _34311_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1307),
    .D(_01001_),
    .Q_N(_16016_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mip[3] ));
 sg13g2_dfrbp_1 _34312_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1306),
    .D(_01002_),
    .Q_N(_16015_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mip[7] ));
 sg13g2_dfrbp_1 _34313_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1305),
    .D(_01003_),
    .Q_N(_16014_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[0] ));
 sg13g2_dfrbp_1 _34314_ (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1303),
    .D(_01004_),
    .Q_N(_16013_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[1] ));
 sg13g2_dfrbp_1 _34315_ (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1301),
    .D(net4323),
    .Q_N(_16012_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[2] ));
 sg13g2_dfrbp_1 _34316_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1299),
    .D(net4145),
    .Q_N(_16011_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[3] ));
 sg13g2_dfrbp_1 _34317_ (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1297),
    .D(_01007_),
    .Q_N(_16010_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[4] ));
 sg13g2_dfrbp_1 _34318_ (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1295),
    .D(_01008_),
    .Q_N(_16009_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[5] ));
 sg13g2_dfrbp_1 _34319_ (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1293),
    .D(net3925),
    .Q_N(_16008_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[6] ));
 sg13g2_dfrbp_1 _34320_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1291),
    .D(net4230),
    .Q_N(_16007_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[7] ));
 sg13g2_dfrbp_1 _34321_ (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1289),
    .D(_01011_),
    .Q_N(_16006_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[8] ));
 sg13g2_dfrbp_1 _34322_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1287),
    .D(_01012_),
    .Q_N(_16005_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[9] ));
 sg13g2_dfrbp_1 _34323_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1285),
    .D(net4057),
    .Q_N(_16004_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[10] ));
 sg13g2_dfrbp_1 _34324_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1283),
    .D(net4179),
    .Q_N(_16003_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[11] ));
 sg13g2_dfrbp_1 _34325_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1281),
    .D(net4135),
    .Q_N(_16002_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[12] ));
 sg13g2_dfrbp_1 _34326_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1279),
    .D(net4125),
    .Q_N(_16001_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[13] ));
 sg13g2_dfrbp_1 _34327_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1277),
    .D(net4340),
    .Q_N(_16000_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[14] ));
 sg13g2_dfrbp_1 _34328_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1275),
    .D(net4141),
    .Q_N(_15999_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[15] ));
 sg13g2_dfrbp_1 _34329_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1273),
    .D(net4205),
    .Q_N(_15998_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[16] ));
 sg13g2_dfrbp_1 _34330_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1271),
    .D(net4248),
    .Q_N(_15997_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[17] ));
 sg13g2_dfrbp_1 _34331_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1269),
    .D(net4417),
    .Q_N(_15996_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[18] ));
 sg13g2_dfrbp_1 _34332_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1267),
    .D(net4552),
    .Q_N(_15995_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[19] ));
 sg13g2_dfrbp_1 _34333_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1265),
    .D(net4234),
    .Q_N(_15994_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[20] ));
 sg13g2_dfrbp_1 _34334_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1263),
    .D(net3970),
    .Q_N(_15993_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[21] ));
 sg13g2_dfrbp_1 _34335_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1261),
    .D(net4405),
    .Q_N(_15992_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[22] ));
 sg13g2_dfrbp_1 _34336_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1259),
    .D(net4424),
    .Q_N(_15991_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[23] ));
 sg13g2_dfrbp_1 _34337_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1257),
    .D(net4121),
    .Q_N(_15990_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[24] ));
 sg13g2_dfrbp_1 _34338_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1255),
    .D(net4088),
    .Q_N(_15989_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[25] ));
 sg13g2_dfrbp_1 _34339_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1253),
    .D(net4265),
    .Q_N(_15988_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[26] ));
 sg13g2_dfrbp_1 _34340_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1251),
    .D(net4964),
    .Q_N(_15987_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[27] ));
 sg13g2_dfrbp_1 _34341_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1249),
    .D(net4691),
    .Q_N(_15986_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[28] ));
 sg13g2_dfrbp_1 _34342_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1247),
    .D(net4875),
    .Q_N(_15985_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[29] ));
 sg13g2_dfrbp_1 _34343_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1245),
    .D(net3887),
    .Q_N(_15984_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[30] ));
 sg13g2_dfrbp_1 _34344_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1243),
    .D(net4791),
    .Q_N(_15983_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[31] ));
 sg13g2_dfrbp_1 _34345_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1241),
    .D(_01035_),
    .Q_N(_15982_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[0] ));
 sg13g2_dfrbp_1 _34346_ (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1239),
    .D(_01036_),
    .Q_N(_15981_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[1] ));
 sg13g2_dfrbp_1 _34347_ (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1237),
    .D(_01037_),
    .Q_N(_15980_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[2] ));
 sg13g2_dfrbp_1 _34348_ (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1235),
    .D(_01038_),
    .Q_N(_15979_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[3] ));
 sg13g2_dfrbp_1 _34349_ (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1233),
    .D(_01039_),
    .Q_N(_15978_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[4] ));
 sg13g2_dfrbp_1 _34350_ (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1231),
    .D(_01040_),
    .Q_N(_15977_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[5] ));
 sg13g2_dfrbp_1 _34351_ (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1229),
    .D(_01041_),
    .Q_N(_15976_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[6] ));
 sg13g2_dfrbp_1 _34352_ (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1227),
    .D(_01042_),
    .Q_N(_15975_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[7] ));
 sg13g2_dfrbp_1 _34353_ (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1225),
    .D(_01043_),
    .Q_N(_15974_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[8] ));
 sg13g2_dfrbp_1 _34354_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1223),
    .D(_01044_),
    .Q_N(_15973_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[9] ));
 sg13g2_dfrbp_1 _34355_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1221),
    .D(_01045_),
    .Q_N(_15972_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[10] ));
 sg13g2_dfrbp_1 _34356_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1219),
    .D(_01046_),
    .Q_N(_15971_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[11] ));
 sg13g2_dfrbp_1 _34357_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1217),
    .D(_01047_),
    .Q_N(_15970_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[12] ));
 sg13g2_dfrbp_1 _34358_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1215),
    .D(_01048_),
    .Q_N(_15969_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[13] ));
 sg13g2_dfrbp_1 _34359_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1213),
    .D(_01049_),
    .Q_N(_15968_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[14] ));
 sg13g2_dfrbp_1 _34360_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1211),
    .D(_01050_),
    .Q_N(_15967_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[15] ));
 sg13g2_dfrbp_1 _34361_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1209),
    .D(_01051_),
    .Q_N(_15966_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[16] ));
 sg13g2_dfrbp_1 _34362_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1207),
    .D(_01052_),
    .Q_N(_15965_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[17] ));
 sg13g2_dfrbp_1 _34363_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1205),
    .D(_01053_),
    .Q_N(_15964_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[18] ));
 sg13g2_dfrbp_1 _34364_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1203),
    .D(_01054_),
    .Q_N(_15963_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[19] ));
 sg13g2_dfrbp_1 _34365_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1201),
    .D(_01055_),
    .Q_N(_15962_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[20] ));
 sg13g2_dfrbp_1 _34366_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1199),
    .D(_01056_),
    .Q_N(_15961_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[21] ));
 sg13g2_dfrbp_1 _34367_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1197),
    .D(_01057_),
    .Q_N(_15960_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[22] ));
 sg13g2_dfrbp_1 _34368_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1195),
    .D(_01058_),
    .Q_N(_15959_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[23] ));
 sg13g2_dfrbp_1 _34369_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1193),
    .D(_01059_),
    .Q_N(_15958_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[24] ));
 sg13g2_dfrbp_1 _34370_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1191),
    .D(_01060_),
    .Q_N(_15957_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[25] ));
 sg13g2_dfrbp_1 _34371_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1189),
    .D(_01061_),
    .Q_N(_15956_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[26] ));
 sg13g2_dfrbp_1 _34372_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1187),
    .D(_01062_),
    .Q_N(_15955_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[27] ));
 sg13g2_dfrbp_1 _34373_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1185),
    .D(_01063_),
    .Q_N(_15954_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[28] ));
 sg13g2_dfrbp_1 _34374_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1183),
    .D(_01064_),
    .Q_N(_15953_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[29] ));
 sg13g2_dfrbp_1 _34375_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1181),
    .D(_01065_),
    .Q_N(_15952_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[30] ));
 sg13g2_dfrbp_1 _34376_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1179),
    .D(_01066_),
    .Q_N(_15951_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[31] ));
 sg13g2_dfrbp_1 _34377_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1177),
    .D(_01067_),
    .Q_N(_15950_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[3] ));
 sg13g2_dfrbp_1 _34378_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1175),
    .D(net4222),
    .Q_N(_15949_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[7] ));
 sg13g2_dfrbp_1 _34379_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1173),
    .D(_01069_),
    .Q_N(_15948_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[11] ));
 sg13g2_dfrbp_1 _34380_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1171),
    .D(_01070_),
    .Q_N(_15947_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[12] ));
 sg13g2_dfrbp_1 _34381_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1169),
    .D(net4560),
    .Q_N(_00240_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.privilege_mode[0] ));
 sg13g2_dfrbp_1 _34382_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1167),
    .D(_01072_),
    .Q_N(_00239_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.privilege_mode[1] ));
 sg13g2_dfrbp_1 _34383_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1165),
    .D(_01073_),
    .Q_N(_15946_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[3][0] ));
 sg13g2_dfrbp_1 _34384_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1164),
    .D(net4181),
    .Q_N(_15945_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[3][1] ));
 sg13g2_dfrbp_1 _34385_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1163),
    .D(_01075_),
    .Q_N(_15944_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[3][2] ));
 sg13g2_dfrbp_1 _34386_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1162),
    .D(net4159),
    .Q_N(_15943_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[3][3] ));
 sg13g2_dfrbp_1 _34387_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1161),
    .D(net4004),
    .Q_N(_15942_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[3][4] ));
 sg13g2_dfrbp_1 _34388_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1160),
    .D(_01078_),
    .Q_N(_15941_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[3][5] ));
 sg13g2_dfrbp_1 _34389_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1159),
    .D(net4208),
    .Q_N(_15940_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[3][6] ));
 sg13g2_dfrbp_1 _34390_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1158),
    .D(_01080_),
    .Q_N(_15939_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[3][7] ));
 sg13g2_dfrbp_1 _34391_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1157),
    .D(net2662),
    .Q_N(_15938_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[2][0] ));
 sg13g2_dfrbp_1 _34392_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1156),
    .D(net4097),
    .Q_N(_15937_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[2][1] ));
 sg13g2_dfrbp_1 _34393_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1155),
    .D(_01083_),
    .Q_N(_15936_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[2][2] ));
 sg13g2_dfrbp_1 _34394_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1154),
    .D(net4153),
    .Q_N(_15935_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[2][3] ));
 sg13g2_dfrbp_1 _34395_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1153),
    .D(net3989),
    .Q_N(_15934_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[2][4] ));
 sg13g2_dfrbp_1 _34396_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1152),
    .D(_01086_),
    .Q_N(_15933_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[2][5] ));
 sg13g2_dfrbp_1 _34397_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1151),
    .D(net4085),
    .Q_N(_15932_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[2][6] ));
 sg13g2_dfrbp_1 _34398_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1150),
    .D(_01088_),
    .Q_N(_15931_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[2][7] ));
 sg13g2_dfrbp_1 _34399_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1149),
    .D(_01089_),
    .Q_N(_15930_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[1][0] ));
 sg13g2_dfrbp_1 _34400_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1148),
    .D(net4035),
    .Q_N(_15929_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[1][1] ));
 sg13g2_dfrbp_1 _34401_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1147),
    .D(_01091_),
    .Q_N(_15928_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[1][2] ));
 sg13g2_dfrbp_1 _34402_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1146),
    .D(net4027),
    .Q_N(_15927_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[1][3] ));
 sg13g2_dfrbp_1 _34403_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1145),
    .D(net4095),
    .Q_N(_15926_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[1][4] ));
 sg13g2_dfrbp_1 _34404_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1144),
    .D(_01094_),
    .Q_N(_15925_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[1][5] ));
 sg13g2_dfrbp_1 _34405_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1143),
    .D(net4132),
    .Q_N(_15924_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[1][6] ));
 sg13g2_dfrbp_1 _34406_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1142),
    .D(_01096_),
    .Q_N(_15923_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[1][7] ));
 sg13g2_dfrbp_1 _34407_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1141),
    .D(net2761),
    .Q_N(_15922_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[15][0] ));
 sg13g2_dfrbp_1 _34408_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1140),
    .D(_01098_),
    .Q_N(_15921_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[15][1] ));
 sg13g2_dfrbp_1 _34409_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1139),
    .D(_01099_),
    .Q_N(_15920_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[15][2] ));
 sg13g2_dfrbp_1 _34410_ (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1138),
    .D(net4093),
    .Q_N(_15919_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[15][3] ));
 sg13g2_dfrbp_1 _34411_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1137),
    .D(net4090),
    .Q_N(_15918_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[15][4] ));
 sg13g2_dfrbp_1 _34412_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1136),
    .D(_01102_),
    .Q_N(_15917_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[15][5] ));
 sg13g2_dfrbp_1 _34413_ (.CLK(clknet_leaf_325_clk),
    .RESET_B(net1135),
    .D(_01103_),
    .Q_N(_15916_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[15][6] ));
 sg13g2_dfrbp_1 _34414_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1134),
    .D(net3975),
    .Q_N(_15915_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[15][7] ));
 sg13g2_dfrbp_1 _34415_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1133),
    .D(_01105_),
    .Q_N(_15914_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][0] ));
 sg13g2_dfrbp_1 _34416_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1132),
    .D(_01106_),
    .Q_N(_15913_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][1] ));
 sg13g2_dfrbp_1 _34417_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1131),
    .D(_01107_),
    .Q_N(_15912_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][2] ));
 sg13g2_dfrbp_1 _34418_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1130),
    .D(_01108_),
    .Q_N(_15911_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][3] ));
 sg13g2_dfrbp_1 _34419_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1129),
    .D(_01109_),
    .Q_N(_15910_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][4] ));
 sg13g2_dfrbp_1 _34420_ (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1128),
    .D(_01110_),
    .Q_N(_15909_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][5] ));
 sg13g2_dfrbp_1 _34421_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1127),
    .D(_01111_),
    .Q_N(_15908_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][6] ));
 sg13g2_dfrbp_1 _34422_ (.CLK(clknet_leaf_319_clk),
    .RESET_B(net1126),
    .D(_01112_),
    .Q_N(_15907_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][7] ));
 sg13g2_dfrbp_1 _34423_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1125),
    .D(_01113_),
    .Q_N(_15906_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][8] ));
 sg13g2_dfrbp_1 _34424_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1124),
    .D(_01114_),
    .Q_N(_15905_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][9] ));
 sg13g2_dfrbp_1 _34425_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1123),
    .D(_01115_),
    .Q_N(_15904_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][10] ));
 sg13g2_dfrbp_1 _34426_ (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1122),
    .D(_01116_),
    .Q_N(_15903_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][11] ));
 sg13g2_dfrbp_1 _34427_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1121),
    .D(_01117_),
    .Q_N(_15902_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][12] ));
 sg13g2_dfrbp_1 _34428_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1120),
    .D(_01118_),
    .Q_N(_15901_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][13] ));
 sg13g2_dfrbp_1 _34429_ (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1119),
    .D(_01119_),
    .Q_N(_15900_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][14] ));
 sg13g2_dfrbp_1 _34430_ (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1118),
    .D(_01120_),
    .Q_N(_15899_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][15] ));
 sg13g2_dfrbp_1 _34431_ (.CLK(clknet_leaf_320_clk),
    .RESET_B(net1117),
    .D(_01121_),
    .Q_N(_15898_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][16] ));
 sg13g2_dfrbp_1 _34432_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1116),
    .D(_01122_),
    .Q_N(_15897_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][17] ));
 sg13g2_dfrbp_1 _34433_ (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1115),
    .D(_01123_),
    .Q_N(_15896_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][18] ));
 sg13g2_dfrbp_1 _34434_ (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1114),
    .D(_01124_),
    .Q_N(_15895_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][19] ));
 sg13g2_dfrbp_1 _34435_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1113),
    .D(_01125_),
    .Q_N(_15894_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][20] ));
 sg13g2_dfrbp_1 _34436_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1112),
    .D(_01126_),
    .Q_N(_15893_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][21] ));
 sg13g2_dfrbp_1 _34437_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1111),
    .D(_01127_),
    .Q_N(_15892_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][22] ));
 sg13g2_dfrbp_1 _34438_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1110),
    .D(_01128_),
    .Q_N(_15891_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][23] ));
 sg13g2_dfrbp_1 _34439_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1109),
    .D(_01129_),
    .Q_N(_15890_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][24] ));
 sg13g2_dfrbp_1 _34440_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1108),
    .D(_01130_),
    .Q_N(_15889_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][25] ));
 sg13g2_dfrbp_1 _34441_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1107),
    .D(_01131_),
    .Q_N(_15888_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][26] ));
 sg13g2_dfrbp_1 _34442_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1106),
    .D(_01132_),
    .Q_N(_15887_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][27] ));
 sg13g2_dfrbp_1 _34443_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1105),
    .D(_01133_),
    .Q_N(_15886_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][28] ));
 sg13g2_dfrbp_1 _34444_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1104),
    .D(_01134_),
    .Q_N(_15885_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][29] ));
 sg13g2_dfrbp_1 _34445_ (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1103),
    .D(_01135_),
    .Q_N(_15884_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][30] ));
 sg13g2_dfrbp_1 _34446_ (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1102),
    .D(_01136_),
    .Q_N(_15883_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][31] ));
 sg13g2_dfrbp_1 _34447_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1101),
    .D(net2681),
    .Q_N(_00305_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[0] ));
 sg13g2_dfrbp_1 _34448_ (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1099),
    .D(_01138_),
    .Q_N(_15882_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[1] ));
 sg13g2_dfrbp_1 _34449_ (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1097),
    .D(net4130),
    .Q_N(_15881_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[2] ));
 sg13g2_dfrbp_1 _34450_ (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1095),
    .D(_01140_),
    .Q_N(_15880_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[3] ));
 sg13g2_dfrbp_1 _34451_ (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1093),
    .D(_01141_),
    .Q_N(_15879_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[4] ));
 sg13g2_dfrbp_1 _34452_ (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1091),
    .D(_01142_),
    .Q_N(_15878_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[5] ));
 sg13g2_dfrbp_1 _34453_ (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1089),
    .D(net5497),
    .Q_N(_15877_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[6] ));
 sg13g2_dfrbp_1 _34454_ (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1087),
    .D(_01144_),
    .Q_N(_15876_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[7] ));
 sg13g2_dfrbp_1 _34455_ (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1085),
    .D(_01145_),
    .Q_N(_15875_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[8] ));
 sg13g2_dfrbp_1 _34456_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1083),
    .D(net4116),
    .Q_N(_15874_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[9] ));
 sg13g2_dfrbp_1 _34457_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1081),
    .D(net3099),
    .Q_N(_15873_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[10] ));
 sg13g2_dfrbp_1 _34458_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1079),
    .D(_01148_),
    .Q_N(_15872_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[11] ));
 sg13g2_dfrbp_1 _34459_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1077),
    .D(_01149_),
    .Q_N(_15871_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[12] ));
 sg13g2_dfrbp_1 _34460_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1075),
    .D(net4485),
    .Q_N(_15870_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[13] ));
 sg13g2_dfrbp_1 _34461_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1073),
    .D(_01151_),
    .Q_N(_15869_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[14] ));
 sg13g2_dfrbp_1 _34462_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1071),
    .D(_01152_),
    .Q_N(_15868_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[15] ));
 sg13g2_dfrbp_1 _34463_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1069),
    .D(_01153_),
    .Q_N(_15867_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[16] ));
 sg13g2_dfrbp_1 _34464_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1067),
    .D(_01154_),
    .Q_N(_15866_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[17] ));
 sg13g2_dfrbp_1 _34465_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1065),
    .D(_01155_),
    .Q_N(_15865_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[18] ));
 sg13g2_dfrbp_1 _34466_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1063),
    .D(_01156_),
    .Q_N(_15864_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[19] ));
 sg13g2_dfrbp_1 _34467_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1061),
    .D(_01157_),
    .Q_N(_15863_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[20] ));
 sg13g2_dfrbp_1 _34468_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1059),
    .D(_01158_),
    .Q_N(_15862_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[21] ));
 sg13g2_dfrbp_1 _34469_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1057),
    .D(_01159_),
    .Q_N(_15861_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[22] ));
 sg13g2_dfrbp_1 _34470_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1055),
    .D(_01160_),
    .Q_N(_15860_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[23] ));
 sg13g2_dfrbp_1 _34471_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1053),
    .D(_01161_),
    .Q_N(_15859_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[24] ));
 sg13g2_dfrbp_1 _34472_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1051),
    .D(_01162_),
    .Q_N(_15858_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[25] ));
 sg13g2_dfrbp_1 _34473_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1049),
    .D(_01163_),
    .Q_N(_15857_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[26] ));
 sg13g2_dfrbp_1 _34474_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1047),
    .D(_01164_),
    .Q_N(_15856_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[27] ));
 sg13g2_dfrbp_1 _34475_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1045),
    .D(_01165_),
    .Q_N(_15855_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[28] ));
 sg13g2_dfrbp_1 _34476_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1043),
    .D(net4476),
    .Q_N(_15854_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[29] ));
 sg13g2_dfrbp_1 _34477_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1041),
    .D(_01167_),
    .Q_N(_15853_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[30] ));
 sg13g2_dfrbp_1 _34478_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1039),
    .D(_01168_),
    .Q_N(_15852_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[31] ));
 sg13g2_dfrbp_1 _34479_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1037),
    .D(_01169_),
    .Q_N(_15851_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[32] ));
 sg13g2_dfrbp_1 _34480_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1035),
    .D(_01170_),
    .Q_N(_15850_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[33] ));
 sg13g2_dfrbp_1 _34481_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1033),
    .D(net5342),
    .Q_N(_15849_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[34] ));
 sg13g2_dfrbp_1 _34482_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1031),
    .D(_01172_),
    .Q_N(_15848_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[35] ));
 sg13g2_dfrbp_1 _34483_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1029),
    .D(_01173_),
    .Q_N(_15847_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[36] ));
 sg13g2_dfrbp_1 _34484_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1027),
    .D(_01174_),
    .Q_N(_15846_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[37] ));
 sg13g2_dfrbp_1 _34485_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1025),
    .D(_01175_),
    .Q_N(_15845_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[38] ));
 sg13g2_dfrbp_1 _34486_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1023),
    .D(_01176_),
    .Q_N(_15844_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[39] ));
 sg13g2_dfrbp_1 _34487_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1021),
    .D(_01177_),
    .Q_N(_15843_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[40] ));
 sg13g2_dfrbp_1 _34488_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1019),
    .D(_01178_),
    .Q_N(_15842_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[41] ));
 sg13g2_dfrbp_1 _34489_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1017),
    .D(net5345),
    .Q_N(_15841_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[42] ));
 sg13g2_dfrbp_1 _34490_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1015),
    .D(net4060),
    .Q_N(_15840_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[43] ));
 sg13g2_dfrbp_1 _34491_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1013),
    .D(_01181_),
    .Q_N(_15839_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[44] ));
 sg13g2_dfrbp_1 _34492_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1011),
    .D(_01182_),
    .Q_N(_15838_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[45] ));
 sg13g2_dfrbp_1 _34493_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1009),
    .D(_01183_),
    .Q_N(_15837_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[46] ));
 sg13g2_dfrbp_1 _34494_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1007),
    .D(net5480),
    .Q_N(_15836_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[47] ));
 sg13g2_dfrbp_1 _34495_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1005),
    .D(net3792),
    .Q_N(_15835_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[48] ));
 sg13g2_dfrbp_1 _34496_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1003),
    .D(_01186_),
    .Q_N(_15834_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[49] ));
 sg13g2_dfrbp_1 _34497_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1001),
    .D(_01187_),
    .Q_N(_15833_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[50] ));
 sg13g2_dfrbp_1 _34498_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net999),
    .D(_01188_),
    .Q_N(_15832_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[51] ));
 sg13g2_dfrbp_1 _34499_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net997),
    .D(net5094),
    .Q_N(_15831_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[52] ));
 sg13g2_dfrbp_1 _34500_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net995),
    .D(_01190_),
    .Q_N(_15830_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[53] ));
 sg13g2_dfrbp_1 _34501_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net993),
    .D(net4649),
    .Q_N(_15829_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[54] ));
 sg13g2_dfrbp_1 _34502_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net991),
    .D(_01192_),
    .Q_N(_15828_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[55] ));
 sg13g2_dfrbp_1 _34503_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net989),
    .D(net4512),
    .Q_N(_15827_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[56] ));
 sg13g2_dfrbp_1 _34504_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net987),
    .D(_01194_),
    .Q_N(_15826_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[57] ));
 sg13g2_dfrbp_1 _34505_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net985),
    .D(_01195_),
    .Q_N(_15825_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[58] ));
 sg13g2_dfrbp_1 _34506_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net983),
    .D(net4960),
    .Q_N(_15824_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[59] ));
 sg13g2_dfrbp_1 _34507_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net981),
    .D(_01197_),
    .Q_N(_15823_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[60] ));
 sg13g2_dfrbp_1 _34508_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net979),
    .D(_01198_),
    .Q_N(_15822_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[61] ));
 sg13g2_dfrbp_1 _34509_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net977),
    .D(net3194),
    .Q_N(_15821_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[62] ));
 sg13g2_dfrbp_1 _34510_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net975),
    .D(net4029),
    .Q_N(_15820_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[63] ));
 sg13g2_dfrbp_1 _34511_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net973),
    .D(_01201_),
    .Q_N(_15819_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[0] ));
 sg13g2_dfrbp_1 _34512_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net971),
    .D(_01202_),
    .Q_N(_15818_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[1] ));
 sg13g2_dfrbp_1 _34513_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net969),
    .D(net5403),
    .Q_N(_15817_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[2] ));
 sg13g2_dfrbp_1 _34514_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net967),
    .D(net5326),
    .Q_N(_15816_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[3] ));
 sg13g2_dfrbp_1 _34515_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net965),
    .D(net5291),
    .Q_N(_15815_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[4] ));
 sg13g2_dfrbp_1 _34516_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net963),
    .D(net5448),
    .Q_N(_15814_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[5] ));
 sg13g2_dfrbp_1 _34517_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net961),
    .D(net5257),
    .Q_N(_15813_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[6] ));
 sg13g2_dfrbp_1 _34518_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net959),
    .D(net5284),
    .Q_N(_15812_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[7] ));
 sg13g2_dfrbp_1 _34519_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net957),
    .D(net5231),
    .Q_N(_15811_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[8] ));
 sg13g2_dfrbp_1 _34520_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net955),
    .D(_01210_),
    .Q_N(_15810_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[9] ));
 sg13g2_dfrbp_1 _34521_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net953),
    .D(net5225),
    .Q_N(_15809_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[10] ));
 sg13g2_dfrbp_1 _34522_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net951),
    .D(_01212_),
    .Q_N(_15808_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[11] ));
 sg13g2_dfrbp_1 _34523_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net949),
    .D(_01213_),
    .Q_N(_15807_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[12] ));
 sg13g2_dfrbp_1 _34524_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net947),
    .D(_01214_),
    .Q_N(_15806_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[13] ));
 sg13g2_dfrbp_1 _34525_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net945),
    .D(_01215_),
    .Q_N(_15805_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[14] ));
 sg13g2_dfrbp_1 _34526_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net943),
    .D(_01216_),
    .Q_N(_15804_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[15] ));
 sg13g2_dfrbp_1 _34527_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net941),
    .D(net5306),
    .Q_N(_15803_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[16] ));
 sg13g2_dfrbp_1 _34528_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net939),
    .D(_01218_),
    .Q_N(_15802_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[17] ));
 sg13g2_dfrbp_1 _34529_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net937),
    .D(_01219_),
    .Q_N(_15801_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[18] ));
 sg13g2_dfrbp_1 _34530_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net935),
    .D(net5213),
    .Q_N(_15800_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[19] ));
 sg13g2_dfrbp_1 _34531_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net933),
    .D(net5464),
    .Q_N(_15799_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[20] ));
 sg13g2_dfrbp_1 _34532_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net931),
    .D(net5393),
    .Q_N(_15798_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[21] ));
 sg13g2_dfrbp_1 _34533_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net929),
    .D(net5249),
    .Q_N(_15797_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[22] ));
 sg13g2_dfrbp_1 _34534_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net927),
    .D(_01224_),
    .Q_N(_15796_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[23] ));
 sg13g2_dfrbp_1 _34535_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net925),
    .D(net5374),
    .Q_N(_15795_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[24] ));
 sg13g2_dfrbp_1 _34536_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net923),
    .D(net5316),
    .Q_N(_15794_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[25] ));
 sg13g2_dfrbp_1 _34537_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net921),
    .D(net5505),
    .Q_N(_15793_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[26] ));
 sg13g2_dfrbp_1 _34538_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net919),
    .D(_01228_),
    .Q_N(_15792_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[27] ));
 sg13g2_dfrbp_1 _34539_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net917),
    .D(net5223),
    .Q_N(_15791_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[28] ));
 sg13g2_dfrbp_1 _34540_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net915),
    .D(net5410),
    .Q_N(_15790_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[29] ));
 sg13g2_dfrbp_1 _34541_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net913),
    .D(net5262),
    .Q_N(_15789_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[30] ));
 sg13g2_dfrbp_1 _34542_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net911),
    .D(_01232_),
    .Q_N(_15788_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[31] ));
 sg13g2_dfrbp_1 _34543_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net909),
    .D(_01233_),
    .Q_N(_15787_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[0] ));
 sg13g2_dfrbp_1 _34544_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net907),
    .D(_01234_),
    .Q_N(_00183_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[1] ));
 sg13g2_dfrbp_1 _34545_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net905),
    .D(_01235_),
    .Q_N(_15786_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[2] ));
 sg13g2_dfrbp_1 _34546_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net903),
    .D(_01236_),
    .Q_N(_00182_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[3] ));
 sg13g2_dfrbp_1 _34547_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net901),
    .D(_01237_),
    .Q_N(_00181_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[4] ));
 sg13g2_dfrbp_1 _34548_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net899),
    .D(_01238_),
    .Q_N(_00180_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[5] ));
 sg13g2_dfrbp_1 _34549_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net897),
    .D(_01239_),
    .Q_N(_15785_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[6] ));
 sg13g2_dfrbp_1 _34550_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net895),
    .D(_01240_),
    .Q_N(_00179_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[7] ));
 sg13g2_dfrbp_1 _34551_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net893),
    .D(_01241_),
    .Q_N(_00178_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[8] ));
 sg13g2_dfrbp_1 _34552_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net891),
    .D(_01242_),
    .Q_N(_00177_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[9] ));
 sg13g2_dfrbp_1 _34553_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net889),
    .D(_01243_),
    .Q_N(_00176_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[10] ));
 sg13g2_dfrbp_1 _34554_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net887),
    .D(_01244_),
    .Q_N(_00175_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[11] ));
 sg13g2_dfrbp_1 _34555_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net885),
    .D(_01245_),
    .Q_N(_00174_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[12] ));
 sg13g2_dfrbp_1 _34556_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net883),
    .D(_01246_),
    .Q_N(_00173_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[13] ));
 sg13g2_dfrbp_1 _34557_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net881),
    .D(_01247_),
    .Q_N(_15784_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[14] ));
 sg13g2_dfrbp_1 _34558_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net879),
    .D(_01248_),
    .Q_N(_00172_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[15] ));
 sg13g2_dfrbp_1 _34559_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net877),
    .D(_01249_),
    .Q_N(_00171_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[16] ));
 sg13g2_dfrbp_1 _34560_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net875),
    .D(_01250_),
    .Q_N(_00170_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[17] ));
 sg13g2_dfrbp_1 _34561_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net873),
    .D(_01251_),
    .Q_N(_00169_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[18] ));
 sg13g2_dfrbp_1 _34562_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net871),
    .D(_01252_),
    .Q_N(_00168_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[19] ));
 sg13g2_dfrbp_1 _34563_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net869),
    .D(_01253_),
    .Q_N(_00167_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[20] ));
 sg13g2_dfrbp_1 _34564_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net867),
    .D(_01254_),
    .Q_N(_00166_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[21] ));
 sg13g2_dfrbp_1 _34565_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net865),
    .D(_01255_),
    .Q_N(_00165_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[22] ));
 sg13g2_dfrbp_1 _34566_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net863),
    .D(_01256_),
    .Q_N(_00164_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[23] ));
 sg13g2_dfrbp_1 _34567_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net861),
    .D(net5187),
    .Q_N(_00163_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[24] ));
 sg13g2_dfrbp_1 _34568_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net859),
    .D(_01258_),
    .Q_N(_00162_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[25] ));
 sg13g2_dfrbp_1 _34569_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net857),
    .D(_01259_),
    .Q_N(_00161_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[26] ));
 sg13g2_dfrbp_1 _34570_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net855),
    .D(_01260_),
    .Q_N(_00160_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[27] ));
 sg13g2_dfrbp_1 _34571_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net853),
    .D(_01261_),
    .Q_N(_00159_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[28] ));
 sg13g2_dfrbp_1 _34572_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net851),
    .D(_01262_),
    .Q_N(_00158_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[29] ));
 sg13g2_dfrbp_1 _34573_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net849),
    .D(_01263_),
    .Q_N(_15783_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[30] ));
 sg13g2_dfrbp_1 _34574_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net847),
    .D(_01264_),
    .Q_N(_15782_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[31] ));
 sg13g2_dfrbp_1 _34575_ (.CLK(clknet_leaf_289_clk),
    .RESET_B(net845),
    .D(_01265_),
    .Q_N(_00304_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[0] ));
 sg13g2_dfrbp_1 _34576_ (.CLK(clknet_leaf_289_clk),
    .RESET_B(net844),
    .D(net4285),
    .Q_N(_15781_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[1] ));
 sg13g2_dfrbp_1 _34577_ (.CLK(clknet_leaf_290_clk),
    .RESET_B(net843),
    .D(net3461),
    .Q_N(_15780_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[2] ));
 sg13g2_dfrbp_1 _34578_ (.CLK(clknet_leaf_282_clk),
    .RESET_B(net842),
    .D(_01268_),
    .Q_N(_15779_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[3] ));
 sg13g2_dfrbp_1 _34579_ (.CLK(clknet_leaf_286_clk),
    .RESET_B(net841),
    .D(_01269_),
    .Q_N(_15778_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[4] ));
 sg13g2_dfrbp_1 _34580_ (.CLK(clknet_leaf_287_clk),
    .RESET_B(net840),
    .D(_01270_),
    .Q_N(_15777_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[5] ));
 sg13g2_dfrbp_1 _34581_ (.CLK(clknet_leaf_286_clk),
    .RESET_B(net839),
    .D(_01271_),
    .Q_N(_15776_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[6] ));
 sg13g2_dfrbp_1 _34582_ (.CLK(clknet_leaf_283_clk),
    .RESET_B(net838),
    .D(_01272_),
    .Q_N(_15775_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[7] ));
 sg13g2_dfrbp_1 _34583_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net837),
    .D(_01273_),
    .Q_N(_15774_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[8] ));
 sg13g2_dfrbp_1 _34584_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net836),
    .D(_01274_),
    .Q_N(_15773_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[9] ));
 sg13g2_dfrbp_1 _34585_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net835),
    .D(net3366),
    .Q_N(_15772_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[10] ));
 sg13g2_dfrbp_1 _34586_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net834),
    .D(_01276_),
    .Q_N(_15771_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[11] ));
 sg13g2_dfrbp_1 _34587_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net833),
    .D(net3797),
    .Q_N(_15770_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[12] ));
 sg13g2_dfrbp_1 _34588_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net832),
    .D(_01278_),
    .Q_N(_15769_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[13] ));
 sg13g2_dfrbp_1 _34589_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net831),
    .D(_01279_),
    .Q_N(_15768_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[14] ));
 sg13g2_dfrbp_1 _34590_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net830),
    .D(_01280_),
    .Q_N(_15767_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[15] ));
 sg13g2_dfrbp_1 _34591_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net829),
    .D(net3421),
    .Q_N(_15766_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[16] ));
 sg13g2_dfrbp_1 _34592_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net828),
    .D(_01282_),
    .Q_N(_15765_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[17] ));
 sg13g2_dfrbp_1 _34593_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net827),
    .D(net3935),
    .Q_N(_15764_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[18] ));
 sg13g2_dfrbp_1 _34594_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net826),
    .D(_01284_),
    .Q_N(_15763_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[19] ));
 sg13g2_dfrbp_1 _34595_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net825),
    .D(_01285_),
    .Q_N(_15762_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[20] ));
 sg13g2_dfrbp_1 _34596_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net824),
    .D(_01286_),
    .Q_N(_15761_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[21] ));
 sg13g2_dfrbp_1 _34597_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net823),
    .D(_01287_),
    .Q_N(_15760_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[22] ));
 sg13g2_dfrbp_1 _34598_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net822),
    .D(_01288_),
    .Q_N(_15759_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[23] ));
 sg13g2_dfrbp_1 _34599_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net821),
    .D(net3762),
    .Q_N(_15758_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[24] ));
 sg13g2_dfrbp_1 _34600_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net820),
    .D(_01290_),
    .Q_N(_15757_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[25] ));
 sg13g2_dfrbp_1 _34601_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net819),
    .D(_01291_),
    .Q_N(_15756_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[26] ));
 sg13g2_dfrbp_1 _34602_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net818),
    .D(_01292_),
    .Q_N(_15755_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[27] ));
 sg13g2_dfrbp_1 _34603_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net817),
    .D(net2830),
    .Q_N(_15754_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[28] ));
 sg13g2_dfrbp_1 _34604_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net816),
    .D(_01294_),
    .Q_N(_15753_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[29] ));
 sg13g2_dfrbp_1 _34605_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net815),
    .D(net3256),
    .Q_N(_15752_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[30] ));
 sg13g2_dfrbp_1 _34606_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net814),
    .D(_01296_),
    .Q_N(_15751_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[31] ));
 sg13g2_dfrbp_1 _34607_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net813),
    .D(_01297_),
    .Q_N(_15750_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[32] ));
 sg13g2_dfrbp_1 _34608_ (.CLK(clknet_leaf_281_clk),
    .RESET_B(net812),
    .D(_01298_),
    .Q_N(_15749_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[33] ));
 sg13g2_dfrbp_1 _34609_ (.CLK(clknet_leaf_281_clk),
    .RESET_B(net811),
    .D(net3690),
    .Q_N(_15748_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[34] ));
 sg13g2_dfrbp_1 _34610_ (.CLK(clknet_leaf_282_clk),
    .RESET_B(net810),
    .D(_01300_),
    .Q_N(_15747_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[35] ));
 sg13g2_dfrbp_1 _34611_ (.CLK(clknet_leaf_282_clk),
    .RESET_B(net809),
    .D(net4345),
    .Q_N(_15746_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[36] ));
 sg13g2_dfrbp_1 _34612_ (.CLK(clknet_leaf_286_clk),
    .RESET_B(net808),
    .D(_01302_),
    .Q_N(_15745_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[37] ));
 sg13g2_dfrbp_1 _34613_ (.CLK(clknet_leaf_283_clk),
    .RESET_B(net807),
    .D(_01303_),
    .Q_N(_15744_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[38] ));
 sg13g2_dfrbp_1 _34614_ (.CLK(clknet_leaf_283_clk),
    .RESET_B(net806),
    .D(_01304_),
    .Q_N(_15743_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[39] ));
 sg13g2_dfrbp_1 _34615_ (.CLK(clknet_leaf_283_clk),
    .RESET_B(net805),
    .D(_01305_),
    .Q_N(_15742_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[40] ));
 sg13g2_dfrbp_1 _34616_ (.CLK(clknet_leaf_283_clk),
    .RESET_B(net804),
    .D(_01306_),
    .Q_N(_15741_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[41] ));
 sg13g2_dfrbp_1 _34617_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net803),
    .D(net3712),
    .Q_N(_15740_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[42] ));
 sg13g2_dfrbp_1 _34618_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net802),
    .D(_01308_),
    .Q_N(_15739_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[43] ));
 sg13g2_dfrbp_1 _34619_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net801),
    .D(_01309_),
    .Q_N(_15738_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[44] ));
 sg13g2_dfrbp_1 _34620_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net800),
    .D(_01310_),
    .Q_N(_15737_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[45] ));
 sg13g2_dfrbp_1 _34621_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net799),
    .D(net3311),
    .Q_N(_15736_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[46] ));
 sg13g2_dfrbp_1 _34622_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net798),
    .D(_01312_),
    .Q_N(_15735_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[47] ));
 sg13g2_dfrbp_1 _34623_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net797),
    .D(net3776),
    .Q_N(_15734_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[48] ));
 sg13g2_dfrbp_1 _34624_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net796),
    .D(_01314_),
    .Q_N(_15733_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[49] ));
 sg13g2_dfrbp_1 _34625_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net795),
    .D(_01315_),
    .Q_N(_15732_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[50] ));
 sg13g2_dfrbp_1 _34626_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net794),
    .D(_01316_),
    .Q_N(_15731_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[51] ));
 sg13g2_dfrbp_1 _34627_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net793),
    .D(net3486),
    .Q_N(_15730_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[52] ));
 sg13g2_dfrbp_1 _34628_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net792),
    .D(_01318_),
    .Q_N(_15729_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[53] ));
 sg13g2_dfrbp_1 _34629_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net791),
    .D(_01319_),
    .Q_N(_15728_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[54] ));
 sg13g2_dfrbp_1 _34630_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net790),
    .D(_01320_),
    .Q_N(_15727_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[55] ));
 sg13g2_dfrbp_1 _34631_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net789),
    .D(_01321_),
    .Q_N(_15726_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[56] ));
 sg13g2_dfrbp_1 _34632_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net788),
    .D(_01322_),
    .Q_N(_15725_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[57] ));
 sg13g2_dfrbp_1 _34633_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net787),
    .D(net3207),
    .Q_N(_15724_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[58] ));
 sg13g2_dfrbp_1 _34634_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net786),
    .D(_01324_),
    .Q_N(_15723_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[59] ));
 sg13g2_dfrbp_1 _34635_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net785),
    .D(_01325_),
    .Q_N(_15722_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[60] ));
 sg13g2_dfrbp_1 _34636_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net784),
    .D(_01326_),
    .Q_N(_15721_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[61] ));
 sg13g2_dfrbp_1 _34637_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net783),
    .D(_01327_),
    .Q_N(_15720_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[62] ));
 sg13g2_dfrbp_1 _34638_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net782),
    .D(net3671),
    .Q_N(_15719_),
    .Q(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[63] ));
 sg13g2_dfrbp_1 _34639_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net781),
    .D(_01329_),
    .Q_N(_15718_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.bit_idx[0] ));
 sg13g2_dfrbp_1 _34640_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net779),
    .D(_01330_),
    .Q_N(_15717_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.bit_idx[1] ));
 sg13g2_dfrbp_1 _34641_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net777),
    .D(net3979),
    .Q_N(_15716_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.bit_idx[2] ));
 sg13g2_dfrbp_1 _34642_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net775),
    .D(_01332_),
    .Q_N(_15715_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.bit_idx[3] ));
 sg13g2_dfrbp_1 _34643_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net773),
    .D(net4299),
    .Q_N(_00283_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.bit_idx[4] ));
 sg13g2_dfrbp_1 _34644_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net771),
    .D(_01334_),
    .Q_N(_15714_),
    .Q(\soc_I.kianv_I.control_unit_I.div_ready ));
 sg13g2_dfrbp_1 _34645_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net769),
    .D(_01335_),
    .Q_N(_15713_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[0] ));
 sg13g2_dfrbp_1 _34646_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net768),
    .D(_01336_),
    .Q_N(_15712_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[1] ));
 sg13g2_dfrbp_1 _34647_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net767),
    .D(_01337_),
    .Q_N(_15711_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[2] ));
 sg13g2_dfrbp_1 _34648_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net766),
    .D(_01338_),
    .Q_N(_15710_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[3] ));
 sg13g2_dfrbp_1 _34649_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net765),
    .D(_01339_),
    .Q_N(_15709_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[4] ));
 sg13g2_dfrbp_1 _34650_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net764),
    .D(_01340_),
    .Q_N(_15708_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[5] ));
 sg13g2_dfrbp_1 _34651_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net763),
    .D(_01341_),
    .Q_N(_15707_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[6] ));
 sg13g2_dfrbp_1 _34652_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net762),
    .D(_01342_),
    .Q_N(_15706_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[7] ));
 sg13g2_dfrbp_1 _34653_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net761),
    .D(_01343_),
    .Q_N(_15705_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[8] ));
 sg13g2_dfrbp_1 _34654_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net760),
    .D(_01344_),
    .Q_N(_15704_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[9] ));
 sg13g2_dfrbp_1 _34655_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net759),
    .D(_01345_),
    .Q_N(_15703_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[10] ));
 sg13g2_dfrbp_1 _34656_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net758),
    .D(_01346_),
    .Q_N(_15702_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[11] ));
 sg13g2_dfrbp_1 _34657_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net757),
    .D(_01347_),
    .Q_N(_15701_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[12] ));
 sg13g2_dfrbp_1 _34658_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net756),
    .D(_01348_),
    .Q_N(_15700_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[13] ));
 sg13g2_dfrbp_1 _34659_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net755),
    .D(_01349_),
    .Q_N(_15699_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[14] ));
 sg13g2_dfrbp_1 _34660_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net754),
    .D(_01350_),
    .Q_N(_15698_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[15] ));
 sg13g2_dfrbp_1 _34661_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net753),
    .D(_01351_),
    .Q_N(_15697_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[16] ));
 sg13g2_dfrbp_1 _34662_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net752),
    .D(_01352_),
    .Q_N(_15696_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[17] ));
 sg13g2_dfrbp_1 _34663_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net751),
    .D(_01353_),
    .Q_N(_15695_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[18] ));
 sg13g2_dfrbp_1 _34664_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net750),
    .D(_01354_),
    .Q_N(_15694_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[19] ));
 sg13g2_dfrbp_1 _34665_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net749),
    .D(_01355_),
    .Q_N(_15693_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[20] ));
 sg13g2_dfrbp_1 _34666_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net748),
    .D(_01356_),
    .Q_N(_15692_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[21] ));
 sg13g2_dfrbp_1 _34667_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net747),
    .D(_01357_),
    .Q_N(_15691_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[22] ));
 sg13g2_dfrbp_1 _34668_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net746),
    .D(_01358_),
    .Q_N(_15690_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[23] ));
 sg13g2_dfrbp_1 _34669_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net745),
    .D(_01359_),
    .Q_N(_15689_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[24] ));
 sg13g2_dfrbp_1 _34670_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net744),
    .D(_01360_),
    .Q_N(_15688_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[25] ));
 sg13g2_dfrbp_1 _34671_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net743),
    .D(_01361_),
    .Q_N(_15687_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[26] ));
 sg13g2_dfrbp_1 _34672_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net742),
    .D(_01362_),
    .Q_N(_15686_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[27] ));
 sg13g2_dfrbp_1 _34673_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net741),
    .D(_01363_),
    .Q_N(_15685_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[28] ));
 sg13g2_dfrbp_1 _34674_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net740),
    .D(_01364_),
    .Q_N(_15684_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[29] ));
 sg13g2_dfrbp_1 _34675_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net739),
    .D(_01365_),
    .Q_N(_15683_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[30] ));
 sg13g2_dfrbp_1 _34676_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net738),
    .D(_01366_),
    .Q_N(_15682_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[31] ));
 sg13g2_dfrbp_1 _34677_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net737),
    .D(_01367_),
    .Q_N(_00252_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.state[0] ));
 sg13g2_dfrbp_1 _34678_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net736),
    .D(_01368_),
    .Q_N(_15681_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.bit_idx[0] ));
 sg13g2_dfrbp_1 _34679_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net734),
    .D(_01369_),
    .Q_N(_00256_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.bit_idx[1] ));
 sg13g2_dfrbp_1 _34680_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net732),
    .D(net5519),
    .Q_N(_00255_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.bit_idx[2] ));
 sg13g2_dfrbp_1 _34681_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net730),
    .D(net5470),
    .Q_N(_00254_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.bit_idx[3] ));
 sg13g2_dfrbp_1 _34682_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net728),
    .D(_01372_),
    .Q_N(_00251_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.bit_idx[4] ));
 sg13g2_dfrbp_1 _34683_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net726),
    .D(_01373_),
    .Q_N(_00284_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_state[0] ));
 sg13g2_dfrbp_1 _34684_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net725),
    .D(_01374_),
    .Q_N(_15680_),
    .Q(\soc_I.kianv_I.control_unit_I.mul_ready ));
 sg13g2_dfrbp_1 _34685_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net723),
    .D(_01375_),
    .Q_N(_00208_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[0] ));
 sg13g2_dfrbp_1 _34686_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net721),
    .D(_01376_),
    .Q_N(_00204_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[1] ));
 sg13g2_dfrbp_1 _34687_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net719),
    .D(_01377_),
    .Q_N(_00200_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[2] ));
 sg13g2_dfrbp_1 _34688_ (.CLK(clknet_leaf_271_clk),
    .RESET_B(net717),
    .D(_01378_),
    .Q_N(_15679_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[3] ));
 sg13g2_dfrbp_1 _34689_ (.CLK(clknet_leaf_271_clk),
    .RESET_B(net715),
    .D(_01379_),
    .Q_N(_00196_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[4] ));
 sg13g2_dfrbp_1 _34690_ (.CLK(clknet_leaf_270_clk),
    .RESET_B(net713),
    .D(_01380_),
    .Q_N(_00192_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[5] ));
 sg13g2_dfrbp_1 _34691_ (.CLK(clknet_leaf_270_clk),
    .RESET_B(net711),
    .D(_01381_),
    .Q_N(_00186_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[6] ));
 sg13g2_dfrbp_1 _34692_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net709),
    .D(_01382_),
    .Q_N(_15678_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[7] ));
 sg13g2_dfrbp_1 _34693_ (.CLK(clknet_leaf_270_clk),
    .RESET_B(net707),
    .D(_01383_),
    .Q_N(_00210_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[8] ));
 sg13g2_dfrbp_1 _34694_ (.CLK(clknet_leaf_271_clk),
    .RESET_B(net705),
    .D(_01384_),
    .Q_N(_00206_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[9] ));
 sg13g2_dfrbp_1 _34695_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net703),
    .D(_01385_),
    .Q_N(_00202_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[10] ));
 sg13g2_dfrbp_1 _34696_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net701),
    .D(_01386_),
    .Q_N(_15677_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[11] ));
 sg13g2_dfrbp_1 _34697_ (.CLK(clknet_leaf_271_clk),
    .RESET_B(net699),
    .D(_01387_),
    .Q_N(_00198_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[12] ));
 sg13g2_dfrbp_1 _34698_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net697),
    .D(_01388_),
    .Q_N(_00194_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[13] ));
 sg13g2_dfrbp_1 _34699_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net695),
    .D(_01389_),
    .Q_N(_00190_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[14] ));
 sg13g2_dfrbp_1 _34700_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net693),
    .D(_01390_),
    .Q_N(_15676_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[15] ));
 sg13g2_dfrbp_1 _34701_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net691),
    .D(_01391_),
    .Q_N(_15675_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[16] ));
 sg13g2_dfrbp_1 _34702_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net689),
    .D(_01392_),
    .Q_N(_15674_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[17] ));
 sg13g2_dfrbp_1 _34703_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net687),
    .D(_01393_),
    .Q_N(_15673_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[18] ));
 sg13g2_dfrbp_1 _34704_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net685),
    .D(_01394_),
    .Q_N(_15672_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[19] ));
 sg13g2_dfrbp_1 _34705_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net683),
    .D(_01395_),
    .Q_N(_15671_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[20] ));
 sg13g2_dfrbp_1 _34706_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net681),
    .D(_01396_),
    .Q_N(_15670_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[21] ));
 sg13g2_dfrbp_1 _34707_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net679),
    .D(_01397_),
    .Q_N(_15669_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[22] ));
 sg13g2_dfrbp_1 _34708_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net677),
    .D(_01398_),
    .Q_N(_15668_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[23] ));
 sg13g2_dfrbp_1 _34709_ (.CLK(clknet_leaf_271_clk),
    .RESET_B(net675),
    .D(_01399_),
    .Q_N(_15667_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[24] ));
 sg13g2_dfrbp_1 _34710_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net673),
    .D(_01400_),
    .Q_N(_15666_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[25] ));
 sg13g2_dfrbp_1 _34711_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net671),
    .D(_01401_),
    .Q_N(_15665_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[26] ));
 sg13g2_dfrbp_1 _34712_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net669),
    .D(_01402_),
    .Q_N(_15664_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[27] ));
 sg13g2_dfrbp_1 _34713_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net667),
    .D(_01403_),
    .Q_N(_15663_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[28] ));
 sg13g2_dfrbp_1 _34714_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net665),
    .D(_01404_),
    .Q_N(_15662_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[29] ));
 sg13g2_dfrbp_1 _34715_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net663),
    .D(_01405_),
    .Q_N(_15661_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[30] ));
 sg13g2_dfrbp_1 _34716_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net661),
    .D(_01406_),
    .Q_N(_15660_),
    .Q(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[31] ));
 sg13g2_dfrbp_1 _34717_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net659),
    .D(_01407_),
    .Q_N(_15659_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[0] ));
 sg13g2_dfrbp_1 _34718_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net657),
    .D(_01408_),
    .Q_N(_15658_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[1] ));
 sg13g2_dfrbp_1 _34719_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net655),
    .D(_01409_),
    .Q_N(_15657_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[2] ));
 sg13g2_dfrbp_1 _34720_ (.CLK(clknet_leaf_268_clk),
    .RESET_B(net653),
    .D(_01410_),
    .Q_N(_15656_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[3] ));
 sg13g2_dfrbp_1 _34721_ (.CLK(clknet_leaf_264_clk),
    .RESET_B(net651),
    .D(_01411_),
    .Q_N(_15655_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[4] ));
 sg13g2_dfrbp_1 _34722_ (.CLK(clknet_leaf_265_clk),
    .RESET_B(net649),
    .D(_01412_),
    .Q_N(_15654_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[5] ));
 sg13g2_dfrbp_1 _34723_ (.CLK(clknet_leaf_268_clk),
    .RESET_B(net647),
    .D(_01413_),
    .Q_N(_15653_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[6] ));
 sg13g2_dfrbp_1 _34724_ (.CLK(clknet_leaf_267_clk),
    .RESET_B(net645),
    .D(_01414_),
    .Q_N(_15652_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[7] ));
 sg13g2_dfrbp_1 _34725_ (.CLK(clknet_leaf_266_clk),
    .RESET_B(net643),
    .D(_01415_),
    .Q_N(_15651_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[8] ));
 sg13g2_dfrbp_1 _34726_ (.CLK(clknet_leaf_267_clk),
    .RESET_B(net641),
    .D(_01416_),
    .Q_N(_15650_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[9] ));
 sg13g2_dfrbp_1 _34727_ (.CLK(clknet_leaf_270_clk),
    .RESET_B(net639),
    .D(_01417_),
    .Q_N(_15649_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[10] ));
 sg13g2_dfrbp_1 _34728_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net637),
    .D(_01418_),
    .Q_N(_15648_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[11] ));
 sg13g2_dfrbp_1 _34729_ (.CLK(clknet_leaf_263_clk),
    .RESET_B(net635),
    .D(_01419_),
    .Q_N(_15647_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[12] ));
 sg13g2_dfrbp_1 _34730_ (.CLK(clknet_leaf_268_clk),
    .RESET_B(net633),
    .D(_01420_),
    .Q_N(_15646_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[13] ));
 sg13g2_dfrbp_1 _34731_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net631),
    .D(_01421_),
    .Q_N(_15645_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[14] ));
 sg13g2_dfrbp_1 _34732_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net629),
    .D(_01422_),
    .Q_N(_15644_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[15] ));
 sg13g2_dfrbp_1 _34733_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net627),
    .D(_01423_),
    .Q_N(_15643_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[16] ));
 sg13g2_dfrbp_1 _34734_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net625),
    .D(_01424_),
    .Q_N(_15642_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[17] ));
 sg13g2_dfrbp_1 _34735_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net623),
    .D(_01425_),
    .Q_N(_15641_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[18] ));
 sg13g2_dfrbp_1 _34736_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net621),
    .D(_01426_),
    .Q_N(_15640_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[19] ));
 sg13g2_dfrbp_1 _34737_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net619),
    .D(_01427_),
    .Q_N(_15639_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[20] ));
 sg13g2_dfrbp_1 _34738_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net617),
    .D(_01428_),
    .Q_N(_15638_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[21] ));
 sg13g2_dfrbp_1 _34739_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net615),
    .D(_01429_),
    .Q_N(_15637_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[22] ));
 sg13g2_dfrbp_1 _34740_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net613),
    .D(_01430_),
    .Q_N(_15636_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[23] ));
 sg13g2_dfrbp_1 _34741_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net611),
    .D(_01431_),
    .Q_N(_15635_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[24] ));
 sg13g2_dfrbp_1 _34742_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net609),
    .D(_01432_),
    .Q_N(_15634_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[25] ));
 sg13g2_dfrbp_1 _34743_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net607),
    .D(_01433_),
    .Q_N(_15633_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[26] ));
 sg13g2_dfrbp_1 _34744_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net605),
    .D(_01434_),
    .Q_N(_15632_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[27] ));
 sg13g2_dfrbp_1 _34745_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net603),
    .D(_01435_),
    .Q_N(_15631_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[28] ));
 sg13g2_dfrbp_1 _34746_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net601),
    .D(_01436_),
    .Q_N(_15630_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[29] ));
 sg13g2_dfrbp_1 _34747_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net599),
    .D(_01437_),
    .Q_N(_15629_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[30] ));
 sg13g2_dfrbp_1 _34748_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net597),
    .D(_01438_),
    .Q_N(_15628_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ALUOut[31] ));
 sg13g2_dfrbp_1 _34749_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net595),
    .D(_01439_),
    .Q_N(_15627_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[0] ));
 sg13g2_dfrbp_1 _34750_ (.CLK(clknet_leaf_273_clk),
    .RESET_B(net593),
    .D(net4542),
    .Q_N(_15626_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[1] ));
 sg13g2_dfrbp_1 _34751_ (.CLK(clknet_leaf_273_clk),
    .RESET_B(net591),
    .D(net4591),
    .Q_N(_15625_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[2] ));
 sg13g2_dfrbp_1 _34752_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net589),
    .D(_01442_),
    .Q_N(_15624_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[3] ));
 sg13g2_dfrbp_1 _34753_ (.CLK(clknet_leaf_275_clk),
    .RESET_B(net587),
    .D(net4973),
    .Q_N(_15623_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[4] ));
 sg13g2_dfrbp_1 _34754_ (.CLK(clknet_leaf_275_clk),
    .RESET_B(net585),
    .D(net5242),
    .Q_N(_15622_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[5] ));
 sg13g2_dfrbp_1 _34755_ (.CLK(clknet_leaf_275_clk),
    .RESET_B(net583),
    .D(net5158),
    .Q_N(_15621_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[6] ));
 sg13g2_dfrbp_1 _34756_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net581),
    .D(net4527),
    .Q_N(_15620_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[7] ));
 sg13g2_dfrbp_1 _34757_ (.CLK(clknet_leaf_273_clk),
    .RESET_B(net579),
    .D(net5329),
    .Q_N(_15619_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[8] ));
 sg13g2_dfrbp_1 _34758_ (.CLK(clknet_leaf_273_clk),
    .RESET_B(net577),
    .D(net5451),
    .Q_N(_15618_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[9] ));
 sg13g2_dfrbp_1 _34759_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net575),
    .D(_01449_),
    .Q_N(_15617_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[10] ));
 sg13g2_dfrbp_1 _34760_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net573),
    .D(net4331),
    .Q_N(_15616_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[11] ));
 sg13g2_dfrbp_1 _34761_ (.CLK(clknet_leaf_273_clk),
    .RESET_B(net571),
    .D(net5440),
    .Q_N(_15615_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[12] ));
 sg13g2_dfrbp_1 _34762_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net569),
    .D(_01452_),
    .Q_N(_15614_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[13] ));
 sg13g2_dfrbp_1 _34763_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net567),
    .D(_01453_),
    .Q_N(_15613_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[14] ));
 sg13g2_dfrbp_1 _34764_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net565),
    .D(net4227),
    .Q_N(_15612_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[15] ));
 sg13g2_dfrbp_1 _34765_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net563),
    .D(net5227),
    .Q_N(_15611_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[16] ));
 sg13g2_dfrbp_1 _34766_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net561),
    .D(_01456_),
    .Q_N(_15610_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[17] ));
 sg13g2_dfrbp_1 _34767_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net559),
    .D(net5371),
    .Q_N(_15609_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[18] ));
 sg13g2_dfrbp_1 _34768_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net557),
    .D(net5309),
    .Q_N(_15608_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[19] ));
 sg13g2_dfrbp_1 _34769_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net555),
    .D(_01459_),
    .Q_N(_15607_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[20] ));
 sg13g2_dfrbp_1 _34770_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net553),
    .D(net4786),
    .Q_N(_15606_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[21] ));
 sg13g2_dfrbp_1 _34771_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net551),
    .D(net5128),
    .Q_N(_15605_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[22] ));
 sg13g2_dfrbp_1 _34772_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net549),
    .D(net4589),
    .Q_N(_15604_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[23] ));
 sg13g2_dfrbp_1 _34773_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net547),
    .D(_01463_),
    .Q_N(_15603_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[24] ));
 sg13g2_dfrbp_1 _34774_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net545),
    .D(net5312),
    .Q_N(_15602_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[25] ));
 sg13g2_dfrbp_1 _34775_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net543),
    .D(net5090),
    .Q_N(_15601_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[26] ));
 sg13g2_dfrbp_1 _34776_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net541),
    .D(net4784),
    .Q_N(_15600_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[27] ));
 sg13g2_dfrbp_1 _34777_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net539),
    .D(net5025),
    .Q_N(_15599_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[28] ));
 sg13g2_dfrbp_1 _34778_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net537),
    .D(net4354),
    .Q_N(_15598_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[29] ));
 sg13g2_dfrbp_1 _34779_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net535),
    .D(net4243),
    .Q_N(_15597_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[30] ));
 sg13g2_dfrbp_1 _34780_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net533),
    .D(net4982),
    .Q_N(_15596_),
    .Q(\soc_I.kianv_I.datapath_unit_I.OldPC[31] ));
 sg13g2_dfrbp_1 _34781_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net531),
    .D(_01471_),
    .Q_N(_15595_),
    .Q(\soc_I.kianv_I.amo_reserved_state_load ));
 sg13g2_dfrbp_1 _34782_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net529),
    .D(_01472_),
    .Q_N(_15594_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[0] ));
 sg13g2_dfrbp_1 _34783_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net527),
    .D(_01473_),
    .Q_N(_15593_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[1] ));
 sg13g2_dfrbp_1 _34784_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net525),
    .D(_01474_),
    .Q_N(_15592_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[2] ));
 sg13g2_dfrbp_1 _34785_ (.CLK(clknet_leaf_269_clk),
    .RESET_B(net523),
    .D(_01475_),
    .Q_N(_15591_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[3] ));
 sg13g2_dfrbp_1 _34786_ (.CLK(clknet_leaf_268_clk),
    .RESET_B(net521),
    .D(_01476_),
    .Q_N(_15590_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[4] ));
 sg13g2_dfrbp_1 _34787_ (.CLK(clknet_leaf_266_clk),
    .RESET_B(net519),
    .D(_01477_),
    .Q_N(_15589_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[5] ));
 sg13g2_dfrbp_1 _34788_ (.CLK(clknet_leaf_269_clk),
    .RESET_B(net517),
    .D(_01478_),
    .Q_N(_15588_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[6] ));
 sg13g2_dfrbp_1 _34789_ (.CLK(clknet_leaf_270_clk),
    .RESET_B(net515),
    .D(_01479_),
    .Q_N(_15587_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[7] ));
 sg13g2_dfrbp_1 _34790_ (.CLK(clknet_leaf_265_clk),
    .RESET_B(net513),
    .D(_01480_),
    .Q_N(_15586_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[8] ));
 sg13g2_dfrbp_1 _34791_ (.CLK(clknet_leaf_266_clk),
    .RESET_B(net511),
    .D(_01481_),
    .Q_N(_15585_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[9] ));
 sg13g2_dfrbp_1 _34792_ (.CLK(clknet_leaf_270_clk),
    .RESET_B(net509),
    .D(_01482_),
    .Q_N(_15584_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[10] ));
 sg13g2_dfrbp_1 _34793_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net507),
    .D(_01483_),
    .Q_N(_15583_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[11] ));
 sg13g2_dfrbp_1 _34794_ (.CLK(clknet_leaf_268_clk),
    .RESET_B(net505),
    .D(_01484_),
    .Q_N(_15582_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[12] ));
 sg13g2_dfrbp_1 _34795_ (.CLK(clknet_leaf_268_clk),
    .RESET_B(net503),
    .D(_01485_),
    .Q_N(_15581_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[13] ));
 sg13g2_dfrbp_1 _34796_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net501),
    .D(_01486_),
    .Q_N(_15580_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[14] ));
 sg13g2_dfrbp_1 _34797_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net499),
    .D(_01487_),
    .Q_N(_15579_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[15] ));
 sg13g2_dfrbp_1 _34798_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net497),
    .D(_01488_),
    .Q_N(_15578_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[16] ));
 sg13g2_dfrbp_1 _34799_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net495),
    .D(_01489_),
    .Q_N(_15577_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[17] ));
 sg13g2_dfrbp_1 _34800_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net493),
    .D(_01490_),
    .Q_N(_15576_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[18] ));
 sg13g2_dfrbp_1 _34801_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net491),
    .D(_01491_),
    .Q_N(_15575_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[19] ));
 sg13g2_dfrbp_1 _34802_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net489),
    .D(_01492_),
    .Q_N(_15574_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[20] ));
 sg13g2_dfrbp_1 _34803_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net487),
    .D(_01493_),
    .Q_N(_15573_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[21] ));
 sg13g2_dfrbp_1 _34804_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net485),
    .D(_01494_),
    .Q_N(_15572_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[22] ));
 sg13g2_dfrbp_1 _34805_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net483),
    .D(_01495_),
    .Q_N(_15571_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[23] ));
 sg13g2_dfrbp_1 _34806_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net481),
    .D(_01496_),
    .Q_N(_15570_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[24] ));
 sg13g2_dfrbp_1 _34807_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net479),
    .D(_01497_),
    .Q_N(_15569_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[25] ));
 sg13g2_dfrbp_1 _34808_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net477),
    .D(_01498_),
    .Q_N(_15568_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[26] ));
 sg13g2_dfrbp_1 _34809_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net475),
    .D(_01499_),
    .Q_N(_15567_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[27] ));
 sg13g2_dfrbp_1 _34810_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net473),
    .D(_01500_),
    .Q_N(_15566_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[28] ));
 sg13g2_dfrbp_1 _34811_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net471),
    .D(_01501_),
    .Q_N(_15565_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[29] ));
 sg13g2_dfrbp_1 _34812_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net469),
    .D(_01502_),
    .Q_N(_15564_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[30] ));
 sg13g2_dfrbp_1 _34813_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net467),
    .D(_01503_),
    .Q_N(_15563_),
    .Q(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[31] ));
 sg13g2_dfrbp_1 _34814_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net465),
    .D(_01504_),
    .Q_N(_15562_),
    .Q(\soc_I.kianv_I.Instr[0] ));
 sg13g2_dfrbp_1 _34815_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net463),
    .D(_01505_),
    .Q_N(_15561_),
    .Q(\soc_I.kianv_I.Instr[1] ));
 sg13g2_dfrbp_1 _34816_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net461),
    .D(_01506_),
    .Q_N(_15560_),
    .Q(\soc_I.kianv_I.Instr[2] ));
 sg13g2_dfrbp_1 _34817_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net459),
    .D(_01507_),
    .Q_N(_15559_),
    .Q(\soc_I.kianv_I.Instr[3] ));
 sg13g2_dfrbp_1 _34818_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net457),
    .D(_01508_),
    .Q_N(_15558_),
    .Q(\soc_I.kianv_I.Instr[4] ));
 sg13g2_dfrbp_1 _34819_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net455),
    .D(_01509_),
    .Q_N(_15557_),
    .Q(\soc_I.kianv_I.Instr[5] ));
 sg13g2_dfrbp_1 _34820_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net453),
    .D(_01510_),
    .Q_N(_00214_),
    .Q(\soc_I.kianv_I.Instr[6] ));
 sg13g2_dfrbp_1 _34821_ (.CLK(clknet_leaf_277_clk),
    .RESET_B(net451),
    .D(_01511_),
    .Q_N(_15556_),
    .Q(\soc_I.kianv_I.Instr[7] ));
 sg13g2_dfrbp_1 _34822_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net449),
    .D(_01512_),
    .Q_N(_15555_),
    .Q(\soc_I.kianv_I.Instr[8] ));
 sg13g2_dfrbp_1 _34823_ (.CLK(clknet_leaf_265_clk),
    .RESET_B(net447),
    .D(_01513_),
    .Q_N(_00185_),
    .Q(\soc_I.kianv_I.Instr[9] ));
 sg13g2_dfrbp_1 _34824_ (.CLK(clknet_leaf_272_clk),
    .RESET_B(net445),
    .D(_01514_),
    .Q_N(_15554_),
    .Q(\soc_I.kianv_I.Instr[10] ));
 sg13g2_dfrbp_1 _34825_ (.CLK(clknet_leaf_271_clk),
    .RESET_B(net443),
    .D(_01515_),
    .Q_N(_15553_),
    .Q(\soc_I.kianv_I.Instr[11] ));
 sg13g2_dfrbp_1 _34826_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net441),
    .D(_01516_),
    .Q_N(_00212_),
    .Q(\soc_I.kianv_I.Instr[12] ));
 sg13g2_dfrbp_1 _34827_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net439),
    .D(_01517_),
    .Q_N(_15552_),
    .Q(\soc_I.kianv_I.Instr[13] ));
 sg13g2_dfrbp_1 _34828_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net437),
    .D(_01518_),
    .Q_N(_00188_),
    .Q(\soc_I.kianv_I.Instr[14] ));
 sg13g2_dfrbp_1 _34829_ (.CLK(clknet_leaf_284_clk),
    .RESET_B(net435),
    .D(_01519_),
    .Q_N(_15551_),
    .Q(\soc_I.kianv_I.Instr[15] ));
 sg13g2_dfrbp_1 _34830_ (.CLK(clknet_leaf_280_clk),
    .RESET_B(net433),
    .D(_01520_),
    .Q_N(_00293_),
    .Q(\soc_I.kianv_I.Instr[16] ));
 sg13g2_dfrbp_1 _34831_ (.CLK(clknet_leaf_266_clk),
    .RESET_B(net431),
    .D(_01521_),
    .Q_N(_00294_),
    .Q(\soc_I.kianv_I.Instr[17] ));
 sg13g2_dfrbp_1 _34832_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net429),
    .D(_01522_),
    .Q_N(_00295_),
    .Q(\soc_I.kianv_I.Instr[18] ));
 sg13g2_dfrbp_1 _34833_ (.CLK(clknet_leaf_277_clk),
    .RESET_B(net427),
    .D(_01523_),
    .Q_N(_00296_),
    .Q(\soc_I.kianv_I.Instr[19] ));
 sg13g2_dfrbp_1 _34834_ (.CLK(clknet_leaf_290_clk),
    .RESET_B(net425),
    .D(_01524_),
    .Q_N(_15550_),
    .Q(\soc_I.kianv_I.Instr[20] ));
 sg13g2_dfrbp_1 _34835_ (.CLK(clknet_leaf_277_clk),
    .RESET_B(net423),
    .D(_01525_),
    .Q_N(_00216_),
    .Q(\soc_I.kianv_I.Instr[21] ));
 sg13g2_dfrbp_1 _34836_ (.CLK(clknet_leaf_275_clk),
    .RESET_B(net421),
    .D(_01526_),
    .Q_N(_00215_),
    .Q(\soc_I.kianv_I.Instr[22] ));
 sg13g2_dfrbp_1 _34837_ (.CLK(clknet_leaf_276_clk),
    .RESET_B(net419),
    .D(_01527_),
    .Q_N(_00238_),
    .Q(\soc_I.kianv_I.Instr[23] ));
 sg13g2_dfrbp_1 _34838_ (.CLK(clknet_leaf_272_clk),
    .RESET_B(net417),
    .D(_01528_),
    .Q_N(_00236_),
    .Q(\soc_I.kianv_I.Instr[24] ));
 sg13g2_dfrbp_1 _34839_ (.CLK(clknet_leaf_271_clk),
    .RESET_B(net415),
    .D(_01529_),
    .Q_N(_00285_),
    .Q(\soc_I.kianv_I.Instr[25] ));
 sg13g2_dfrbp_1 _34840_ (.CLK(clknet_leaf_271_clk),
    .RESET_B(net413),
    .D(_01530_),
    .Q_N(_15549_),
    .Q(\soc_I.kianv_I.Instr[26] ));
 sg13g2_dfrbp_1 _34841_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net411),
    .D(_01531_),
    .Q_N(_15548_),
    .Q(\soc_I.kianv_I.Instr[27] ));
 sg13g2_dfrbp_1 _34842_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net409),
    .D(_01532_),
    .Q_N(_15547_),
    .Q(\soc_I.kianv_I.Instr[28] ));
 sg13g2_dfrbp_1 _34843_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net407),
    .D(_01533_),
    .Q_N(_15546_),
    .Q(\soc_I.kianv_I.Instr[29] ));
 sg13g2_dfrbp_1 _34844_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net405),
    .D(_01534_),
    .Q_N(_00213_),
    .Q(\soc_I.kianv_I.Instr[30] ));
 sg13g2_dfrbp_1 _34845_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net403),
    .D(_01535_),
    .Q_N(_00189_),
    .Q(\soc_I.kianv_I.Instr[31] ));
 sg13g2_dfrbp_1 _34846_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net401),
    .D(_01536_),
    .Q_N(_15545_),
    .Q(\soc_I.PC[0] ));
 sg13g2_dfrbp_1 _34847_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net399),
    .D(_01537_),
    .Q_N(_15544_),
    .Q(\soc_I.PC[1] ));
 sg13g2_dfrbp_1 _34848_ (.CLK(clknet_leaf_272_clk),
    .RESET_B(net397),
    .D(_01538_),
    .Q_N(_15543_),
    .Q(\soc_I.PC[2] ));
 sg13g2_dfrbp_1 _34849_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net395),
    .D(_01539_),
    .Q_N(_15542_),
    .Q(\soc_I.PC[3] ));
 sg13g2_dfrbp_1 _34850_ (.CLK(clknet_leaf_277_clk),
    .RESET_B(net393),
    .D(_01540_),
    .Q_N(_15541_),
    .Q(\soc_I.PC[4] ));
 sg13g2_dfrbp_1 _34851_ (.CLK(clknet_leaf_276_clk),
    .RESET_B(net391),
    .D(net5324),
    .Q_N(_15540_),
    .Q(\soc_I.PC[5] ));
 sg13g2_dfrbp_1 _34852_ (.CLK(clknet_leaf_276_clk),
    .RESET_B(net389),
    .D(_01542_),
    .Q_N(_15539_),
    .Q(\soc_I.PC[6] ));
 sg13g2_dfrbp_1 _34853_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net387),
    .D(_01543_),
    .Q_N(_15538_),
    .Q(\soc_I.PC[7] ));
 sg13g2_dfrbp_1 _34854_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net385),
    .D(_01544_),
    .Q_N(_15537_),
    .Q(\soc_I.PC[8] ));
 sg13g2_dfrbp_1 _34855_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net383),
    .D(net5331),
    .Q_N(_15536_),
    .Q(\soc_I.PC[9] ));
 sg13g2_dfrbp_1 _34856_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net381),
    .D(_01546_),
    .Q_N(_15535_),
    .Q(\soc_I.PC[10] ));
 sg13g2_dfrbp_1 _34857_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net379),
    .D(_01547_),
    .Q_N(_15534_),
    .Q(\soc_I.PC[11] ));
 sg13g2_dfrbp_1 _34858_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net377),
    .D(_01548_),
    .Q_N(_15533_),
    .Q(\soc_I.PC[12] ));
 sg13g2_dfrbp_1 _34859_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net375),
    .D(_01549_),
    .Q_N(_15532_),
    .Q(\soc_I.PC[13] ));
 sg13g2_dfrbp_1 _34860_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net373),
    .D(_01550_),
    .Q_N(_15531_),
    .Q(\soc_I.PC[14] ));
 sg13g2_dfrbp_1 _34861_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net371),
    .D(_01551_),
    .Q_N(_15530_),
    .Q(\soc_I.PC[15] ));
 sg13g2_dfrbp_1 _34862_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net369),
    .D(_01552_),
    .Q_N(_15529_),
    .Q(\led[0] ));
 sg13g2_dfrbp_1 _34863_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net367),
    .D(_01553_),
    .Q_N(_15528_),
    .Q(\led[1] ));
 sg13g2_dfrbp_1 _34864_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net365),
    .D(_01554_),
    .Q_N(_15527_),
    .Q(\led[2] ));
 sg13g2_dfrbp_1 _34865_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net363),
    .D(_01555_),
    .Q_N(_15526_),
    .Q(\led[3] ));
 sg13g2_dfrbp_1 _34866_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net361),
    .D(_01556_),
    .Q_N(_15525_),
    .Q(\soc_I.PC[20] ));
 sg13g2_dfrbp_1 _34867_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net359),
    .D(_01557_),
    .Q_N(_15524_),
    .Q(\soc_I.PC[21] ));
 sg13g2_dfrbp_1 _34868_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net357),
    .D(_01558_),
    .Q_N(_15523_),
    .Q(\soc_I.PC[22] ));
 sg13g2_dfrbp_1 _34869_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net355),
    .D(net5259),
    .Q_N(_15522_),
    .Q(\soc_I.PC[23] ));
 sg13g2_dfrbp_1 _34870_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net353),
    .D(_01560_),
    .Q_N(_15521_),
    .Q(\soc_I.PC[24] ));
 sg13g2_dfrbp_1 _34871_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net351),
    .D(_01561_),
    .Q_N(_15520_),
    .Q(\soc_I.PC[25] ));
 sg13g2_dfrbp_1 _34872_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net349),
    .D(_01562_),
    .Q_N(_15519_),
    .Q(\soc_I.PC[26] ));
 sg13g2_dfrbp_1 _34873_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net347),
    .D(_01563_),
    .Q_N(_15518_),
    .Q(\soc_I.PC[27] ));
 sg13g2_dfrbp_1 _34874_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net345),
    .D(_01564_),
    .Q_N(_15517_),
    .Q(\soc_I.PC[28] ));
 sg13g2_dfrbp_1 _34875_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net343),
    .D(_01565_),
    .Q_N(_15516_),
    .Q(\soc_I.PC[29] ));
 sg13g2_dfrbp_1 _34876_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net341),
    .D(_01566_),
    .Q_N(_15515_),
    .Q(\soc_I.PC[30] ));
 sg13g2_dfrbp_1 _34877_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net339),
    .D(_01567_),
    .Q_N(_15514_),
    .Q(\soc_I.PC[31] ));
 sg13g2_dfrbp_1 _34878_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net337),
    .D(_01568_),
    .Q_N(_15513_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][0] ));
 sg13g2_dfrbp_1 _34879_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net336),
    .D(_01569_),
    .Q_N(_15512_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][1] ));
 sg13g2_dfrbp_1 _34880_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net335),
    .D(_01570_),
    .Q_N(_15511_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][2] ));
 sg13g2_dfrbp_1 _34881_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net334),
    .D(_01571_),
    .Q_N(_15510_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][3] ));
 sg13g2_dfrbp_1 _34882_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net333),
    .D(_01572_),
    .Q_N(_15509_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][4] ));
 sg13g2_dfrbp_1 _34883_ (.CLK(clknet_leaf_265_clk),
    .RESET_B(net332),
    .D(_01573_),
    .Q_N(_15508_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][5] ));
 sg13g2_dfrbp_1 _34884_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net331),
    .D(_01574_),
    .Q_N(_15507_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][6] ));
 sg13g2_dfrbp_1 _34885_ (.CLK(clknet_leaf_305_clk),
    .RESET_B(net330),
    .D(_01575_),
    .Q_N(_15506_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][7] ));
 sg13g2_dfrbp_1 _34886_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net329),
    .D(_01576_),
    .Q_N(_15505_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][8] ));
 sg13g2_dfrbp_1 _34887_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net328),
    .D(_01577_),
    .Q_N(_15504_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][9] ));
 sg13g2_dfrbp_1 _34888_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net327),
    .D(_01578_),
    .Q_N(_15503_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][10] ));
 sg13g2_dfrbp_1 _34889_ (.CLK(clknet_leaf_316_clk),
    .RESET_B(net326),
    .D(_01579_),
    .Q_N(_15502_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][11] ));
 sg13g2_dfrbp_1 _34890_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net325),
    .D(_01580_),
    .Q_N(_15501_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][12] ));
 sg13g2_dfrbp_1 _34891_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net324),
    .D(_01581_),
    .Q_N(_15500_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][13] ));
 sg13g2_dfrbp_1 _34892_ (.CLK(clknet_leaf_289_clk),
    .RESET_B(net323),
    .D(_01582_),
    .Q_N(_15499_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][14] ));
 sg13g2_dfrbp_1 _34893_ (.CLK(clknet_leaf_309_clk),
    .RESET_B(net322),
    .D(_01583_),
    .Q_N(_15498_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][15] ));
 sg13g2_dfrbp_1 _34894_ (.CLK(clknet_leaf_317_clk),
    .RESET_B(net321),
    .D(_01584_),
    .Q_N(_15497_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][16] ));
 sg13g2_dfrbp_1 _34895_ (.CLK(clknet_leaf_312_clk),
    .RESET_B(net320),
    .D(_01585_),
    .Q_N(_15496_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][17] ));
 sg13g2_dfrbp_1 _34896_ (.CLK(clknet_leaf_308_clk),
    .RESET_B(net319),
    .D(_01586_),
    .Q_N(_15495_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][18] ));
 sg13g2_dfrbp_1 _34897_ (.CLK(clknet_leaf_288_clk),
    .RESET_B(net318),
    .D(_01587_),
    .Q_N(_15494_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][19] ));
 sg13g2_dfrbp_1 _34898_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net317),
    .D(_01588_),
    .Q_N(_15493_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][20] ));
 sg13g2_dfrbp_1 _34899_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net316),
    .D(_01589_),
    .Q_N(_15492_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][21] ));
 sg13g2_dfrbp_1 _34900_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net315),
    .D(_01590_),
    .Q_N(_15491_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][22] ));
 sg13g2_dfrbp_1 _34901_ (.CLK(clknet_leaf_305_clk),
    .RESET_B(net314),
    .D(_01591_),
    .Q_N(_15490_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][23] ));
 sg13g2_dfrbp_1 _34902_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net313),
    .D(_01592_),
    .Q_N(_15489_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][24] ));
 sg13g2_dfrbp_1 _34903_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net312),
    .D(_01593_),
    .Q_N(_15488_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][25] ));
 sg13g2_dfrbp_1 _34904_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net311),
    .D(_01594_),
    .Q_N(_15487_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][26] ));
 sg13g2_dfrbp_1 _34905_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net310),
    .D(_01595_),
    .Q_N(_15486_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][27] ));
 sg13g2_dfrbp_1 _34906_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net309),
    .D(_01596_),
    .Q_N(_15485_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][28] ));
 sg13g2_dfrbp_1 _34907_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net308),
    .D(_01597_),
    .Q_N(_15484_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][29] ));
 sg13g2_dfrbp_1 _34908_ (.CLK(clknet_leaf_291_clk),
    .RESET_B(net307),
    .D(_01598_),
    .Q_N(_15483_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][30] ));
 sg13g2_dfrbp_1 _34909_ (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1309),
    .D(_01599_),
    .Q_N(_16655_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][31] ));
 sg13g2_dfrbp_1 _34910_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1310),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[0] ),
    .Q_N(_16656_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[0] ));
 sg13g2_dfrbp_1 _34911_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1311),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[1] ),
    .Q_N(_16657_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[1] ));
 sg13g2_dfrbp_1 _34912_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1312),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[2] ),
    .Q_N(_16658_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[2] ));
 sg13g2_dfrbp_1 _34913_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1313),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[3] ),
    .Q_N(_16659_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[3] ));
 sg13g2_dfrbp_1 _34914_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1314),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[4] ),
    .Q_N(_16660_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[4] ));
 sg13g2_dfrbp_1 _34915_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1315),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[5] ),
    .Q_N(_16661_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[5] ));
 sg13g2_dfrbp_1 _34916_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1316),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[6] ),
    .Q_N(_16662_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[6] ));
 sg13g2_dfrbp_1 _34917_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1317),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[7] ),
    .Q_N(_16663_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[7] ));
 sg13g2_dfrbp_1 _34918_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1318),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[8] ),
    .Q_N(_16664_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[8] ));
 sg13g2_dfrbp_1 _34919_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1319),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[9] ),
    .Q_N(_16665_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[9] ));
 sg13g2_dfrbp_1 _34920_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1320),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[10] ),
    .Q_N(_16666_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[10] ));
 sg13g2_dfrbp_1 _34921_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1321),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[11] ),
    .Q_N(_16667_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[11] ));
 sg13g2_dfrbp_1 _34922_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1322),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[12] ),
    .Q_N(_16668_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[12] ));
 sg13g2_dfrbp_1 _34923_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1323),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[13] ),
    .Q_N(_16669_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[13] ));
 sg13g2_dfrbp_1 _34924_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1324),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[14] ),
    .Q_N(_16670_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[14] ));
 sg13g2_dfrbp_1 _34925_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1325),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[15] ),
    .Q_N(_16671_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[15] ));
 sg13g2_dfrbp_1 _34926_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1326),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[16] ),
    .Q_N(_16672_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[16] ));
 sg13g2_dfrbp_1 _34927_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1327),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[17] ),
    .Q_N(_16673_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[17] ));
 sg13g2_dfrbp_1 _34928_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1328),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[18] ),
    .Q_N(_16674_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[18] ));
 sg13g2_dfrbp_1 _34929_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1329),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[19] ),
    .Q_N(_16675_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[19] ));
 sg13g2_dfrbp_1 _34930_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1330),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[20] ),
    .Q_N(_16676_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[20] ));
 sg13g2_dfrbp_1 _34931_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1331),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[21] ),
    .Q_N(_16677_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[21] ));
 sg13g2_dfrbp_1 _34932_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1332),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[22] ),
    .Q_N(_16678_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[22] ));
 sg13g2_dfrbp_1 _34933_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1333),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[23] ),
    .Q_N(_16679_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[23] ));
 sg13g2_dfrbp_1 _34934_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1334),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[24] ),
    .Q_N(_16680_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[24] ));
 sg13g2_dfrbp_1 _34935_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1335),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[25] ),
    .Q_N(_16681_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[25] ));
 sg13g2_dfrbp_1 _34936_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1336),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[26] ),
    .Q_N(_16682_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[26] ));
 sg13g2_dfrbp_1 _34937_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1337),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[27] ),
    .Q_N(_16683_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[27] ));
 sg13g2_dfrbp_1 _34938_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1338),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[28] ),
    .Q_N(_16684_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[28] ));
 sg13g2_dfrbp_1 _34939_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1339),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[29] ),
    .Q_N(_16685_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[29] ));
 sg13g2_dfrbp_1 _34940_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1340),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[30] ),
    .Q_N(_16686_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[30] ));
 sg13g2_dfrbp_1 _34941_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1341),
    .D(\soc_I.kianv_I.datapath_unit_I.MULExtResult[31] ),
    .Q_N(_16687_),
    .Q(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[31] ));
 sg13g2_dfrbp_1 _34942_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1342),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[0] ),
    .Q_N(_16688_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[0] ));
 sg13g2_dfrbp_1 _34943_ (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1343),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[1] ),
    .Q_N(_16689_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[1] ));
 sg13g2_dfrbp_1 _34944_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1344),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[2] ),
    .Q_N(_16690_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[2] ));
 sg13g2_dfrbp_1 _34945_ (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1345),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[3] ),
    .Q_N(_16691_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[3] ));
 sg13g2_dfrbp_1 _34946_ (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1346),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[4] ),
    .Q_N(_16692_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[4] ));
 sg13g2_dfrbp_1 _34947_ (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1347),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[5] ),
    .Q_N(_16693_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[5] ));
 sg13g2_dfrbp_1 _34948_ (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1348),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[6] ),
    .Q_N(_16694_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[6] ));
 sg13g2_dfrbp_1 _34949_ (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1349),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[7] ),
    .Q_N(_16695_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[7] ));
 sg13g2_dfrbp_1 _34950_ (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1350),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[8] ),
    .Q_N(_16696_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[8] ));
 sg13g2_dfrbp_1 _34951_ (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1351),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[9] ),
    .Q_N(_16697_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[9] ));
 sg13g2_dfrbp_1 _34952_ (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1352),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[10] ),
    .Q_N(_16698_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[10] ));
 sg13g2_dfrbp_1 _34953_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1353),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[11] ),
    .Q_N(_16699_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[11] ));
 sg13g2_dfrbp_1 _34954_ (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1354),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[12] ),
    .Q_N(_16700_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[12] ));
 sg13g2_dfrbp_1 _34955_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1355),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[13] ),
    .Q_N(_16701_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[13] ));
 sg13g2_dfrbp_1 _34956_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1356),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[14] ),
    .Q_N(_16702_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[14] ));
 sg13g2_dfrbp_1 _34957_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1357),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[15] ),
    .Q_N(_16703_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[15] ));
 sg13g2_dfrbp_1 _34958_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1358),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[16] ),
    .Q_N(_16704_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[16] ));
 sg13g2_dfrbp_1 _34959_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1359),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[17] ),
    .Q_N(_16705_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[17] ));
 sg13g2_dfrbp_1 _34960_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1360),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[18] ),
    .Q_N(_16706_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[18] ));
 sg13g2_dfrbp_1 _34961_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1361),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[19] ),
    .Q_N(_16707_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[19] ));
 sg13g2_dfrbp_1 _34962_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1362),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[20] ),
    .Q_N(_16708_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[20] ));
 sg13g2_dfrbp_1 _34963_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1363),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[21] ),
    .Q_N(_16709_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[21] ));
 sg13g2_dfrbp_1 _34964_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1364),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[22] ),
    .Q_N(_16710_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[22] ));
 sg13g2_dfrbp_1 _34965_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1365),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[23] ),
    .Q_N(_16711_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[23] ));
 sg13g2_dfrbp_1 _34966_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1366),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[24] ),
    .Q_N(_16712_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[24] ));
 sg13g2_dfrbp_1 _34967_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1367),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[25] ),
    .Q_N(_16713_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[25] ));
 sg13g2_dfrbp_1 _34968_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1368),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[26] ),
    .Q_N(_16714_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[26] ));
 sg13g2_dfrbp_1 _34969_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1369),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[27] ),
    .Q_N(_16715_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[27] ));
 sg13g2_dfrbp_1 _34970_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1370),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[28] ),
    .Q_N(_16716_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[28] ));
 sg13g2_dfrbp_1 _34971_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1371),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[29] ),
    .Q_N(_16717_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[29] ));
 sg13g2_dfrbp_1 _34972_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1372),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[30] ),
    .Q_N(_16718_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[30] ));
 sg13g2_dfrbp_1 _34973_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1373),
    .D(\soc_I.kianv_I.datapath_unit_I.CSRData[31] ),
    .Q_N(_16719_),
    .Q(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[31] ));
 sg13g2_dfrbp_1 _34974_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1374),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[0] ),
    .Q_N(_16720_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[0] ));
 sg13g2_dfrbp_1 _34975_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1375),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[1] ),
    .Q_N(_16721_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[1] ));
 sg13g2_dfrbp_1 _34976_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1376),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[2] ),
    .Q_N(_16722_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[2] ));
 sg13g2_dfrbp_1 _34977_ (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1377),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[3] ),
    .Q_N(_16723_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[3] ));
 sg13g2_dfrbp_1 _34978_ (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1378),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[4] ),
    .Q_N(_16724_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[4] ));
 sg13g2_dfrbp_1 _34979_ (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1379),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[5] ),
    .Q_N(_16725_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[5] ));
 sg13g2_dfrbp_1 _34980_ (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1380),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[6] ),
    .Q_N(_16726_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[6] ));
 sg13g2_dfrbp_1 _34981_ (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1381),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[7] ),
    .Q_N(_16727_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[7] ));
 sg13g2_dfrbp_1 _34982_ (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1382),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[8] ),
    .Q_N(_16728_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[8] ));
 sg13g2_dfrbp_1 _34983_ (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1383),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[9] ),
    .Q_N(_16729_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[9] ));
 sg13g2_dfrbp_1 _34984_ (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1384),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[10] ),
    .Q_N(_16730_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[10] ));
 sg13g2_dfrbp_1 _34985_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1385),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[11] ),
    .Q_N(_16731_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[11] ));
 sg13g2_dfrbp_1 _34986_ (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1386),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[12] ),
    .Q_N(_16732_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[12] ));
 sg13g2_dfrbp_1 _34987_ (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1387),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[13] ),
    .Q_N(_16733_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[13] ));
 sg13g2_dfrbp_1 _34988_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1388),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[14] ),
    .Q_N(_16734_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[14] ));
 sg13g2_dfrbp_1 _34989_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1389),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[15] ),
    .Q_N(_16735_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[15] ));
 sg13g2_dfrbp_1 _34990_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1390),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[16] ),
    .Q_N(_16736_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[16] ));
 sg13g2_dfrbp_1 _34991_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1391),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[17] ),
    .Q_N(_16737_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[17] ));
 sg13g2_dfrbp_1 _34992_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1392),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[18] ),
    .Q_N(_16738_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[18] ));
 sg13g2_dfrbp_1 _34993_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1393),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[19] ),
    .Q_N(_16739_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[19] ));
 sg13g2_dfrbp_1 _34994_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1394),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[20] ),
    .Q_N(_16740_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[20] ));
 sg13g2_dfrbp_1 _34995_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1395),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[21] ),
    .Q_N(_16741_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[21] ));
 sg13g2_dfrbp_1 _34996_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1396),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[22] ),
    .Q_N(_16742_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[22] ));
 sg13g2_dfrbp_1 _34997_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1397),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[23] ),
    .Q_N(_16743_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[23] ));
 sg13g2_dfrbp_1 _34998_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1398),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[24] ),
    .Q_N(_16744_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[24] ));
 sg13g2_dfrbp_1 _34999_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1399),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[25] ),
    .Q_N(_16745_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[25] ));
 sg13g2_dfrbp_1 _35000_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1400),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[26] ),
    .Q_N(_16746_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[26] ));
 sg13g2_dfrbp_1 _35001_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1401),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[27] ),
    .Q_N(_16747_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[27] ));
 sg13g2_dfrbp_1 _35002_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1402),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[28] ),
    .Q_N(_16748_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[28] ));
 sg13g2_dfrbp_1 _35003_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1403),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[29] ),
    .Q_N(_16749_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[29] ));
 sg13g2_dfrbp_1 _35004_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1405),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[30] ),
    .Q_N(_16750_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[30] ));
 sg13g2_dfrbp_1 _35005_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net306),
    .D(\soc_I.kianv_I.datapath_unit_I.Data[31] ),
    .Q_N(_15482_),
    .Q(\soc_I.kianv_I.datapath_unit_I.DataLatched[31] ));
 sg13g2_dfrbp_1 _35006_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1406),
    .D(_01600_),
    .Q_N(_16751_),
    .Q(\soc_I.gpio0_I.ready ));
 sg13g2_dfrbp_1 _35007_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net2333),
    .D(\soc_I.clint_I.addr[0] ),
    .Q_N(_16752_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ADDR_I.q[0] ));
 sg13g2_dfrbp_1 _35008_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net305),
    .D(\soc_I.clint_I.addr[1] ),
    .Q_N(_15481_),
    .Q(\soc_I.kianv_I.datapath_unit_I.ADDR_I.q[1] ));
 sg13g2_dfrbp_1 _35009_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net304),
    .D(_01601_),
    .Q_N(_00303_),
    .Q(\soc_I.clint_I.tick_cnt[0] ));
 sg13g2_dfrbp_1 _35010_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net303),
    .D(_01602_),
    .Q_N(_15480_),
    .Q(\soc_I.clint_I.tick_cnt[1] ));
 sg13g2_dfrbp_1 _35011_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net302),
    .D(net3627),
    .Q_N(_15479_),
    .Q(\soc_I.clint_I.tick_cnt[2] ));
 sg13g2_dfrbp_1 _35012_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net301),
    .D(_01604_),
    .Q_N(_15478_),
    .Q(\soc_I.clint_I.tick_cnt[3] ));
 sg13g2_dfrbp_1 _35013_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net300),
    .D(_01605_),
    .Q_N(_15477_),
    .Q(\soc_I.clint_I.tick_cnt[4] ));
 sg13g2_dfrbp_1 _35014_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net299),
    .D(_01606_),
    .Q_N(_15476_),
    .Q(\soc_I.clint_I.tick_cnt[5] ));
 sg13g2_dfrbp_1 _35015_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net298),
    .D(_01607_),
    .Q_N(_15475_),
    .Q(\soc_I.clint_I.tick_cnt[6] ));
 sg13g2_dfrbp_1 _35016_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net297),
    .D(_01608_),
    .Q_N(_15474_),
    .Q(\soc_I.clint_I.tick_cnt[7] ));
 sg13g2_dfrbp_1 _35017_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net296),
    .D(_01609_),
    .Q_N(_15473_),
    .Q(\soc_I.clint_I.tick_cnt[8] ));
 sg13g2_dfrbp_1 _35018_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net295),
    .D(_01610_),
    .Q_N(_15472_),
    .Q(\soc_I.clint_I.tick_cnt[9] ));
 sg13g2_dfrbp_1 _35019_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net294),
    .D(_01611_),
    .Q_N(_15471_),
    .Q(\soc_I.clint_I.tick_cnt[10] ));
 sg13g2_dfrbp_1 _35020_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net293),
    .D(_01612_),
    .Q_N(_15470_),
    .Q(\soc_I.clint_I.tick_cnt[11] ));
 sg13g2_dfrbp_1 _35021_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net292),
    .D(_01613_),
    .Q_N(_15469_),
    .Q(\soc_I.clint_I.tick_cnt[12] ));
 sg13g2_dfrbp_1 _35022_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net291),
    .D(_01614_),
    .Q_N(_15468_),
    .Q(\soc_I.clint_I.tick_cnt[13] ));
 sg13g2_dfrbp_1 _35023_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net290),
    .D(_01615_),
    .Q_N(_15467_),
    .Q(\soc_I.clint_I.tick_cnt[14] ));
 sg13g2_dfrbp_1 _35024_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net289),
    .D(_01616_),
    .Q_N(_15466_),
    .Q(\soc_I.clint_I.tick_cnt[15] ));
 sg13g2_dfrbp_1 _35025_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net288),
    .D(_01617_),
    .Q_N(_15465_),
    .Q(\soc_I.clint_I.tick_cnt[16] ));
 sg13g2_dfrbp_1 _35026_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net287),
    .D(_01618_),
    .Q_N(_15464_),
    .Q(\soc_I.clint_I.tick_cnt[17] ));
 sg13g2_dfrbp_1 _35027_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net286),
    .D(_01619_),
    .Q_N(_15463_),
    .Q(\soc_I.IRQ3 ));
 sg13g2_dfrbp_1 _35028_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net284),
    .D(_01620_),
    .Q_N(_00111_),
    .Q(\soc_I.clint_I.mtimecmp[32] ));
 sg13g2_dfrbp_1 _35029_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net282),
    .D(_01621_),
    .Q_N(_00116_),
    .Q(\soc_I.clint_I.mtimecmp[33] ));
 sg13g2_dfrbp_1 _35030_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net280),
    .D(_01622_),
    .Q_N(_00121_),
    .Q(\soc_I.clint_I.mtimecmp[34] ));
 sg13g2_dfrbp_1 _35031_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net278),
    .D(_01623_),
    .Q_N(_00126_),
    .Q(\soc_I.clint_I.mtimecmp[35] ));
 sg13g2_dfrbp_1 _35032_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net276),
    .D(_01624_),
    .Q_N(_00131_),
    .Q(\soc_I.clint_I.mtimecmp[36] ));
 sg13g2_dfrbp_1 _35033_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net274),
    .D(_01625_),
    .Q_N(_00136_),
    .Q(\soc_I.clint_I.mtimecmp[37] ));
 sg13g2_dfrbp_1 _35034_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net272),
    .D(_01626_),
    .Q_N(_00141_),
    .Q(\soc_I.clint_I.mtimecmp[38] ));
 sg13g2_dfrbp_1 _35035_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net270),
    .D(_01627_),
    .Q_N(_00146_),
    .Q(\soc_I.clint_I.mtimecmp[39] ));
 sg13g2_dfrbp_1 _35036_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net268),
    .D(_01628_),
    .Q_N(_15462_),
    .Q(\soc_I.rst_cnt[0] ));
 sg13g2_dfrbp_1 _35037_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net267),
    .D(_01629_),
    .Q_N(_15461_),
    .Q(\soc_I.rst_cnt[1] ));
 sg13g2_dfrbp_1 _35038_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net266),
    .D(_01630_),
    .Q_N(_15460_),
    .Q(\soc_I.rst_cnt[2] ));
 sg13g2_dfrbp_1 _35039_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net265),
    .D(_01631_),
    .Q_N(_00245_),
    .Q(\soc_I.clint_I.resetn ));
 sg13g2_dfrbp_1 _35040_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net264),
    .D(net3911),
    .Q_N(_00302_),
    .Q(\soc_I.clint_I.mtime[0] ));
 sg13g2_dfrbp_1 _35041_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net262),
    .D(_01633_),
    .Q_N(_00117_),
    .Q(\soc_I.clint_I.mtime[1] ));
 sg13g2_dfrbp_1 _35042_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net260),
    .D(net5516),
    .Q_N(_00122_),
    .Q(\soc_I.clint_I.mtime[2] ));
 sg13g2_dfrbp_1 _35043_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net258),
    .D(net3695),
    .Q_N(_00127_),
    .Q(\soc_I.clint_I.mtime[3] ));
 sg13g2_dfrbp_1 _35044_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net256),
    .D(net4490),
    .Q_N(_00132_),
    .Q(\soc_I.clint_I.mtime[4] ));
 sg13g2_dfrbp_1 _35045_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net254),
    .D(net3594),
    .Q_N(_00137_),
    .Q(\soc_I.clint_I.mtime[5] ));
 sg13g2_dfrbp_1 _35046_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net252),
    .D(_01638_),
    .Q_N(_00142_),
    .Q(\soc_I.clint_I.mtime[6] ));
 sg13g2_dfrbp_1 _35047_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net250),
    .D(net3414),
    .Q_N(_00147_),
    .Q(\soc_I.clint_I.mtime[7] ));
 sg13g2_dfrbp_1 _35048_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net248),
    .D(_01640_),
    .Q_N(_00077_),
    .Q(\soc_I.clint_I.mtime[8] ));
 sg13g2_dfrbp_1 _35049_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net246),
    .D(net4333),
    .Q_N(_00081_),
    .Q(\soc_I.clint_I.mtime[9] ));
 sg13g2_dfrbp_1 _35050_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net244),
    .D(_01642_),
    .Q_N(_00085_),
    .Q(\soc_I.clint_I.mtime[10] ));
 sg13g2_dfrbp_1 _35051_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net242),
    .D(net4519),
    .Q_N(_00089_),
    .Q(\soc_I.clint_I.mtime[11] ));
 sg13g2_dfrbp_1 _35052_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net240),
    .D(net5189),
    .Q_N(_00093_),
    .Q(\soc_I.clint_I.mtime[12] ));
 sg13g2_dfrbp_1 _35053_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net238),
    .D(net4503),
    .Q_N(_00097_),
    .Q(\soc_I.clint_I.mtime[13] ));
 sg13g2_dfrbp_1 _35054_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net236),
    .D(net5244),
    .Q_N(_00101_),
    .Q(\soc_I.clint_I.mtime[14] ));
 sg13g2_dfrbp_1 _35055_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net234),
    .D(net4603),
    .Q_N(_00105_),
    .Q(\soc_I.clint_I.mtime[15] ));
 sg13g2_dfrbp_1 _35056_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net232),
    .D(net5429),
    .Q_N(_00015_),
    .Q(\soc_I.clint_I.mtime[16] ));
 sg13g2_dfrbp_1 _35057_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net230),
    .D(net4498),
    .Q_N(_00022_),
    .Q(\soc_I.clint_I.mtime[17] ));
 sg13g2_dfrbp_1 _35058_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net228),
    .D(_01650_),
    .Q_N(_00030_),
    .Q(\soc_I.clint_I.mtime[18] ));
 sg13g2_dfrbp_1 _35059_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net226),
    .D(net3944),
    .Q_N(_00038_),
    .Q(\soc_I.clint_I.mtime[19] ));
 sg13g2_dfrbp_1 _35060_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net224),
    .D(net5120),
    .Q_N(_00045_),
    .Q(\soc_I.clint_I.mtime[20] ));
 sg13g2_dfrbp_1 _35061_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net222),
    .D(net5004),
    .Q_N(_00052_),
    .Q(\soc_I.clint_I.mtime[21] ));
 sg13g2_dfrbp_1 _35062_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net220),
    .D(_01654_),
    .Q_N(_00060_),
    .Q(\soc_I.clint_I.mtime[22] ));
 sg13g2_dfrbp_1 _35063_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net218),
    .D(net4726),
    .Q_N(_00068_),
    .Q(\soc_I.clint_I.mtime[23] ));
 sg13g2_dfrbp_1 _35064_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net216),
    .D(_01656_),
    .Q_N(_00018_),
    .Q(\soc_I.clint_I.mtime[24] ));
 sg13g2_dfrbp_1 _35065_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net214),
    .D(net4173),
    .Q_N(_00026_),
    .Q(\soc_I.clint_I.mtime[25] ));
 sg13g2_dfrbp_1 _35066_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net212),
    .D(net5196),
    .Q_N(_00034_),
    .Q(\soc_I.clint_I.mtime[26] ));
 sg13g2_dfrbp_1 _35067_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net210),
    .D(net4902),
    .Q_N(_00042_),
    .Q(\soc_I.clint_I.mtime[27] ));
 sg13g2_dfrbp_1 _35068_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net208),
    .D(_01660_),
    .Q_N(_00048_),
    .Q(\soc_I.clint_I.mtime[28] ));
 sg13g2_dfrbp_1 _35069_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net206),
    .D(net4556),
    .Q_N(_00056_),
    .Q(\soc_I.clint_I.mtime[29] ));
 sg13g2_dfrbp_1 _35070_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net204),
    .D(_01662_),
    .Q_N(_00064_),
    .Q(\soc_I.clint_I.mtime[30] ));
 sg13g2_dfrbp_1 _35071_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net202),
    .D(net4583),
    .Q_N(_00073_),
    .Q(\soc_I.clint_I.mtime[31] ));
 sg13g2_dfrbp_1 _35072_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net200),
    .D(_01664_),
    .Q_N(_00112_),
    .Q(\soc_I.clint_I.mtime[32] ));
 sg13g2_dfrbp_1 _35073_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net198),
    .D(net4496),
    .Q_N(_15459_),
    .Q(\soc_I.clint_I.mtime[33] ));
 sg13g2_dfrbp_1 _35074_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net196),
    .D(net4998),
    .Q_N(_15458_),
    .Q(\soc_I.clint_I.mtime[34] ));
 sg13g2_dfrbp_1 _35075_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net194),
    .D(net5538),
    .Q_N(_15457_),
    .Q(\soc_I.clint_I.mtime[35] ));
 sg13g2_dfrbp_1 _35076_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net192),
    .D(net5547),
    .Q_N(_15456_),
    .Q(\soc_I.clint_I.mtime[36] ));
 sg13g2_dfrbp_1 _35077_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net190),
    .D(net5167),
    .Q_N(_15455_),
    .Q(\soc_I.clint_I.mtime[37] ));
 sg13g2_dfrbp_1 _35078_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net188),
    .D(net5483),
    .Q_N(_15454_),
    .Q(\soc_I.clint_I.mtime[38] ));
 sg13g2_dfrbp_1 _35079_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net186),
    .D(_01671_),
    .Q_N(_15453_),
    .Q(\soc_I.clint_I.mtime[39] ));
 sg13g2_dfrbp_1 _35080_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net184),
    .D(_01672_),
    .Q_N(_15452_),
    .Q(\soc_I.clint_I.mtime[40] ));
 sg13g2_dfrbp_1 _35081_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net182),
    .D(net5318),
    .Q_N(_15451_),
    .Q(\soc_I.clint_I.mtime[41] ));
 sg13g2_dfrbp_1 _35082_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net180),
    .D(_01674_),
    .Q_N(_15450_),
    .Q(\soc_I.clint_I.mtime[42] ));
 sg13g2_dfrbp_1 _35083_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net178),
    .D(_01675_),
    .Q_N(_15449_),
    .Q(\soc_I.clint_I.mtime[43] ));
 sg13g2_dfrbp_1 _35084_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net176),
    .D(net5170),
    .Q_N(_15448_),
    .Q(\soc_I.clint_I.mtime[44] ));
 sg13g2_dfrbp_1 _35085_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net174),
    .D(net5500),
    .Q_N(_15447_),
    .Q(\soc_I.clint_I.mtime[45] ));
 sg13g2_dfrbp_1 _35086_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net172),
    .D(net5553),
    .Q_N(_15446_),
    .Q(\soc_I.clint_I.mtime[46] ));
 sg13g2_dfrbp_1 _35087_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net170),
    .D(_01679_),
    .Q_N(_15445_),
    .Q(\soc_I.clint_I.mtime[47] ));
 sg13g2_dfrbp_1 _35088_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net168),
    .D(_01680_),
    .Q_N(_15444_),
    .Q(\soc_I.clint_I.mtime[48] ));
 sg13g2_dfrbp_1 _35089_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net166),
    .D(_01681_),
    .Q_N(_15443_),
    .Q(\soc_I.clint_I.mtime[49] ));
 sg13g2_dfrbp_1 _35090_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net164),
    .D(net5445),
    .Q_N(_15442_),
    .Q(\soc_I.clint_I.mtime[50] ));
 sg13g2_dfrbp_1 _35091_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net162),
    .D(_01683_),
    .Q_N(_15441_),
    .Q(\soc_I.clint_I.mtime[51] ));
 sg13g2_dfrbp_1 _35092_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net160),
    .D(_01684_),
    .Q_N(_15440_),
    .Q(\soc_I.clint_I.mtime[52] ));
 sg13g2_dfrbp_1 _35093_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net158),
    .D(_01685_),
    .Q_N(_15439_),
    .Q(\soc_I.clint_I.mtime[53] ));
 sg13g2_dfrbp_1 _35094_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net156),
    .D(net4276),
    .Q_N(_15438_),
    .Q(\soc_I.clint_I.mtime[54] ));
 sg13g2_dfrbp_1 _35095_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net154),
    .D(_01687_),
    .Q_N(_15437_),
    .Q(\soc_I.clint_I.mtime[55] ));
 sg13g2_dfrbp_1 _35096_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net152),
    .D(_01688_),
    .Q_N(_15436_),
    .Q(\soc_I.clint_I.mtime[56] ));
 sg13g2_dfrbp_1 _35097_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net150),
    .D(_01689_),
    .Q_N(_15435_),
    .Q(\soc_I.clint_I.mtime[57] ));
 sg13g2_dfrbp_1 _35098_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net148),
    .D(_01690_),
    .Q_N(_15434_),
    .Q(\soc_I.clint_I.mtime[58] ));
 sg13g2_dfrbp_1 _35099_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net146),
    .D(net4827),
    .Q_N(_15433_),
    .Q(\soc_I.clint_I.mtime[59] ));
 sg13g2_dfrbp_1 _35100_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net144),
    .D(net4306),
    .Q_N(_15432_),
    .Q(\soc_I.clint_I.mtime[60] ));
 sg13g2_dfrbp_1 _35101_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net142),
    .D(_01693_),
    .Q_N(_15431_),
    .Q(\soc_I.clint_I.mtime[61] ));
 sg13g2_dfrbp_1 _35102_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net140),
    .D(net4565),
    .Q_N(_15430_),
    .Q(\soc_I.clint_I.mtime[62] ));
 sg13g2_dfrbp_1 _35103_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net138),
    .D(net4777),
    .Q_N(_15429_),
    .Q(\soc_I.clint_I.mtime[63] ));
 sg13g2_dfrbp_1 _35104_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net136),
    .D(_01696_),
    .Q_N(_15428_),
    .Q(\gpio_uo_out[0] ));
 sg13g2_dfrbp_1 _35105_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net134),
    .D(_01697_),
    .Q_N(_15427_),
    .Q(\gpio_uo_out[1] ));
 sg13g2_dfrbp_1 _35106_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net132),
    .D(_01698_),
    .Q_N(_15426_),
    .Q(\gpio_uo_out[2] ));
 sg13g2_dfrbp_1 _35107_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net130),
    .D(_01699_),
    .Q_N(_15425_),
    .Q(\gpio_uo_out[3] ));
 sg13g2_dfrbp_1 _35108_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net128),
    .D(_01700_),
    .Q_N(_15424_),
    .Q(\gpio_uo_out[4] ));
 sg13g2_dfrbp_1 _35109_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net126),
    .D(_01701_),
    .Q_N(_15423_),
    .Q(\gpio_uo_out[5] ));
 sg13g2_dfrbp_1 _35110_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net124),
    .D(_01702_),
    .Q_N(_15422_),
    .Q(\gpio_uo_out[6] ));
 sg13g2_dfrbp_1 _35111_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net122),
    .D(_01703_),
    .Q_N(_15421_),
    .Q(\gpio_uo_out[7] ));
 sg13g2_dfrbp_1 _35112_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net120),
    .D(_01704_),
    .Q_N(_15420_),
    .Q(\soc_I.clint_I.ready ));
 sg13g2_dfrbp_1 _35113_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net119),
    .D(_01705_),
    .Q_N(_15419_),
    .Q(\gpio_uo_en[0] ));
 sg13g2_dfrbp_1 _35114_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net117),
    .D(_01706_),
    .Q_N(_15418_),
    .Q(\gpio_uo_en[1] ));
 sg13g2_dfrbp_1 _35115_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net115),
    .D(_01707_),
    .Q_N(_15417_),
    .Q(\gpio_uo_en[2] ));
 sg13g2_dfrbp_1 _35116_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net113),
    .D(_01708_),
    .Q_N(_15416_),
    .Q(\gpio_uo_en[3] ));
 sg13g2_dfrbp_1 _35117_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net111),
    .D(_01709_),
    .Q_N(_15415_),
    .Q(\gpio_uo_en[4] ));
 sg13g2_dfrbp_1 _35118_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net109),
    .D(_01710_),
    .Q_N(_15414_),
    .Q(\gpio_uo_en[5] ));
 sg13g2_dfrbp_1 _35119_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net107),
    .D(_01711_),
    .Q_N(_15413_),
    .Q(\gpio_uo_en[6] ));
 sg13g2_dfrbp_1 _35120_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net105),
    .D(_01712_),
    .Q_N(_15412_),
    .Q(\gpio_uo_en[7] ));
 sg13g2_dfrbp_1 _35121_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net103),
    .D(_01713_),
    .Q_N(_15411_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][0] ));
 sg13g2_dfrbp_1 _35122_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net102),
    .D(_01714_),
    .Q_N(_15410_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][1] ));
 sg13g2_dfrbp_1 _35123_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net101),
    .D(_01715_),
    .Q_N(_15409_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][2] ));
 sg13g2_dfrbp_1 _35124_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net100),
    .D(_01716_),
    .Q_N(_15408_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][3] ));
 sg13g2_dfrbp_1 _35125_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net99),
    .D(_01717_),
    .Q_N(_15407_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][4] ));
 sg13g2_dfrbp_1 _35126_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net98),
    .D(_01718_),
    .Q_N(_15406_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][5] ));
 sg13g2_dfrbp_1 _35127_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net97),
    .D(_01719_),
    .Q_N(_15405_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][6] ));
 sg13g2_dfrbp_1 _35128_ (.CLK(clknet_leaf_304_clk),
    .RESET_B(net96),
    .D(_01720_),
    .Q_N(_15404_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][7] ));
 sg13g2_dfrbp_1 _35129_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net95),
    .D(_01721_),
    .Q_N(_15403_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][8] ));
 sg13g2_dfrbp_1 _35130_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net94),
    .D(_01722_),
    .Q_N(_15402_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][9] ));
 sg13g2_dfrbp_1 _35131_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net93),
    .D(_01723_),
    .Q_N(_15401_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][10] ));
 sg13g2_dfrbp_1 _35132_ (.CLK(clknet_leaf_318_clk),
    .RESET_B(net92),
    .D(_01724_),
    .Q_N(_15400_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][11] ));
 sg13g2_dfrbp_1 _35133_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net91),
    .D(_01725_),
    .Q_N(_15399_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][12] ));
 sg13g2_dfrbp_1 _35134_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net90),
    .D(_01726_),
    .Q_N(_15398_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][13] ));
 sg13g2_dfrbp_1 _35135_ (.CLK(clknet_leaf_289_clk),
    .RESET_B(net89),
    .D(_01727_),
    .Q_N(_15397_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][14] ));
 sg13g2_dfrbp_1 _35136_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net88),
    .D(net3826),
    .Q_N(_15396_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][15] ));
 sg13g2_dfrbp_1 _35137_ (.CLK(clknet_leaf_318_clk),
    .RESET_B(net87),
    .D(_01729_),
    .Q_N(_15395_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][16] ));
 sg13g2_dfrbp_1 _35138_ (.CLK(clknet_leaf_312_clk),
    .RESET_B(net86),
    .D(_01730_),
    .Q_N(_15394_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][17] ));
 sg13g2_dfrbp_1 _35139_ (.CLK(clknet_leaf_302_clk),
    .RESET_B(net85),
    .D(_01731_),
    .Q_N(_15393_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][18] ));
 sg13g2_dfrbp_1 _35140_ (.CLK(clknet_leaf_301_clk),
    .RESET_B(net84),
    .D(_01732_),
    .Q_N(_15392_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][19] ));
 sg13g2_dfrbp_1 _35141_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net83),
    .D(_01733_),
    .Q_N(_15391_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][20] ));
 sg13g2_dfrbp_1 _35142_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net82),
    .D(_01734_),
    .Q_N(_15390_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][21] ));
 sg13g2_dfrbp_1 _35143_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net81),
    .D(_01735_),
    .Q_N(_15389_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][22] ));
 sg13g2_dfrbp_1 _35144_ (.CLK(clknet_leaf_315_clk),
    .RESET_B(net80),
    .D(_01736_),
    .Q_N(_15388_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][23] ));
 sg13g2_dfrbp_1 _35145_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net79),
    .D(_01737_),
    .Q_N(_15387_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][24] ));
 sg13g2_dfrbp_1 _35146_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net78),
    .D(_01738_),
    .Q_N(_15386_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][25] ));
 sg13g2_dfrbp_1 _35147_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net77),
    .D(_01739_),
    .Q_N(_15385_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][26] ));
 sg13g2_dfrbp_1 _35148_ (.CLK(clknet_leaf_277_clk),
    .RESET_B(net76),
    .D(_01740_),
    .Q_N(_15384_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][27] ));
 sg13g2_dfrbp_1 _35149_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net75),
    .D(_01741_),
    .Q_N(_15383_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][28] ));
 sg13g2_dfrbp_1 _35150_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net74),
    .D(_01742_),
    .Q_N(_15382_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][29] ));
 sg13g2_dfrbp_1 _35151_ (.CLK(clknet_leaf_291_clk),
    .RESET_B(net73),
    .D(_01743_),
    .Q_N(_15381_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][30] ));
 sg13g2_dfrbp_1 _35152_ (.CLK(clknet_leaf_307_clk),
    .RESET_B(net72),
    .D(_01744_),
    .Q_N(_15380_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][31] ));
 sg13g2_dfrbp_1 _35153_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net71),
    .D(_01745_),
    .Q_N(_15379_),
    .Q(\soc_I.spi0_I.sclk ));
 sg13g2_dfrbp_1 _35154_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net69),
    .D(_01746_),
    .Q_N(_15378_),
    .Q(\soc_I.spi0_I.xfer_cycles[0] ));
 sg13g2_dfrbp_1 _35155_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net67),
    .D(_01747_),
    .Q_N(_15377_),
    .Q(\soc_I.spi0_I.xfer_cycles[1] ));
 sg13g2_dfrbp_1 _35156_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net65),
    .D(net4677),
    .Q_N(_15376_),
    .Q(\soc_I.spi0_I.xfer_cycles[2] ));
 sg13g2_dfrbp_1 _35157_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net63),
    .D(net3191),
    .Q_N(_15375_),
    .Q(\soc_I.spi0_I.xfer_cycles[3] ));
 sg13g2_dfrbp_1 _35158_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net61),
    .D(net4293),
    .Q_N(_00148_),
    .Q(\soc_I.spi0_I.xfer_cycles[4] ));
 sg13g2_dfrbp_1 _35159_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net59),
    .D(net4740),
    .Q_N(_15374_),
    .Q(\soc_I.spi0_I.xfer_cycles[5] ));
 sg13g2_dfrbp_1 _35160_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net57),
    .D(_01752_),
    .Q_N(_15373_),
    .Q(\soc_I.spi0_I.ready_xfer ));
 sg13g2_dfrbp_1 _35161_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net55),
    .D(net2840),
    .Q_N(_15372_),
    .Q(\soc_I.spi0_I.sio0_si_mosi ));
 sg13g2_dfrbp_1 _35162_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net53),
    .D(_01754_),
    .Q_N(_00286_),
    .Q(\soc_I.spi0_I.state ));
 sg13g2_dfrbp_1 _35163_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net51),
    .D(_01755_),
    .Q_N(_15371_),
    .Q(\soc_I.spi0_I.spi_buf[0] ));
 sg13g2_dfrbp_1 _35164_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net49),
    .D(_01756_),
    .Q_N(_15370_),
    .Q(\soc_I.spi0_I.spi_buf[1] ));
 sg13g2_dfrbp_1 _35165_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net47),
    .D(_01757_),
    .Q_N(_15369_),
    .Q(\soc_I.spi0_I.spi_buf[2] ));
 sg13g2_dfrbp_1 _35166_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net45),
    .D(_01758_),
    .Q_N(_15368_),
    .Q(\soc_I.spi0_I.spi_buf[3] ));
 sg13g2_dfrbp_1 _35167_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net43),
    .D(_01759_),
    .Q_N(_15367_),
    .Q(\soc_I.spi0_I.spi_buf[4] ));
 sg13g2_dfrbp_1 _35168_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net41),
    .D(_01760_),
    .Q_N(_15366_),
    .Q(\soc_I.spi0_I.spi_buf[5] ));
 sg13g2_dfrbp_1 _35169_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net39),
    .D(_01761_),
    .Q_N(_15365_),
    .Q(\soc_I.spi0_I.spi_buf[6] ));
 sg13g2_dfrbp_1 _35170_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net37),
    .D(_01762_),
    .Q_N(_15364_),
    .Q(\soc_I.spi0_I.spi_buf[7] ));
 sg13g2_dfrbp_1 _35171_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net35),
    .D(net2599),
    .Q_N(_00301_),
    .Q(\soc_I.spi0_I.tick_cnt[0] ));
 sg13g2_dfrbp_1 _35172_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net33),
    .D(_01764_),
    .Q_N(_15363_),
    .Q(\soc_I.spi0_I.tick_cnt[1] ));
 sg13g2_dfrbp_1 _35173_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net31),
    .D(net3821),
    .Q_N(_15362_),
    .Q(\soc_I.spi0_I.tick_cnt[2] ));
 sg13g2_dfrbp_1 _35174_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net29),
    .D(_01766_),
    .Q_N(_15361_),
    .Q(\soc_I.spi0_I.tick_cnt[3] ));
 sg13g2_dfrbp_1 _35175_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net27),
    .D(_01767_),
    .Q_N(_15360_),
    .Q(\soc_I.spi0_I.tick_cnt[4] ));
 sg13g2_dfrbp_1 _35176_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net25),
    .D(_01768_),
    .Q_N(_15359_),
    .Q(\soc_I.spi0_I.tick_cnt[5] ));
 sg13g2_dfrbp_1 _35177_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net23),
    .D(net3427),
    .Q_N(_15358_),
    .Q(\soc_I.spi0_I.tick_cnt[6] ));
 sg13g2_dfrbp_1 _35178_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net21),
    .D(_01770_),
    .Q_N(_15357_),
    .Q(\soc_I.spi0_I.tick_cnt[7] ));
 sg13g2_dfrbp_1 _35179_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net19),
    .D(_01771_),
    .Q_N(_15356_),
    .Q(\soc_I.spi0_I.tick_cnt[8] ));
 sg13g2_dfrbp_1 _35180_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net17),
    .D(_01772_),
    .Q_N(_15355_),
    .Q(\soc_I.spi0_I.tick_cnt[9] ));
 sg13g2_dfrbp_1 _35181_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net15),
    .D(_01773_),
    .Q_N(_15354_),
    .Q(\soc_I.spi0_I.tick_cnt[10] ));
 sg13g2_dfrbp_1 _35182_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net2593),
    .D(_01774_),
    .Q_N(_15353_),
    .Q(\soc_I.spi0_I.tick_cnt[11] ));
 sg13g2_dfrbp_1 _35183_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net2591),
    .D(_01775_),
    .Q_N(_15352_),
    .Q(\soc_I.spi0_I.tick_cnt[12] ));
 sg13g2_dfrbp_1 _35184_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net2589),
    .D(_01776_),
    .Q_N(_15351_),
    .Q(\soc_I.spi0_I.tick_cnt[13] ));
 sg13g2_dfrbp_1 _35185_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net2587),
    .D(_01777_),
    .Q_N(_15350_),
    .Q(\soc_I.spi0_I.tick_cnt[14] ));
 sg13g2_dfrbp_1 _35186_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net2585),
    .D(_01778_),
    .Q_N(_15349_),
    .Q(\soc_I.spi0_I.tick_cnt[15] ));
 sg13g2_dfrbp_1 _35187_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net2583),
    .D(_01779_),
    .Q_N(_15348_),
    .Q(\soc_I.spi0_I.tick_cnt[16] ));
 sg13g2_dfrbp_1 _35188_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net2581),
    .D(_01780_),
    .Q_N(_15347_),
    .Q(\soc_I.spi0_I.tick_cnt[17] ));
 sg13g2_dfrbp_1 _35189_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net2579),
    .D(_01781_),
    .Q_N(_00108_),
    .Q(\soc_I.spi0_I.cen ));
 sg13g2_dfrbp_1 _35190_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net2577),
    .D(net4165),
    .Q_N(_00149_),
    .Q(\soc_I.rx_uart_i.fifo_i.cnt[0] ));
 sg13g2_dfrbp_1 _35191_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net2576),
    .D(net5205),
    .Q_N(_15346_),
    .Q(\soc_I.rx_uart_i.fifo_i.cnt[1] ));
 sg13g2_dfrbp_1 _35192_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net2575),
    .D(_01784_),
    .Q_N(_15345_),
    .Q(\soc_I.rx_uart_i.fifo_i.cnt[2] ));
 sg13g2_dfrbp_1 _35193_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net2574),
    .D(_01785_),
    .Q_N(_15344_),
    .Q(\soc_I.rx_uart_i.fifo_i.cnt[3] ));
 sg13g2_dfrbp_1 _35194_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net2573),
    .D(_01786_),
    .Q_N(_15343_),
    .Q(\soc_I.rx_uart_i.fifo_i.cnt[4] ));
 sg13g2_dfrbp_1 _35195_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net2572),
    .D(net4217),
    .Q_N(_15342_),
    .Q(\soc_I.gpio0_I.rdata[0] ));
 sg13g2_dfrbp_1 _35196_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net2570),
    .D(net3406),
    .Q_N(_15341_),
    .Q(\soc_I.gpio0_I.rdata[1] ));
 sg13g2_dfrbp_1 _35197_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net2568),
    .D(net4641),
    .Q_N(_15340_),
    .Q(\soc_I.gpio0_I.rdata[2] ));
 sg13g2_dfrbp_1 _35198_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net2566),
    .D(net4635),
    .Q_N(_15339_),
    .Q(\soc_I.gpio0_I.rdata[3] ));
 sg13g2_dfrbp_1 _35199_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net2564),
    .D(net3919),
    .Q_N(_15338_),
    .Q(\soc_I.gpio0_I.rdata[4] ));
 sg13g2_dfrbp_1 _35200_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net2562),
    .D(net3803),
    .Q_N(_15337_),
    .Q(\soc_I.gpio0_I.rdata[5] ));
 sg13g2_dfrbp_1 _35201_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net2560),
    .D(net4278),
    .Q_N(_15336_),
    .Q(\soc_I.gpio0_I.rdata[6] ));
 sg13g2_dfrbp_1 _35202_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net2558),
    .D(net4062),
    .Q_N(_15335_),
    .Q(\soc_I.gpio0_I.rdata[7] ));
 sg13g2_dfrbp_1 _35203_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net2556),
    .D(net5216),
    .Q_N(_15334_),
    .Q(\soc_I.rx_uart_i.ready ));
 sg13g2_dfrbp_1 _35204_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2554),
    .D(net2860),
    .Q_N(_15333_),
    .Q(\soc_I.qqspi_I.rdata[0] ));
 sg13g2_dfrbp_1 _35205_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net2553),
    .D(net2850),
    .Q_N(_15332_),
    .Q(\soc_I.qqspi_I.rdata[1] ));
 sg13g2_dfrbp_1 _35206_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2552),
    .D(net2678),
    .Q_N(_15331_),
    .Q(\soc_I.qqspi_I.rdata[2] ));
 sg13g2_dfrbp_1 _35207_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net2551),
    .D(net3445),
    .Q_N(_15330_),
    .Q(\soc_I.qqspi_I.rdata[3] ));
 sg13g2_dfrbp_1 _35208_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net2550),
    .D(net2814),
    .Q_N(_15329_),
    .Q(\soc_I.qqspi_I.rdata[4] ));
 sg13g2_dfrbp_1 _35209_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net2549),
    .D(net2784),
    .Q_N(_15328_),
    .Q(\soc_I.qqspi_I.rdata[5] ));
 sg13g2_dfrbp_1 _35210_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net2548),
    .D(net2698),
    .Q_N(_15327_),
    .Q(\soc_I.qqspi_I.rdata[6] ));
 sg13g2_dfrbp_1 _35211_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net2547),
    .D(net2950),
    .Q_N(_15326_),
    .Q(\soc_I.qqspi_I.rdata[7] ));
 sg13g2_dfrbp_1 _35212_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2546),
    .D(net3746),
    .Q_N(_15325_),
    .Q(\soc_I.qqspi_I.rdata[8] ));
 sg13g2_dfrbp_1 _35213_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2545),
    .D(net3884),
    .Q_N(_15324_),
    .Q(\soc_I.qqspi_I.rdata[9] ));
 sg13g2_dfrbp_1 _35214_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2544),
    .D(net3977),
    .Q_N(_15323_),
    .Q(\soc_I.qqspi_I.rdata[10] ));
 sg13g2_dfrbp_1 _35215_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2543),
    .D(net2655),
    .Q_N(_15322_),
    .Q(\soc_I.qqspi_I.rdata[11] ));
 sg13g2_dfrbp_1 _35216_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2542),
    .D(net3652),
    .Q_N(_15321_),
    .Q(\soc_I.qqspi_I.rdata[12] ));
 sg13g2_dfrbp_1 _35217_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2541),
    .D(net3146),
    .Q_N(_15320_),
    .Q(\soc_I.qqspi_I.rdata[13] ));
 sg13g2_dfrbp_1 _35218_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2540),
    .D(net4167),
    .Q_N(_15319_),
    .Q(\soc_I.qqspi_I.rdata[14] ));
 sg13g2_dfrbp_1 _35219_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2539),
    .D(net2641),
    .Q_N(_15318_),
    .Q(\soc_I.qqspi_I.rdata[15] ));
 sg13g2_dfrbp_1 _35220_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2538),
    .D(net2706),
    .Q_N(_15317_),
    .Q(\soc_I.qqspi_I.rdata[16] ));
 sg13g2_dfrbp_1 _35221_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2537),
    .D(net3495),
    .Q_N(_15316_),
    .Q(\soc_I.qqspi_I.rdata[17] ));
 sg13g2_dfrbp_1 _35222_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2536),
    .D(net2782),
    .Q_N(_15315_),
    .Q(\soc_I.qqspi_I.rdata[18] ));
 sg13g2_dfrbp_1 _35223_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2535),
    .D(net2720),
    .Q_N(_15314_),
    .Q(\soc_I.qqspi_I.rdata[19] ));
 sg13g2_dfrbp_1 _35224_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2534),
    .D(net3630),
    .Q_N(_15313_),
    .Q(\soc_I.qqspi_I.rdata[20] ));
 sg13g2_dfrbp_1 _35225_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2533),
    .D(net2768),
    .Q_N(_15312_),
    .Q(\soc_I.qqspi_I.rdata[21] ));
 sg13g2_dfrbp_1 _35226_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2532),
    .D(net3086),
    .Q_N(_15311_),
    .Q(\soc_I.qqspi_I.rdata[22] ));
 sg13g2_dfrbp_1 _35227_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2531),
    .D(net4383),
    .Q_N(_15310_),
    .Q(\soc_I.qqspi_I.rdata[23] ));
 sg13g2_dfrbp_1 _35228_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net2530),
    .D(net3093),
    .Q_N(_15309_),
    .Q(\soc_I.qqspi_I.rdata[24] ));
 sg13g2_dfrbp_1 _35229_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net2529),
    .D(net2670),
    .Q_N(_15308_),
    .Q(\soc_I.qqspi_I.rdata[25] ));
 sg13g2_dfrbp_1 _35230_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net2528),
    .D(net2780),
    .Q_N(_15307_),
    .Q(\soc_I.qqspi_I.rdata[26] ));
 sg13g2_dfrbp_1 _35231_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net2527),
    .D(net2691),
    .Q_N(_15306_),
    .Q(\soc_I.qqspi_I.rdata[27] ));
 sg13g2_dfrbp_1 _35232_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net2526),
    .D(net2694),
    .Q_N(_15305_),
    .Q(\soc_I.qqspi_I.rdata[28] ));
 sg13g2_dfrbp_1 _35233_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net2525),
    .D(net2857),
    .Q_N(_15304_),
    .Q(\soc_I.qqspi_I.rdata[29] ));
 sg13g2_dfrbp_1 _35234_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net2524),
    .D(net2774),
    .Q_N(_15303_),
    .Q(\soc_I.qqspi_I.rdata[30] ));
 sg13g2_dfrbp_1 _35235_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net2523),
    .D(net2791),
    .Q_N(_15302_),
    .Q(\soc_I.qqspi_I.rdata[31] ));
 sg13g2_dfrbp_1 _35236_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net2522),
    .D(net5144),
    .Q_N(_15301_),
    .Q(\soc_I.rx_uart_i.fifo_i.din[0] ));
 sg13g2_dfrbp_1 _35237_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net2520),
    .D(_01829_),
    .Q_N(_15300_),
    .Q(\soc_I.rx_uart_i.fifo_i.din[1] ));
 sg13g2_dfrbp_1 _35238_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net2518),
    .D(_01830_),
    .Q_N(_15299_),
    .Q(\soc_I.rx_uart_i.fifo_i.din[2] ));
 sg13g2_dfrbp_1 _35239_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net2516),
    .D(_01831_),
    .Q_N(_15298_),
    .Q(\soc_I.rx_uart_i.fifo_i.din[3] ));
 sg13g2_dfrbp_1 _35240_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net2514),
    .D(_01832_),
    .Q_N(_15297_),
    .Q(\soc_I.rx_uart_i.fifo_i.din[4] ));
 sg13g2_dfrbp_1 _35241_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net2512),
    .D(_01833_),
    .Q_N(_15296_),
    .Q(\soc_I.rx_uart_i.fifo_i.din[5] ));
 sg13g2_dfrbp_1 _35242_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net2510),
    .D(_01834_),
    .Q_N(_15295_),
    .Q(\soc_I.rx_uart_i.fifo_i.din[6] ));
 sg13g2_dfrbp_1 _35243_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net2508),
    .D(_01835_),
    .Q_N(_15294_),
    .Q(\soc_I.rx_uart_i.fifo_i.din[7] ));
 sg13g2_dfrbp_1 _35244_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2506),
    .D(_01836_),
    .Q_N(_15293_),
    .Q(\soc_I.rx_uart_i.state[0] ));
 sg13g2_dfrbp_1 _35245_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2504),
    .D(_01837_),
    .Q_N(_15292_),
    .Q(\soc_I.rx_uart_i.state[1] ));
 sg13g2_dfrbp_1 _35246_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2502),
    .D(_01838_),
    .Q_N(_00249_),
    .Q(\soc_I.rx_uart_i.state[2] ));
 sg13g2_dfrbp_1 _35247_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net2500),
    .D(net3096),
    .Q_N(_00300_),
    .Q(\soc_I.rx_uart_i.bit_idx[0] ));
 sg13g2_dfrbp_1 _35248_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net2498),
    .D(_01840_),
    .Q_N(_15291_),
    .Q(\soc_I.rx_uart_i.bit_idx[1] ));
 sg13g2_dfrbp_1 _35249_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net2496),
    .D(_01841_),
    .Q_N(_15290_),
    .Q(\soc_I.rx_uart_i.bit_idx[2] ));
 sg13g2_dfrbp_1 _35250_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2494),
    .D(net5221),
    .Q_N(_15289_),
    .Q(\soc_I.rx_uart_i.wait_states[0] ));
 sg13g2_dfrbp_1 _35251_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2492),
    .D(net5247),
    .Q_N(_15288_),
    .Q(\soc_I.rx_uart_i.wait_states[1] ));
 sg13g2_dfrbp_1 _35252_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2490),
    .D(net4535),
    .Q_N(_00153_),
    .Q(\soc_I.rx_uart_i.wait_states[2] ));
 sg13g2_dfrbp_1 _35253_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2488),
    .D(_01845_),
    .Q_N(_15287_),
    .Q(\soc_I.rx_uart_i.wait_states[3] ));
 sg13g2_dfrbp_1 _35254_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2486),
    .D(net5016),
    .Q_N(_00154_),
    .Q(\soc_I.rx_uart_i.wait_states[4] ));
 sg13g2_dfrbp_1 _35255_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2484),
    .D(_01847_),
    .Q_N(_15286_),
    .Q(\soc_I.rx_uart_i.wait_states[5] ));
 sg13g2_dfrbp_1 _35256_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2482),
    .D(net4889),
    .Q_N(_00155_),
    .Q(\soc_I.rx_uart_i.wait_states[6] ));
 sg13g2_dfrbp_1 _35257_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2480),
    .D(net5163),
    .Q_N(_15285_),
    .Q(\soc_I.rx_uart_i.wait_states[7] ));
 sg13g2_dfrbp_1 _35258_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2478),
    .D(net4851),
    .Q_N(_15284_),
    .Q(\soc_I.rx_uart_i.wait_states[8] ));
 sg13g2_dfrbp_1 _35259_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2476),
    .D(net5110),
    .Q_N(_15283_),
    .Q(\soc_I.rx_uart_i.wait_states[9] ));
 sg13g2_dfrbp_1 _35260_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2474),
    .D(net4760),
    .Q_N(_00156_),
    .Q(\soc_I.rx_uart_i.wait_states[10] ));
 sg13g2_dfrbp_1 _35261_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2472),
    .D(_01853_),
    .Q_N(_15282_),
    .Q(\soc_I.rx_uart_i.wait_states[11] ));
 sg13g2_dfrbp_1 _35262_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2470),
    .D(_01854_),
    .Q_N(_15281_),
    .Q(\soc_I.rx_uart_i.wait_states[12] ));
 sg13g2_dfrbp_1 _35263_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2468),
    .D(net5178),
    .Q_N(_15280_),
    .Q(\soc_I.rx_uart_i.wait_states[13] ));
 sg13g2_dfrbp_1 _35264_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2466),
    .D(net4867),
    .Q_N(_00157_),
    .Q(\soc_I.rx_uart_i.wait_states[14] ));
 sg13g2_dfrbp_1 _35265_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2464),
    .D(_01857_),
    .Q_N(_15279_),
    .Q(\soc_I.rx_uart_i.wait_states[15] ));
 sg13g2_dfrbp_1 _35266_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2462),
    .D(net2634),
    .Q_N(_00290_),
    .Q(\soc_I.rx_uart_i.wait_states[16] ));
 sg13g2_dfrbp_1 _35267_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net2460),
    .D(net2605),
    .Q_N(_00299_),
    .Q(\soc_I.rx_uart_i.fifo_i.wr_ptr[0] ));
 sg13g2_dfrbp_1 _35268_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net2458),
    .D(_01860_),
    .Q_N(_15278_),
    .Q(\soc_I.rx_uart_i.fifo_i.wr_ptr[1] ));
 sg13g2_dfrbp_1 _35269_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net2456),
    .D(_01861_),
    .Q_N(_15277_),
    .Q(\soc_I.rx_uart_i.fifo_i.wr_ptr[2] ));
 sg13g2_dfrbp_1 _35270_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net2454),
    .D(_01862_),
    .Q_N(_15276_),
    .Q(\soc_I.rx_uart_i.fifo_i.wr_ptr[3] ));
 sg13g2_dfrbp_1 _35271_ (.CLK(clknet_leaf_325_clk),
    .RESET_B(net2452),
    .D(net2607),
    .Q_N(_00298_),
    .Q(\soc_I.rx_uart_i.fifo_i.rd_ptr[0] ));
 sg13g2_dfrbp_1 _35272_ (.CLK(clknet_leaf_325_clk),
    .RESET_B(net2450),
    .D(net3909),
    .Q_N(_15275_),
    .Q(\soc_I.rx_uart_i.fifo_i.rd_ptr[1] ));
 sg13g2_dfrbp_1 _35273_ (.CLK(clknet_leaf_325_clk),
    .RESET_B(net2448),
    .D(_01865_),
    .Q_N(_15274_),
    .Q(\soc_I.rx_uart_i.fifo_i.rd_ptr[2] ));
 sg13g2_dfrbp_1 _35274_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net2446),
    .D(_01866_),
    .Q_N(_15273_),
    .Q(\soc_I.rx_uart_i.fifo_i.rd_ptr[3] ));
 sg13g2_dfrbp_1 _35275_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2444),
    .D(_01867_),
    .Q_N(_15272_),
    .Q(\soc_I.rx_uart_i.rx_in_sync[0] ));
 sg13g2_dfrbp_1 _35276_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2443),
    .D(_01868_),
    .Q_N(_15271_),
    .Q(\soc_I.rx_uart_i.rx_in_sync[1] ));
 sg13g2_dfrbp_1 _35277_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net2442),
    .D(_01869_),
    .Q_N(_00289_),
    .Q(\soc_I.rx_uart_i.rx_in_sync[2] ));
 sg13g2_dfrbp_1 _35278_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net2441),
    .D(net4283),
    .Q_N(_15270_),
    .Q(\soc_I.tx_uart_i.ready ));
 sg13g2_dfrbp_1 _35279_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net2439),
    .D(net5208),
    .Q_N(_15269_),
    .Q(\soc_I.tx_uart_i.tx_out ));
 sg13g2_dfrbp_1 _35280_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net2437),
    .D(_01872_),
    .Q_N(_15268_),
    .Q(\soc_I.spi0_I.ready_ctrl ));
 sg13g2_dfrbp_1 _35281_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net2436),
    .D(net2609),
    .Q_N(_00297_),
    .Q(\soc_I.tx_uart_i.bit_idx[0] ));
 sg13g2_dfrbp_1 _35282_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net2434),
    .D(_01874_),
    .Q_N(_15267_),
    .Q(\soc_I.tx_uart_i.bit_idx[1] ));
 sg13g2_dfrbp_1 _35283_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net2432),
    .D(_01875_),
    .Q_N(_00152_),
    .Q(\soc_I.tx_uart_i.bit_idx[2] ));
 sg13g2_dfrbp_1 _35284_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net2430),
    .D(_01876_),
    .Q_N(_15266_),
    .Q(\soc_I.tx_uart_i.tx_data_reg[0] ));
 sg13g2_dfrbp_1 _35285_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net2428),
    .D(_01877_),
    .Q_N(_15265_),
    .Q(\soc_I.tx_uart_i.tx_data_reg[1] ));
 sg13g2_dfrbp_1 _35286_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net2426),
    .D(_01878_),
    .Q_N(_15264_),
    .Q(\soc_I.tx_uart_i.tx_data_reg[2] ));
 sg13g2_dfrbp_1 _35287_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net2424),
    .D(_01879_),
    .Q_N(_15263_),
    .Q(\soc_I.tx_uart_i.tx_data_reg[3] ));
 sg13g2_dfrbp_1 _35288_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net2422),
    .D(net4046),
    .Q_N(_15262_),
    .Q(\soc_I.tx_uart_i.tx_data_reg[4] ));
 sg13g2_dfrbp_1 _35289_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net2420),
    .D(_01881_),
    .Q_N(_15261_),
    .Q(\soc_I.tx_uart_i.tx_data_reg[5] ));
 sg13g2_dfrbp_1 _35290_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net2418),
    .D(_01882_),
    .Q_N(_15260_),
    .Q(\soc_I.tx_uart_i.tx_data_reg[6] ));
 sg13g2_dfrbp_1 _35291_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net2416),
    .D(_01883_),
    .Q_N(_15259_),
    .Q(\soc_I.tx_uart_i.tx_data_reg[7] ));
 sg13g2_dfrbp_1 _35292_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net2414),
    .D(net2800),
    .Q_N(_15258_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[9][0] ));
 sg13g2_dfrbp_1 _35293_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net2413),
    .D(net4185),
    .Q_N(_15257_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[9][1] ));
 sg13g2_dfrbp_1 _35294_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net2412),
    .D(_01886_),
    .Q_N(_15256_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[9][2] ));
 sg13g2_dfrbp_1 _35295_ (.CLK(clknet_leaf_323_clk),
    .RESET_B(net2411),
    .D(_01887_),
    .Q_N(_15255_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[9][3] ));
 sg13g2_dfrbp_1 _35296_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net2410),
    .D(net3940),
    .Q_N(_15254_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[9][4] ));
 sg13g2_dfrbp_1 _35297_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net2409),
    .D(_01889_),
    .Q_N(_15253_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[9][5] ));
 sg13g2_dfrbp_1 _35298_ (.CLK(clknet_leaf_321_clk),
    .RESET_B(net2408),
    .D(net4151),
    .Q_N(_15252_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[9][6] ));
 sg13g2_dfrbp_1 _35299_ (.CLK(clknet_leaf_323_clk),
    .RESET_B(net2407),
    .D(_01891_),
    .Q_N(_15251_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[9][7] ));
 sg13g2_dfrbp_1 _35300_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2406),
    .D(_01892_),
    .Q_N(_15250_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][0] ));
 sg13g2_dfrbp_1 _35301_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2405),
    .D(_01893_),
    .Q_N(_15249_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][1] ));
 sg13g2_dfrbp_1 _35302_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2404),
    .D(_01894_),
    .Q_N(_15248_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][2] ));
 sg13g2_dfrbp_1 _35303_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2403),
    .D(_01895_),
    .Q_N(_15247_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][3] ));
 sg13g2_dfrbp_1 _35304_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2402),
    .D(_01896_),
    .Q_N(_15246_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][4] ));
 sg13g2_dfrbp_1 _35305_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2401),
    .D(_01897_),
    .Q_N(_15245_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][5] ));
 sg13g2_dfrbp_1 _35306_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2400),
    .D(_01898_),
    .Q_N(_15244_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][6] ));
 sg13g2_dfrbp_1 _35307_ (.CLK(clknet_leaf_305_clk),
    .RESET_B(net2399),
    .D(_01899_),
    .Q_N(_15243_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][7] ));
 sg13g2_dfrbp_1 _35308_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2398),
    .D(_01900_),
    .Q_N(_15242_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][8] ));
 sg13g2_dfrbp_1 _35309_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2397),
    .D(_01901_),
    .Q_N(_15241_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][9] ));
 sg13g2_dfrbp_1 _35310_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2396),
    .D(_01902_),
    .Q_N(_15240_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][10] ));
 sg13g2_dfrbp_1 _35311_ (.CLK(clknet_leaf_313_clk),
    .RESET_B(net2395),
    .D(_01903_),
    .Q_N(_15239_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][11] ));
 sg13g2_dfrbp_1 _35312_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2394),
    .D(_01904_),
    .Q_N(_15238_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][12] ));
 sg13g2_dfrbp_1 _35313_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2393),
    .D(_01905_),
    .Q_N(_15237_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][13] ));
 sg13g2_dfrbp_1 _35314_ (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2392),
    .D(_01906_),
    .Q_N(_15236_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][14] ));
 sg13g2_dfrbp_1 _35315_ (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2391),
    .D(_01907_),
    .Q_N(_15235_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][15] ));
 sg13g2_dfrbp_1 _35316_ (.CLK(clknet_leaf_317_clk),
    .RESET_B(net2390),
    .D(_01908_),
    .Q_N(_15234_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][16] ));
 sg13g2_dfrbp_1 _35317_ (.CLK(clknet_leaf_314_clk),
    .RESET_B(net2389),
    .D(_01909_),
    .Q_N(_15233_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][17] ));
 sg13g2_dfrbp_1 _35318_ (.CLK(clknet_leaf_306_clk),
    .RESET_B(net2388),
    .D(_01910_),
    .Q_N(_15232_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][18] ));
 sg13g2_dfrbp_1 _35319_ (.CLK(clknet_leaf_303_clk),
    .RESET_B(net2387),
    .D(_01911_),
    .Q_N(_15231_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][19] ));
 sg13g2_dfrbp_1 _35320_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net2386),
    .D(_01912_),
    .Q_N(_15230_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][20] ));
 sg13g2_dfrbp_1 _35321_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2385),
    .D(net3081),
    .Q_N(_15229_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][21] ));
 sg13g2_dfrbp_1 _35322_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2384),
    .D(_01914_),
    .Q_N(_15228_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][22] ));
 sg13g2_dfrbp_1 _35323_ (.CLK(clknet_leaf_306_clk),
    .RESET_B(net2383),
    .D(_01915_),
    .Q_N(_15227_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][23] ));
 sg13g2_dfrbp_1 _35324_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2382),
    .D(_01916_),
    .Q_N(_15226_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][24] ));
 sg13g2_dfrbp_1 _35325_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2381),
    .D(_01917_),
    .Q_N(_15225_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][25] ));
 sg13g2_dfrbp_1 _35326_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2380),
    .D(_01918_),
    .Q_N(_15224_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][26] ));
 sg13g2_dfrbp_1 _35327_ (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2379),
    .D(_01919_),
    .Q_N(_15223_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][27] ));
 sg13g2_dfrbp_1 _35328_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2378),
    .D(_01920_),
    .Q_N(_15222_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][28] ));
 sg13g2_dfrbp_1 _35329_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2377),
    .D(_01921_),
    .Q_N(_15221_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][29] ));
 sg13g2_dfrbp_1 _35330_ (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2376),
    .D(_01922_),
    .Q_N(_15220_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][30] ));
 sg13g2_dfrbp_1 _35331_ (.CLK(clknet_leaf_309_clk),
    .RESET_B(net2375),
    .D(_01923_),
    .Q_N(_15219_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][31] ));
 sg13g2_dfrbp_1 _35332_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net2374),
    .D(net4021),
    .Q_N(_15218_),
    .Q(\soc_I.tx_uart_i.wait_states[1] ));
 sg13g2_dfrbp_1 _35333_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net2373),
    .D(_01925_),
    .Q_N(_15217_),
    .Q(\soc_I.tx_uart_i.wait_states[2] ));
 sg13g2_dfrbp_1 _35334_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net2372),
    .D(_01926_),
    .Q_N(_15216_),
    .Q(\soc_I.tx_uart_i.wait_states[3] ));
 sg13g2_dfrbp_1 _35335_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net2371),
    .D(_01927_),
    .Q_N(_15215_),
    .Q(\soc_I.tx_uart_i.wait_states[4] ));
 sg13g2_dfrbp_1 _35336_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net2370),
    .D(net3616),
    .Q_N(_15214_),
    .Q(\soc_I.tx_uart_i.wait_states[5] ));
 sg13g2_dfrbp_1 _35337_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net2369),
    .D(_01929_),
    .Q_N(_15213_),
    .Q(\soc_I.tx_uart_i.wait_states[6] ));
 sg13g2_dfrbp_1 _35338_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net2368),
    .D(_01930_),
    .Q_N(_15212_),
    .Q(\soc_I.tx_uart_i.wait_states[7] ));
 sg13g2_dfrbp_1 _35339_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net2367),
    .D(_01931_),
    .Q_N(_15211_),
    .Q(\soc_I.tx_uart_i.wait_states[8] ));
 sg13g2_dfrbp_1 _35340_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2366),
    .D(net3931),
    .Q_N(_15210_),
    .Q(\soc_I.tx_uart_i.wait_states[9] ));
 sg13g2_dfrbp_1 _35341_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2365),
    .D(net3528),
    .Q_N(_15209_),
    .Q(\soc_I.tx_uart_i.wait_states[10] ));
 sg13g2_dfrbp_1 _35342_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2364),
    .D(_01934_),
    .Q_N(_15208_),
    .Q(\soc_I.tx_uart_i.wait_states[11] ));
 sg13g2_dfrbp_1 _35343_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2363),
    .D(_01935_),
    .Q_N(_15207_),
    .Q(\soc_I.tx_uart_i.wait_states[12] ));
 sg13g2_dfrbp_1 _35344_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net2362),
    .D(net4196),
    .Q_N(_15206_),
    .Q(\soc_I.tx_uart_i.wait_states[13] ));
 sg13g2_dfrbp_1 _35345_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net2361),
    .D(_01937_),
    .Q_N(_15205_),
    .Q(\soc_I.tx_uart_i.wait_states[14] ));
 sg13g2_dfrbp_1 _35346_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net2360),
    .D(_01938_),
    .Q_N(_15204_),
    .Q(\soc_I.tx_uart_i.wait_states[15] ));
 sg13g2_dfrbp_1 _35347_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2359),
    .D(_01939_),
    .Q_N(_15203_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][0] ));
 sg13g2_dfrbp_1 _35348_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2358),
    .D(_01940_),
    .Q_N(_15202_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][1] ));
 sg13g2_dfrbp_1 _35349_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2357),
    .D(_01941_),
    .Q_N(_15201_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][2] ));
 sg13g2_dfrbp_1 _35350_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2356),
    .D(_01942_),
    .Q_N(_15200_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][3] ));
 sg13g2_dfrbp_1 _35351_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2355),
    .D(_01943_),
    .Q_N(_15199_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][4] ));
 sg13g2_dfrbp_1 _35352_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2354),
    .D(_01944_),
    .Q_N(_15198_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][5] ));
 sg13g2_dfrbp_1 _35353_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2353),
    .D(_01945_),
    .Q_N(_15197_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][6] ));
 sg13g2_dfrbp_1 _35354_ (.CLK(clknet_leaf_304_clk),
    .RESET_B(net2352),
    .D(_01946_),
    .Q_N(_15196_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][7] ));
 sg13g2_dfrbp_1 _35355_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2351),
    .D(_01947_),
    .Q_N(_15195_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][8] ));
 sg13g2_dfrbp_1 _35356_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2350),
    .D(_01948_),
    .Q_N(_15194_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][9] ));
 sg13g2_dfrbp_1 _35357_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2349),
    .D(_01949_),
    .Q_N(_15193_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][10] ));
 sg13g2_dfrbp_1 _35358_ (.CLK(clknet_leaf_313_clk),
    .RESET_B(net2348),
    .D(_01950_),
    .Q_N(_15192_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][11] ));
 sg13g2_dfrbp_1 _35359_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2347),
    .D(_01951_),
    .Q_N(_15191_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][12] ));
 sg13g2_dfrbp_1 _35360_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2346),
    .D(_01952_),
    .Q_N(_15190_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][13] ));
 sg13g2_dfrbp_1 _35361_ (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2345),
    .D(_01953_),
    .Q_N(_15189_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][14] ));
 sg13g2_dfrbp_1 _35362_ (.CLK(clknet_leaf_307_clk),
    .RESET_B(net2344),
    .D(_01954_),
    .Q_N(_15188_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][15] ));
 sg13g2_dfrbp_1 _35363_ (.CLK(clknet_leaf_320_clk),
    .RESET_B(net2343),
    .D(_01955_),
    .Q_N(_15187_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][16] ));
 sg13g2_dfrbp_1 _35364_ (.CLK(clknet_leaf_312_clk),
    .RESET_B(net2342),
    .D(_01956_),
    .Q_N(_15186_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][17] ));
 sg13g2_dfrbp_1 _35365_ (.CLK(clknet_leaf_302_clk),
    .RESET_B(net2341),
    .D(_01957_),
    .Q_N(_15185_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][18] ));
 sg13g2_dfrbp_1 _35366_ (.CLK(clknet_leaf_308_clk),
    .RESET_B(net2340),
    .D(_01958_),
    .Q_N(_15184_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][19] ));
 sg13g2_dfrbp_1 _35367_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2332),
    .D(_01959_),
    .Q_N(_15183_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][20] ));
 sg13g2_dfrbp_1 _35368_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2331),
    .D(_01960_),
    .Q_N(_15182_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][21] ));
 sg13g2_dfrbp_1 _35369_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2330),
    .D(_01961_),
    .Q_N(_15181_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][22] ));
 sg13g2_dfrbp_1 _35370_ (.CLK(clknet_leaf_315_clk),
    .RESET_B(net2329),
    .D(_01962_),
    .Q_N(_15180_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][23] ));
 sg13g2_dfrbp_1 _35371_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2328),
    .D(_01963_),
    .Q_N(_15179_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][24] ));
 sg13g2_dfrbp_1 _35372_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2327),
    .D(_01964_),
    .Q_N(_15178_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][25] ));
 sg13g2_dfrbp_1 _35373_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2326),
    .D(_01965_),
    .Q_N(_15177_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][26] ));
 sg13g2_dfrbp_1 _35374_ (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2325),
    .D(_01966_),
    .Q_N(_15176_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][27] ));
 sg13g2_dfrbp_1 _35375_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2324),
    .D(_01967_),
    .Q_N(_15175_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][28] ));
 sg13g2_dfrbp_1 _35376_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2323),
    .D(_01968_),
    .Q_N(_15174_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][29] ));
 sg13g2_dfrbp_1 _35377_ (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2322),
    .D(_01969_),
    .Q_N(_15173_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][30] ));
 sg13g2_dfrbp_1 _35378_ (.CLK(clknet_leaf_307_clk),
    .RESET_B(net2321),
    .D(_01970_),
    .Q_N(_15172_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][31] ));
 sg13g2_dfrbp_1 _35379_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net2319),
    .D(net3868),
    .Q_N(_00109_),
    .Q(\soc_I.spi0_I.rx_data[0] ));
 sg13g2_dfrbp_1 _35380_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net2315),
    .D(net3720),
    .Q_N(_15171_),
    .Q(\soc_I.spi0_I.rx_data[1] ));
 sg13g2_dfrbp_1 _35381_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net2311),
    .D(net3948),
    .Q_N(_15170_),
    .Q(\soc_I.spi0_I.rx_data[2] ));
 sg13g2_dfrbp_1 _35382_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net2307),
    .D(net4317),
    .Q_N(_15169_),
    .Q(\soc_I.spi0_I.rx_data[3] ));
 sg13g2_dfrbp_1 _35383_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net2303),
    .D(net4009),
    .Q_N(_15168_),
    .Q(\soc_I.spi0_I.rx_data[4] ));
 sg13g2_dfrbp_1 _35384_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net2299),
    .D(net4103),
    .Q_N(_15167_),
    .Q(\soc_I.spi0_I.rx_data[5] ));
 sg13g2_dfrbp_1 _35385_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net2295),
    .D(net4628),
    .Q_N(_15166_),
    .Q(\soc_I.spi0_I.rx_data[6] ));
 sg13g2_dfrbp_1 _35386_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net2291),
    .D(net3706),
    .Q_N(_15165_),
    .Q(\soc_I.spi0_I.rx_data[7] ));
 sg13g2_dfrbp_1 _35387_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net2287),
    .D(net5535),
    .Q_N(_15164_),
    .Q(uio_oe[1]));
 sg13g2_dfrbp_1 _35388_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net2283),
    .D(net5382),
    .Q_N(_15163_),
    .Q(uio_oe[5]));
 sg13g2_dfrbp_1 _35389_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net2279),
    .D(net5395),
    .Q_N(_15162_),
    .Q(uio_out[0]));
 sg13g2_dfrbp_1 _35390_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net2275),
    .D(net5514),
    .Q_N(_15161_),
    .Q(uio_out[6]));
 sg13g2_dfrbp_1 _35391_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net2135),
    .D(_01983_),
    .Q_N(_15160_),
    .Q(uio_out[7]));
 sg13g2_dfrbp_1 _35392_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net2131),
    .D(net3053),
    .Q_N(_00011_),
    .Q(sclk));
 sg13g2_dfrbp_1 _35393_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1999),
    .D(_01985_),
    .Q_N(_15159_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[0] ));
 sg13g2_dfrbp_1 _35394_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1997),
    .D(_01986_),
    .Q_N(_15158_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[1] ));
 sg13g2_dfrbp_1 _35395_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1995),
    .D(_01987_),
    .Q_N(_15157_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[2] ));
 sg13g2_dfrbp_1 _35396_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1993),
    .D(_01988_),
    .Q_N(_15156_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[3] ));
 sg13g2_dfrbp_1 _35397_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1991),
    .D(_01989_),
    .Q_N(_15155_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[4] ));
 sg13g2_dfrbp_1 _35398_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1989),
    .D(_01990_),
    .Q_N(_15154_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[5] ));
 sg13g2_dfrbp_1 _35399_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1987),
    .D(_01991_),
    .Q_N(_15153_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[6] ));
 sg13g2_dfrbp_1 _35400_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1985),
    .D(_01992_),
    .Q_N(_15152_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[7] ));
 sg13g2_dfrbp_1 _35401_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1983),
    .D(_01993_),
    .Q_N(_15151_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[8] ));
 sg13g2_dfrbp_1 _35402_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1981),
    .D(_01994_),
    .Q_N(_15150_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[9] ));
 sg13g2_dfrbp_1 _35403_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1979),
    .D(_01995_),
    .Q_N(_15149_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[10] ));
 sg13g2_dfrbp_1 _35404_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1977),
    .D(_01996_),
    .Q_N(_15148_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[11] ));
 sg13g2_dfrbp_1 _35405_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1975),
    .D(_01997_),
    .Q_N(_15147_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[12] ));
 sg13g2_dfrbp_1 _35406_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1973),
    .D(_01998_),
    .Q_N(_15146_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[13] ));
 sg13g2_dfrbp_1 _35407_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1971),
    .D(_01999_),
    .Q_N(_15145_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[14] ));
 sg13g2_dfrbp_1 _35408_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1969),
    .D(_02000_),
    .Q_N(_15144_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[15] ));
 sg13g2_dfrbp_1 _35409_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1967),
    .D(_02001_),
    .Q_N(_15143_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[16] ));
 sg13g2_dfrbp_1 _35410_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1965),
    .D(_02002_),
    .Q_N(_15142_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[17] ));
 sg13g2_dfrbp_1 _35411_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1963),
    .D(_02003_),
    .Q_N(_15141_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[18] ));
 sg13g2_dfrbp_1 _35412_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1961),
    .D(_02004_),
    .Q_N(_15140_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[19] ));
 sg13g2_dfrbp_1 _35413_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1959),
    .D(_02005_),
    .Q_N(_15139_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[20] ));
 sg13g2_dfrbp_1 _35414_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1957),
    .D(_02006_),
    .Q_N(_15138_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[21] ));
 sg13g2_dfrbp_1 _35415_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1955),
    .D(_02007_),
    .Q_N(_15137_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[22] ));
 sg13g2_dfrbp_1 _35416_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1953),
    .D(_02008_),
    .Q_N(_15136_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[23] ));
 sg13g2_dfrbp_1 _35417_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1951),
    .D(_02009_),
    .Q_N(_15135_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[24] ));
 sg13g2_dfrbp_1 _35418_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1949),
    .D(_02010_),
    .Q_N(_15134_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[25] ));
 sg13g2_dfrbp_1 _35419_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1947),
    .D(_02011_),
    .Q_N(_15133_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[26] ));
 sg13g2_dfrbp_1 _35420_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1945),
    .D(_02012_),
    .Q_N(_15132_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[27] ));
 sg13g2_dfrbp_1 _35421_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1943),
    .D(_02013_),
    .Q_N(_15131_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[28] ));
 sg13g2_dfrbp_1 _35422_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1941),
    .D(_02014_),
    .Q_N(_15130_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[29] ));
 sg13g2_dfrbp_1 _35423_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1939),
    .D(_02015_),
    .Q_N(_15129_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[30] ));
 sg13g2_dfrbp_1 _35424_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1793),
    .D(_02016_),
    .Q_N(_15128_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[31] ));
 sg13g2_dfrbp_1 _35425_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1791),
    .D(_02017_),
    .Q_N(_00244_),
    .Q(\soc_I.qqspi_I.ready ));
 sg13g2_dfrbp_1 _35426_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1723),
    .D(_02018_),
    .Q_N(_15127_),
    .Q(sio0_si_mosi_o));
 sg13g2_dfrbp_1 _35427_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1719),
    .D(_02019_),
    .Q_N(_15126_),
    .Q(sio1_so_miso_o));
 sg13g2_dfrbp_1 _35428_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1715),
    .D(_02020_),
    .Q_N(_15125_),
    .Q(sio2_o));
 sg13g2_dfrbp_1 _35429_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1711),
    .D(_02021_),
    .Q_N(_15124_),
    .Q(sio3_o));
 sg13g2_dfrbp_1 _35430_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1707),
    .D(_02022_),
    .Q_N(_15123_),
    .Q(\soc_I.qqspi_I.spi_buf[24] ));
 sg13g2_dfrbp_1 _35431_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1703),
    .D(_02023_),
    .Q_N(_15122_),
    .Q(\soc_I.qqspi_I.spi_buf[25] ));
 sg13g2_dfrbp_1 _35432_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1699),
    .D(net5418),
    .Q_N(_15121_),
    .Q(\soc_I.qqspi_I.spi_buf[26] ));
 sg13g2_dfrbp_1 _35433_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1695),
    .D(_02025_),
    .Q_N(_15120_),
    .Q(\soc_I.qqspi_I.spi_buf[27] ));
 sg13g2_dfrbp_1 _35434_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1691),
    .D(net5531),
    .Q_N(_15119_),
    .Q(\soc_I.qqspi_I.spi_buf[28] ));
 sg13g2_dfrbp_1 _35435_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1687),
    .D(_02027_),
    .Q_N(_15118_),
    .Q(\soc_I.qqspi_I.spi_buf[29] ));
 sg13g2_dfrbp_1 _35436_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1683),
    .D(_02028_),
    .Q_N(_15117_),
    .Q(\soc_I.qqspi_I.spi_buf[30] ));
 sg13g2_dfrbp_1 _35437_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1679),
    .D(_02029_),
    .Q_N(_15116_),
    .Q(\soc_I.qqspi_I.spi_buf[31] ));
 sg13g2_dfrbp_1 _35438_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1675),
    .D(_02030_),
    .Q_N(_00241_),
    .Q(\soc_I.qqspi_I.is_quad ));
 sg13g2_dfrbp_1 _35439_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1671),
    .D(_02031_),
    .Q_N(_15115_),
    .Q(\soc_I.div_ready ));
 sg13g2_dfrbp_1 _35440_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1669),
    .D(_02032_),
    .Q_N(_15114_),
    .Q(\soc_I.spi_div_ready ));
 sg13g2_dfrbp_1 _35441_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1667),
    .D(_02033_),
    .Q_N(_00106_),
    .Q(\soc_I.div_reg[0] ));
 sg13g2_dfrbp_1 _35442_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1663),
    .D(_02034_),
    .Q_N(_00113_),
    .Q(\soc_I.div_reg[1] ));
 sg13g2_dfrbp_1 _35443_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1659),
    .D(_02035_),
    .Q_N(_00118_),
    .Q(\soc_I.div_reg[2] ));
 sg13g2_dfrbp_1 _35444_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1655),
    .D(_02036_),
    .Q_N(_00123_),
    .Q(\soc_I.div_reg[3] ));
 sg13g2_dfrbp_1 _35445_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1651),
    .D(_02037_),
    .Q_N(_00128_),
    .Q(\soc_I.div_reg[4] ));
 sg13g2_dfrbp_1 _35446_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1647),
    .D(_02038_),
    .Q_N(_00133_),
    .Q(\soc_I.div_reg[5] ));
 sg13g2_dfrbp_1 _35447_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1643),
    .D(_02039_),
    .Q_N(_00138_),
    .Q(\soc_I.div_reg[6] ));
 sg13g2_dfrbp_1 _35448_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1639),
    .D(_02040_),
    .Q_N(_00143_),
    .Q(\soc_I.div_reg[7] ));
 sg13g2_dfrbp_1 _35449_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1635),
    .D(_02041_),
    .Q_N(_00074_),
    .Q(\soc_I.div_reg[8] ));
 sg13g2_dfrbp_1 _35450_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1631),
    .D(_02042_),
    .Q_N(_00078_),
    .Q(\soc_I.div_reg[9] ));
 sg13g2_dfrbp_1 _35451_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1627),
    .D(_02043_),
    .Q_N(_00082_),
    .Q(\soc_I.div_reg[10] ));
 sg13g2_dfrbp_1 _35452_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1623),
    .D(_02044_),
    .Q_N(_00086_),
    .Q(\soc_I.div_reg[11] ));
 sg13g2_dfrbp_1 _35453_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1619),
    .D(_02045_),
    .Q_N(_00090_),
    .Q(\soc_I.div_reg[12] ));
 sg13g2_dfrbp_1 _35454_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1615),
    .D(_02046_),
    .Q_N(_00094_),
    .Q(\soc_I.div_reg[13] ));
 sg13g2_dfrbp_1 _35455_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1611),
    .D(_02047_),
    .Q_N(_00098_),
    .Q(\soc_I.div_reg[14] ));
 sg13g2_dfrbp_1 _35456_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1607),
    .D(_02048_),
    .Q_N(_00102_),
    .Q(\soc_I.div_reg[15] ));
 sg13g2_dfrbp_1 _35457_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1603),
    .D(_02049_),
    .Q_N(_00012_),
    .Q(\soc_I.clint_I.div[0] ));
 sg13g2_dfrbp_1 _35458_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1599),
    .D(_02050_),
    .Q_N(_00019_),
    .Q(\soc_I.clint_I.div[1] ));
 sg13g2_dfrbp_1 _35459_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1595),
    .D(_02051_),
    .Q_N(_00027_),
    .Q(\soc_I.clint_I.div[2] ));
 sg13g2_dfrbp_1 _35460_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1591),
    .D(_02052_),
    .Q_N(_00035_),
    .Q(\soc_I.clint_I.div[3] ));
 sg13g2_dfrbp_1 _35461_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1587),
    .D(_02053_),
    .Q_N(_00246_),
    .Q(\soc_I.clint_I.div[4] ));
 sg13g2_dfrbp_1 _35462_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1583),
    .D(_02054_),
    .Q_N(_00049_),
    .Q(\soc_I.clint_I.div[5] ));
 sg13g2_dfrbp_1 _35463_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1579),
    .D(_02055_),
    .Q_N(_00057_),
    .Q(\soc_I.clint_I.div[6] ));
 sg13g2_dfrbp_1 _35464_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1575),
    .D(_02056_),
    .Q_N(_00065_),
    .Q(\soc_I.clint_I.div[7] ));
 sg13g2_dfrbp_1 _35465_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1571),
    .D(_02057_),
    .Q_N(_00247_),
    .Q(\soc_I.clint_I.div[8] ));
 sg13g2_dfrbp_1 _35466_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1567),
    .D(_02058_),
    .Q_N(_00023_),
    .Q(\soc_I.clint_I.div[9] ));
 sg13g2_dfrbp_1 _35467_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1563),
    .D(_02059_),
    .Q_N(_00031_),
    .Q(\soc_I.clint_I.div[10] ));
 sg13g2_dfrbp_1 _35468_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1559),
    .D(_02060_),
    .Q_N(_00039_),
    .Q(\soc_I.clint_I.div[11] ));
 sg13g2_dfrbp_1 _35469_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1555),
    .D(_02061_),
    .Q_N(_00248_),
    .Q(\soc_I.clint_I.div[12] ));
 sg13g2_dfrbp_1 _35470_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1551),
    .D(_02062_),
    .Q_N(_00053_),
    .Q(\soc_I.clint_I.div[13] ));
 sg13g2_dfrbp_1 _35471_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1547),
    .D(_02063_),
    .Q_N(_00061_),
    .Q(\soc_I.clint_I.div[14] ));
 sg13g2_dfrbp_1 _35472_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1543),
    .D(_02064_),
    .Q_N(_00069_),
    .Q(\soc_I.clint_I.div[15] ));
 sg13g2_dfrbp_1 _35473_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1539),
    .D(_02065_),
    .Q_N(_15113_),
    .Q(\soc_I.uart_tx_ready ));
 sg13g2_dfrbp_1 _35474_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1537),
    .D(_02066_),
    .Q_N(_00107_),
    .Q(\soc_I.spi0_I.div[0] ));
 sg13g2_dfrbp_1 _35475_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1533),
    .D(_02067_),
    .Q_N(_00114_),
    .Q(\soc_I.spi0_I.div[1] ));
 sg13g2_dfrbp_1 _35476_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1529),
    .D(_02068_),
    .Q_N(_00119_),
    .Q(\soc_I.spi0_I.div[2] ));
 sg13g2_dfrbp_1 _35477_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1525),
    .D(_02069_),
    .Q_N(_00124_),
    .Q(\soc_I.spi0_I.div[3] ));
 sg13g2_dfrbp_1 _35478_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1521),
    .D(_02070_),
    .Q_N(_00129_),
    .Q(\soc_I.spi0_I.div[4] ));
 sg13g2_dfrbp_1 _35479_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1517),
    .D(_02071_),
    .Q_N(_00134_),
    .Q(\soc_I.spi0_I.div[5] ));
 sg13g2_dfrbp_1 _35480_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1513),
    .D(_02072_),
    .Q_N(_00139_),
    .Q(\soc_I.spi0_I.div[6] ));
 sg13g2_dfrbp_1 _35481_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1509),
    .D(_02073_),
    .Q_N(_00144_),
    .Q(\soc_I.spi0_I.div[7] ));
 sg13g2_dfrbp_1 _35482_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1505),
    .D(_02074_),
    .Q_N(_00287_),
    .Q(\soc_I.spi0_I.div[8] ));
 sg13g2_dfrbp_1 _35483_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1501),
    .D(_02075_),
    .Q_N(_15112_),
    .Q(\soc_I.spi0_I.div[9] ));
 sg13g2_dfrbp_1 _35484_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1497),
    .D(_02076_),
    .Q_N(_15111_),
    .Q(\soc_I.spi0_I.div[10] ));
 sg13g2_dfrbp_1 _35485_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1493),
    .D(_02077_),
    .Q_N(_15110_),
    .Q(\soc_I.spi0_I.div[11] ));
 sg13g2_dfrbp_1 _35486_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1489),
    .D(_02078_),
    .Q_N(_00288_),
    .Q(\soc_I.spi0_I.div[12] ));
 sg13g2_dfrbp_1 _35487_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1485),
    .D(_02079_),
    .Q_N(_15109_),
    .Q(\soc_I.spi0_I.div[13] ));
 sg13g2_dfrbp_1 _35488_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1481),
    .D(_02080_),
    .Q_N(_15108_),
    .Q(\soc_I.spi0_I.div[14] ));
 sg13g2_dfrbp_1 _35489_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1477),
    .D(_02081_),
    .Q_N(_15107_),
    .Q(\soc_I.spi0_I.div[15] ));
 sg13g2_dfrbp_1 _35490_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1473),
    .D(_02082_),
    .Q_N(_15106_),
    .Q(\soc_I.spi_div_reg[16] ));
 sg13g2_dfrbp_1 _35491_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1469),
    .D(_02083_),
    .Q_N(_15105_),
    .Q(\soc_I.spi_div_reg[17] ));
 sg13g2_dfrbp_1 _35492_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1465),
    .D(_02084_),
    .Q_N(_15104_),
    .Q(\soc_I.spi_div_reg[18] ));
 sg13g2_dfrbp_1 _35493_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1461),
    .D(_02085_),
    .Q_N(_15103_),
    .Q(\soc_I.spi_div_reg[19] ));
 sg13g2_dfrbp_1 _35494_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1457),
    .D(_02086_),
    .Q_N(_15102_),
    .Q(\soc_I.spi_div_reg[20] ));
 sg13g2_dfrbp_1 _35495_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1453),
    .D(_02087_),
    .Q_N(_15101_),
    .Q(\soc_I.spi_div_reg[21] ));
 sg13g2_dfrbp_1 _35496_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1449),
    .D(_02088_),
    .Q_N(_15100_),
    .Q(\soc_I.spi_div_reg[22] ));
 sg13g2_dfrbp_1 _35497_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1445),
    .D(_02089_),
    .Q_N(_15099_),
    .Q(\soc_I.spi_div_reg[23] ));
 sg13g2_dfrbp_1 _35498_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1441),
    .D(_02090_),
    .Q_N(_15098_),
    .Q(\soc_I.spi_div_reg[24] ));
 sg13g2_dfrbp_1 _35499_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1437),
    .D(_02091_),
    .Q_N(_15097_),
    .Q(\soc_I.spi_div_reg[25] ));
 sg13g2_dfrbp_1 _35500_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1433),
    .D(_02092_),
    .Q_N(_15096_),
    .Q(\soc_I.spi_div_reg[26] ));
 sg13g2_dfrbp_1 _35501_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1429),
    .D(_02093_),
    .Q_N(_15095_),
    .Q(\soc_I.spi_div_reg[27] ));
 sg13g2_dfrbp_1 _35502_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1425),
    .D(_02094_),
    .Q_N(_15094_),
    .Q(\soc_I.spi_div_reg[28] ));
 sg13g2_dfrbp_1 _35503_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1421),
    .D(_02095_),
    .Q_N(_15093_),
    .Q(\soc_I.spi_div_reg[29] ));
 sg13g2_dfrbp_1 _35504_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1417),
    .D(_02096_),
    .Q_N(_15092_),
    .Q(\soc_I.spi_div_reg[30] ));
 sg13g2_dfrbp_1 _35505_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1413),
    .D(_02097_),
    .Q_N(_00070_),
    .Q(\soc_I.spi_div_reg[31] ));
 sg13g2_dfrbp_1 _35506_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1409),
    .D(_02098_),
    .Q_N(_00250_),
    .Q(\soc_I.uart_lsr_rdy ));
 sg13g2_dfrbp_1 _35507_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1407),
    .D(_02099_),
    .Q_N(_00292_),
    .Q(\soc_I.rx_uart_i.data_rd ));
 sg13g2_dfrbp_1 _35508_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1304),
    .D(net2622),
    .Q_N(_15091_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[8][0] ));
 sg13g2_dfrbp_1 _35509_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1302),
    .D(net4147),
    .Q_N(_15090_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[8][1] ));
 sg13g2_dfrbp_1 _35510_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1300),
    .D(_02102_),
    .Q_N(_15089_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[8][2] ));
 sg13g2_dfrbp_1 _35511_ (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1298),
    .D(net3692),
    .Q_N(_15088_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[8][3] ));
 sg13g2_dfrbp_1 _35512_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1296),
    .D(net4210),
    .Q_N(_15087_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[8][4] ));
 sg13g2_dfrbp_1 _35513_ (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1294),
    .D(_02105_),
    .Q_N(_15086_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[8][5] ));
 sg13g2_dfrbp_1 _35514_ (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1292),
    .D(net3621),
    .Q_N(_15085_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[8][6] ));
 sg13g2_dfrbp_1 _35515_ (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1290),
    .D(net3533),
    .Q_N(_15084_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[8][7] ));
 sg13g2_dfrbp_1 _35516_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1288),
    .D(_02108_),
    .Q_N(_15083_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[31] ));
 sg13g2_dfrbp_1 _35517_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1284),
    .D(_02109_),
    .Q_N(_15082_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[0] ));
 sg13g2_dfrbp_1 _35518_ (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1280),
    .D(_02110_),
    .Q_N(_15081_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[1] ));
 sg13g2_dfrbp_1 _35519_ (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1276),
    .D(_02111_),
    .Q_N(_15080_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[2] ));
 sg13g2_dfrbp_1 _35520_ (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1272),
    .D(_02112_),
    .Q_N(_15079_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[4] ));
 sg13g2_dfrbp_1 _35521_ (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1268),
    .D(_02113_),
    .Q_N(_15078_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[5] ));
 sg13g2_dfrbp_1 _35522_ (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1264),
    .D(_02114_),
    .Q_N(_15077_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[6] ));
 sg13g2_dfrbp_1 _35523_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1260),
    .D(_02115_),
    .Q_N(_15076_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[8] ));
 sg13g2_dfrbp_1 _35524_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1256),
    .D(_02116_),
    .Q_N(_15075_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[9] ));
 sg13g2_dfrbp_1 _35525_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1252),
    .D(_02117_),
    .Q_N(_15074_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[10] ));
 sg13g2_dfrbp_1 _35526_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1248),
    .D(_02118_),
    .Q_N(_15073_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[13] ));
 sg13g2_dfrbp_1 _35527_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1244),
    .D(_02119_),
    .Q_N(_15072_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[14] ));
 sg13g2_dfrbp_1 _35528_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1240),
    .D(_02120_),
    .Q_N(_15071_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[15] ));
 sg13g2_dfrbp_1 _35529_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1236),
    .D(_02121_),
    .Q_N(_15070_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[16] ));
 sg13g2_dfrbp_1 _35530_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1232),
    .D(_02122_),
    .Q_N(_15069_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[17] ));
 sg13g2_dfrbp_1 _35531_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1228),
    .D(_02123_),
    .Q_N(_15068_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[18] ));
 sg13g2_dfrbp_1 _35532_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1224),
    .D(_02124_),
    .Q_N(_15067_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[19] ));
 sg13g2_dfrbp_1 _35533_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1220),
    .D(_02125_),
    .Q_N(_15066_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[20] ));
 sg13g2_dfrbp_1 _35534_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1216),
    .D(_02126_),
    .Q_N(_15065_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[21] ));
 sg13g2_dfrbp_1 _35535_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1212),
    .D(_02127_),
    .Q_N(_15064_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[22] ));
 sg13g2_dfrbp_1 _35536_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1208),
    .D(_02128_),
    .Q_N(_15063_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[23] ));
 sg13g2_dfrbp_1 _35537_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1204),
    .D(_02129_),
    .Q_N(_15062_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[24] ));
 sg13g2_dfrbp_1 _35538_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1200),
    .D(_02130_),
    .Q_N(_15061_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[25] ));
 sg13g2_dfrbp_1 _35539_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1196),
    .D(_02131_),
    .Q_N(_15060_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[26] ));
 sg13g2_dfrbp_1 _35540_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1192),
    .D(_02132_),
    .Q_N(_15059_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[27] ));
 sg13g2_dfrbp_1 _35541_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1188),
    .D(_02133_),
    .Q_N(_15058_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[28] ));
 sg13g2_dfrbp_1 _35542_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1184),
    .D(_02134_),
    .Q_N(_15057_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[29] ));
 sg13g2_dfrbp_1 _35543_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1180),
    .D(_02135_),
    .Q_N(_15056_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[30] ));
 sg13g2_dfrbp_1 _35544_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1176),
    .D(_02136_),
    .Q_N(_15055_),
    .Q(\soc_I.tx_uart_i.wait_states[0] ));
 sg13g2_dfrbp_1 _35545_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1172),
    .D(_02137_),
    .Q_N(_15054_),
    .Q(\soc_I.tx_uart_i.return_state[1] ));
 sg13g2_dfrbp_1 _35546_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1168),
    .D(net3928),
    .Q_N(_15053_),
    .Q(\soc_I.tx_uart_i.return_state[0] ));
 sg13g2_dfrbp_1 _35547_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1100),
    .D(net3010),
    .Q_N(_15052_),
    .Q(\soc_I.rx_uart_i.return_state[1] ));
 sg13g2_dfrbp_1 _35548_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1096),
    .D(_02140_),
    .Q_N(_15051_),
    .Q(\soc_I.rx_uart_i.return_state[0] ));
 sg13g2_dfrbp_1 _35549_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1092),
    .D(net2602),
    .Q_N(_00184_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_state[2] ));
 sg13g2_dfrbp_1 _35550_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1090),
    .D(net2617),
    .Q_N(_15050_),
    .Q(\soc_I.kianv_I.datapath_unit_I.div_I.div_state[1] ));
 sg13g2_dfrbp_1 _35551_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1088),
    .D(_02143_),
    .Q_N(_15049_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.state[2] ));
 sg13g2_dfrbp_1 _35552_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1086),
    .D(_02144_),
    .Q_N(_15048_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.state[1] ));
 sg13g2_dfrbp_1 _35553_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1084),
    .D(_02145_),
    .Q_N(_15047_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[63] ));
 sg13g2_dfrbp_1 _35554_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1080),
    .D(net4616),
    .Q_N(_15046_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[62] ));
 sg13g2_dfrbp_1 _35555_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1076),
    .D(_02147_),
    .Q_N(_00282_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[61] ));
 sg13g2_dfrbp_1 _35556_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1072),
    .D(net4950),
    .Q_N(_00281_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[60] ));
 sg13g2_dfrbp_1 _35557_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1068),
    .D(net5103),
    .Q_N(_00280_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[59] ));
 sg13g2_dfrbp_1 _35558_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1064),
    .D(_02150_),
    .Q_N(_00279_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[58] ));
 sg13g2_dfrbp_1 _35559_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1060),
    .D(_02151_),
    .Q_N(_00278_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[57] ));
 sg13g2_dfrbp_1 _35560_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1056),
    .D(net4532),
    .Q_N(_00277_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[56] ));
 sg13g2_dfrbp_1 _35561_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1052),
    .D(_02153_),
    .Q_N(_00276_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[55] ));
 sg13g2_dfrbp_1 _35562_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1048),
    .D(_02154_),
    .Q_N(_00275_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[54] ));
 sg13g2_dfrbp_1 _35563_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1044),
    .D(_02155_),
    .Q_N(_00274_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[53] ));
 sg13g2_dfrbp_1 _35564_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1040),
    .D(_02156_),
    .Q_N(_00273_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[52] ));
 sg13g2_dfrbp_1 _35565_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1036),
    .D(_02157_),
    .Q_N(_15045_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[51] ));
 sg13g2_dfrbp_1 _35566_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1032),
    .D(net4835),
    .Q_N(_00272_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[50] ));
 sg13g2_dfrbp_1 _35567_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1028),
    .D(net4368),
    .Q_N(_00271_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[49] ));
 sg13g2_dfrbp_1 _35568_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1024),
    .D(_02160_),
    .Q_N(_00270_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[48] ));
 sg13g2_dfrbp_1 _35569_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1020),
    .D(_02161_),
    .Q_N(_15044_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[47] ));
 sg13g2_dfrbp_1 _35570_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1016),
    .D(_02162_),
    .Q_N(_15043_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[46] ));
 sg13g2_dfrbp_1 _35571_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1012),
    .D(_02163_),
    .Q_N(_15042_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[45] ));
 sg13g2_dfrbp_1 _35572_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1008),
    .D(_02164_),
    .Q_N(_15041_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[44] ));
 sg13g2_dfrbp_1 _35573_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1004),
    .D(_02165_),
    .Q_N(_15040_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[43] ));
 sg13g2_dfrbp_1 _35574_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1000),
    .D(_02166_),
    .Q_N(_15039_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[42] ));
 sg13g2_dfrbp_1 _35575_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net996),
    .D(_02167_),
    .Q_N(_15038_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[41] ));
 sg13g2_dfrbp_1 _35576_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net992),
    .D(_02168_),
    .Q_N(_15037_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[40] ));
 sg13g2_dfrbp_1 _35577_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net988),
    .D(_02169_),
    .Q_N(_15036_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[39] ));
 sg13g2_dfrbp_1 _35578_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net984),
    .D(net5115),
    .Q_N(_15035_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[38] ));
 sg13g2_dfrbp_1 _35579_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net980),
    .D(_02171_),
    .Q_N(_15034_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[37] ));
 sg13g2_dfrbp_1 _35580_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net976),
    .D(_02172_),
    .Q_N(_15033_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[36] ));
 sg13g2_dfrbp_1 _35581_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net972),
    .D(_02173_),
    .Q_N(_15032_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[35] ));
 sg13g2_dfrbp_1 _35582_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net968),
    .D(_02174_),
    .Q_N(_15031_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[34] ));
 sg13g2_dfrbp_1 _35583_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net964),
    .D(_02175_),
    .Q_N(_15030_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[33] ));
 sg13g2_dfrbp_1 _35584_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net960),
    .D(net5432),
    .Q_N(_15029_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[32] ));
 sg13g2_dfrbp_1 _35585_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net956),
    .D(net5336),
    .Q_N(_15028_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[31] ));
 sg13g2_dfrbp_1 _35586_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net952),
    .D(_02178_),
    .Q_N(_15027_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[30] ));
 sg13g2_dfrbp_1 _35587_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net948),
    .D(_02179_),
    .Q_N(_15026_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[29] ));
 sg13g2_dfrbp_1 _35588_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net944),
    .D(_02180_),
    .Q_N(_15025_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[28] ));
 sg13g2_dfrbp_1 _35589_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net940),
    .D(_02181_),
    .Q_N(_15024_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[27] ));
 sg13g2_dfrbp_1 _35590_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net936),
    .D(_02182_),
    .Q_N(_15023_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[26] ));
 sg13g2_dfrbp_1 _35591_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net932),
    .D(net5193),
    .Q_N(_15022_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[25] ));
 sg13g2_dfrbp_1 _35592_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net928),
    .D(_02184_),
    .Q_N(_15021_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[24] ));
 sg13g2_dfrbp_1 _35593_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net924),
    .D(_02185_),
    .Q_N(_15020_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[23] ));
 sg13g2_dfrbp_1 _35594_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net920),
    .D(_02186_),
    .Q_N(_15019_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[22] ));
 sg13g2_dfrbp_1 _35595_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net916),
    .D(_02187_),
    .Q_N(_15018_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[21] ));
 sg13g2_dfrbp_1 _35596_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net912),
    .D(_02188_),
    .Q_N(_15017_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[20] ));
 sg13g2_dfrbp_1 _35597_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net908),
    .D(_02189_),
    .Q_N(_15016_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[19] ));
 sg13g2_dfrbp_1 _35598_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net904),
    .D(_02190_),
    .Q_N(_15015_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[18] ));
 sg13g2_dfrbp_1 _35599_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net900),
    .D(_02191_),
    .Q_N(_15014_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[17] ));
 sg13g2_dfrbp_1 _35600_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net896),
    .D(_02192_),
    .Q_N(_15013_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[16] ));
 sg13g2_dfrbp_1 _35601_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net892),
    .D(_02193_),
    .Q_N(_15012_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[15] ));
 sg13g2_dfrbp_1 _35602_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net888),
    .D(_02194_),
    .Q_N(_00269_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[14] ));
 sg13g2_dfrbp_1 _35603_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net884),
    .D(_02195_),
    .Q_N(_00268_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[13] ));
 sg13g2_dfrbp_1 _35604_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net880),
    .D(_02196_),
    .Q_N(_00267_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[12] ));
 sg13g2_dfrbp_1 _35605_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net876),
    .D(_02197_),
    .Q_N(_15011_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[11] ));
 sg13g2_dfrbp_1 _35606_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net872),
    .D(_02198_),
    .Q_N(_00266_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[10] ));
 sg13g2_dfrbp_1 _35607_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net868),
    .D(net5084),
    .Q_N(_00265_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[9] ));
 sg13g2_dfrbp_1 _35608_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net864),
    .D(_02200_),
    .Q_N(_00264_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[8] ));
 sg13g2_dfrbp_1 _35609_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net860),
    .D(_02201_),
    .Q_N(_00263_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[7] ));
 sg13g2_dfrbp_1 _35610_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net856),
    .D(_02202_),
    .Q_N(_00262_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[6] ));
 sg13g2_dfrbp_1 _35611_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net852),
    .D(net3230),
    .Q_N(_00261_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[5] ));
 sg13g2_dfrbp_1 _35612_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net848),
    .D(net5070),
    .Q_N(_00260_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[4] ));
 sg13g2_dfrbp_1 _35613_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net780),
    .D(_02205_),
    .Q_N(_00259_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[3] ));
 sg13g2_dfrbp_1 _35614_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net776),
    .D(net5202),
    .Q_N(_00258_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[2] ));
 sg13g2_dfrbp_1 _35615_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net772),
    .D(_02207_),
    .Q_N(_00257_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[1] ));
 sg13g2_dfrbp_1 _35616_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net735),
    .D(net4492),
    .Q_N(_00253_),
    .Q(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[0] ));
 sg13g2_dfrbp_1 _35617_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net731),
    .D(_02209_),
    .Q_N(_15010_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[5] ));
 sg13g2_dfrbp_1 _35618_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net729),
    .D(_02210_),
    .Q_N(_15009_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[4] ));
 sg13g2_dfrbp_1 _35619_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net727),
    .D(_02211_),
    .Q_N(_15008_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[3] ));
 sg13g2_dfrbp_1 _35620_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net724),
    .D(_02212_),
    .Q_N(_15007_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[2] ));
 sg13g2_dfrbp_1 _35621_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net722),
    .D(_02213_),
    .Q_N(_15006_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[1] ));
 sg13g2_dfrbp_1 _35622_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net720),
    .D(_02214_),
    .Q_N(_15005_),
    .Q(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[0] ));
 sg13g2_dfrbp_1 _35623_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net718),
    .D(_02215_),
    .Q_N(_15004_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][0] ));
 sg13g2_dfrbp_1 _35624_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net716),
    .D(_02216_),
    .Q_N(_15003_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][1] ));
 sg13g2_dfrbp_1 _35625_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net714),
    .D(_02217_),
    .Q_N(_15002_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][2] ));
 sg13g2_dfrbp_1 _35626_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net712),
    .D(_02218_),
    .Q_N(_15001_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][3] ));
 sg13g2_dfrbp_1 _35627_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net710),
    .D(_02219_),
    .Q_N(_15000_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][4] ));
 sg13g2_dfrbp_1 _35628_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net708),
    .D(_02220_),
    .Q_N(_14999_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][5] ));
 sg13g2_dfrbp_1 _35629_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net706),
    .D(_02221_),
    .Q_N(_14998_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][6] ));
 sg13g2_dfrbp_1 _35630_ (.CLK(clknet_leaf_305_clk),
    .RESET_B(net704),
    .D(_02222_),
    .Q_N(_14997_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][7] ));
 sg13g2_dfrbp_1 _35631_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net702),
    .D(_02223_),
    .Q_N(_14996_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][8] ));
 sg13g2_dfrbp_1 _35632_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net700),
    .D(_02224_),
    .Q_N(_14995_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][9] ));
 sg13g2_dfrbp_1 _35633_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net698),
    .D(_02225_),
    .Q_N(_14994_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][10] ));
 sg13g2_dfrbp_1 _35634_ (.CLK(clknet_leaf_315_clk),
    .RESET_B(net696),
    .D(_02226_),
    .Q_N(_14993_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][11] ));
 sg13g2_dfrbp_1 _35635_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net694),
    .D(_02227_),
    .Q_N(_14992_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][12] ));
 sg13g2_dfrbp_1 _35636_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net692),
    .D(_02228_),
    .Q_N(_14991_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][13] ));
 sg13g2_dfrbp_1 _35637_ (.CLK(clknet_leaf_300_clk),
    .RESET_B(net690),
    .D(_02229_),
    .Q_N(_14990_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][14] ));
 sg13g2_dfrbp_1 _35638_ (.CLK(clknet_leaf_310_clk),
    .RESET_B(net688),
    .D(_02230_),
    .Q_N(_14989_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][15] ));
 sg13g2_dfrbp_1 _35639_ (.CLK(clknet_leaf_316_clk),
    .RESET_B(net686),
    .D(_02231_),
    .Q_N(_14988_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][16] ));
 sg13g2_dfrbp_1 _35640_ (.CLK(clknet_leaf_314_clk),
    .RESET_B(net684),
    .D(net3649),
    .Q_N(_14987_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][17] ));
 sg13g2_dfrbp_1 _35641_ (.CLK(clknet_leaf_306_clk),
    .RESET_B(net682),
    .D(_02233_),
    .Q_N(_14986_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][18] ));
 sg13g2_dfrbp_1 _35642_ (.CLK(clknet_leaf_302_clk),
    .RESET_B(net680),
    .D(_02234_),
    .Q_N(_14985_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][19] ));
 sg13g2_dfrbp_1 _35643_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net678),
    .D(_02235_),
    .Q_N(_14984_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][20] ));
 sg13g2_dfrbp_1 _35644_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net676),
    .D(_02236_),
    .Q_N(_14983_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][21] ));
 sg13g2_dfrbp_1 _35645_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net674),
    .D(_02237_),
    .Q_N(_14982_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][22] ));
 sg13g2_dfrbp_1 _35646_ (.CLK(clknet_leaf_284_clk),
    .RESET_B(net672),
    .D(_02238_),
    .Q_N(_14981_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][23] ));
 sg13g2_dfrbp_1 _35647_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net670),
    .D(_02239_),
    .Q_N(_14980_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][24] ));
 sg13g2_dfrbp_1 _35648_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net668),
    .D(_02240_),
    .Q_N(_14979_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][25] ));
 sg13g2_dfrbp_1 _35649_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net666),
    .D(_02241_),
    .Q_N(_14978_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][26] ));
 sg13g2_dfrbp_1 _35650_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net664),
    .D(_02242_),
    .Q_N(_14977_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][27] ));
 sg13g2_dfrbp_1 _35651_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net662),
    .D(_02243_),
    .Q_N(_14976_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][28] ));
 sg13g2_dfrbp_1 _35652_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net660),
    .D(_02244_),
    .Q_N(_14975_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][29] ));
 sg13g2_dfrbp_1 _35653_ (.CLK(clknet_leaf_291_clk),
    .RESET_B(net658),
    .D(_02245_),
    .Q_N(_14974_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][30] ));
 sg13g2_dfrbp_1 _35654_ (.CLK(clknet_leaf_285_clk),
    .RESET_B(net656),
    .D(_02246_),
    .Q_N(_14973_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][31] ));
 sg13g2_dfrbp_1 _35655_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net654),
    .D(_02247_),
    .Q_N(_14972_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][0] ));
 sg13g2_dfrbp_1 _35656_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net652),
    .D(_02248_),
    .Q_N(_14971_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][1] ));
 sg13g2_dfrbp_1 _35657_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net650),
    .D(_02249_),
    .Q_N(_14970_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][2] ));
 sg13g2_dfrbp_1 _35658_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net648),
    .D(_02250_),
    .Q_N(_14969_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][3] ));
 sg13g2_dfrbp_1 _35659_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net646),
    .D(_02251_),
    .Q_N(_14968_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][4] ));
 sg13g2_dfrbp_1 _35660_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net644),
    .D(_02252_),
    .Q_N(_14967_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][5] ));
 sg13g2_dfrbp_1 _35661_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net642),
    .D(_02253_),
    .Q_N(_14966_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][6] ));
 sg13g2_dfrbp_1 _35662_ (.CLK(clknet_leaf_302_clk),
    .RESET_B(net640),
    .D(_02254_),
    .Q_N(_14965_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][7] ));
 sg13g2_dfrbp_1 _35663_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net638),
    .D(_02255_),
    .Q_N(_14964_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][8] ));
 sg13g2_dfrbp_1 _35664_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net636),
    .D(_02256_),
    .Q_N(_14963_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][9] ));
 sg13g2_dfrbp_1 _35665_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net634),
    .D(_02257_),
    .Q_N(_14962_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][10] ));
 sg13g2_dfrbp_1 _35666_ (.CLK(clknet_leaf_315_clk),
    .RESET_B(net632),
    .D(_02258_),
    .Q_N(_14961_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][11] ));
 sg13g2_dfrbp_1 _35667_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net630),
    .D(_02259_),
    .Q_N(_14960_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][12] ));
 sg13g2_dfrbp_1 _35668_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net628),
    .D(_02260_),
    .Q_N(_14959_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][13] ));
 sg13g2_dfrbp_1 _35669_ (.CLK(clknet_leaf_299_clk),
    .RESET_B(net626),
    .D(_02261_),
    .Q_N(_14958_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][14] ));
 sg13g2_dfrbp_1 _35670_ (.CLK(clknet_leaf_310_clk),
    .RESET_B(net624),
    .D(_02262_),
    .Q_N(_14957_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][15] ));
 sg13g2_dfrbp_1 _35671_ (.CLK(clknet_leaf_317_clk),
    .RESET_B(net622),
    .D(_02263_),
    .Q_N(_14956_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][16] ));
 sg13g2_dfrbp_1 _35672_ (.CLK(clknet_leaf_312_clk),
    .RESET_B(net620),
    .D(_02264_),
    .Q_N(_14955_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][17] ));
 sg13g2_dfrbp_1 _35673_ (.CLK(clknet_leaf_304_clk),
    .RESET_B(net618),
    .D(_02265_),
    .Q_N(_14954_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][18] ));
 sg13g2_dfrbp_1 _35674_ (.CLK(clknet_leaf_302_clk),
    .RESET_B(net616),
    .D(_02266_),
    .Q_N(_14953_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][19] ));
 sg13g2_dfrbp_1 _35675_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net614),
    .D(_02267_),
    .Q_N(_14952_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][20] ));
 sg13g2_dfrbp_1 _35676_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net612),
    .D(_02268_),
    .Q_N(_14951_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][21] ));
 sg13g2_dfrbp_1 _35677_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net610),
    .D(_02269_),
    .Q_N(_14950_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][22] ));
 sg13g2_dfrbp_1 _35678_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net608),
    .D(_02270_),
    .Q_N(_14949_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][23] ));
 sg13g2_dfrbp_1 _35679_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net606),
    .D(_02271_),
    .Q_N(_14948_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][24] ));
 sg13g2_dfrbp_1 _35680_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net604),
    .D(_02272_),
    .Q_N(_14947_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][25] ));
 sg13g2_dfrbp_1 _35681_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net602),
    .D(_02273_),
    .Q_N(_14946_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][26] ));
 sg13g2_dfrbp_1 _35682_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net600),
    .D(_02274_),
    .Q_N(_14945_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][27] ));
 sg13g2_dfrbp_1 _35683_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net598),
    .D(_02275_),
    .Q_N(_14944_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][28] ));
 sg13g2_dfrbp_1 _35684_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net596),
    .D(_02276_),
    .Q_N(_14943_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][29] ));
 sg13g2_dfrbp_1 _35685_ (.CLK(clknet_leaf_298_clk),
    .RESET_B(net594),
    .D(_02277_),
    .Q_N(_14942_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][30] ));
 sg13g2_dfrbp_1 _35686_ (.CLK(clknet_leaf_284_clk),
    .RESET_B(net592),
    .D(_02278_),
    .Q_N(_14941_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][31] ));
 sg13g2_dfrbp_1 _35687_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net590),
    .D(_02279_),
    .Q_N(_14940_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[7][0] ));
 sg13g2_dfrbp_1 _35688_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net588),
    .D(_02280_),
    .Q_N(_14939_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[7][1] ));
 sg13g2_dfrbp_1 _35689_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net586),
    .D(_02281_),
    .Q_N(_14938_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[7][2] ));
 sg13g2_dfrbp_1 _35690_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net584),
    .D(net4255),
    .Q_N(_14937_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[7][3] ));
 sg13g2_dfrbp_1 _35691_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net582),
    .D(net4017),
    .Q_N(_14936_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[7][4] ));
 sg13g2_dfrbp_1 _35692_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net580),
    .D(net4038),
    .Q_N(_14935_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[7][5] ));
 sg13g2_dfrbp_1 _35693_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net578),
    .D(_02285_),
    .Q_N(_14934_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[7][6] ));
 sg13g2_dfrbp_1 _35694_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net576),
    .D(net4113),
    .Q_N(_14933_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[7][7] ));
 sg13g2_dfrbp_1 _35695_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net574),
    .D(_02287_),
    .Q_N(_14932_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[6][0] ));
 sg13g2_dfrbp_1 _35696_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net572),
    .D(_02288_),
    .Q_N(_14931_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[6][1] ));
 sg13g2_dfrbp_1 _35697_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net570),
    .D(net3957),
    .Q_N(_14930_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[6][2] ));
 sg13g2_dfrbp_1 _35698_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net568),
    .D(net4054),
    .Q_N(_14929_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[6][3] ));
 sg13g2_dfrbp_1 _35699_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net566),
    .D(net4011),
    .Q_N(_14928_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[6][4] ));
 sg13g2_dfrbp_1 _35700_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net564),
    .D(net4015),
    .Q_N(_14927_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[6][5] ));
 sg13g2_dfrbp_1 _35701_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net562),
    .D(_02293_),
    .Q_N(_14926_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[6][6] ));
 sg13g2_dfrbp_1 _35702_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net560),
    .D(net4319),
    .Q_N(_14925_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[6][7] ));
 sg13g2_dfrbp_1 _35703_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net558),
    .D(_02295_),
    .Q_N(_14924_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[5][0] ));
 sg13g2_dfrbp_1 _35704_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net556),
    .D(_02296_),
    .Q_N(_14923_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[5][1] ));
 sg13g2_dfrbp_1 _35705_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net554),
    .D(_02297_),
    .Q_N(_14922_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[5][2] ));
 sg13g2_dfrbp_1 _35706_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net552),
    .D(net4548),
    .Q_N(_14921_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[5][3] ));
 sg13g2_dfrbp_1 _35707_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net550),
    .D(net4041),
    .Q_N(_14920_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[5][4] ));
 sg13g2_dfrbp_1 _35708_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net548),
    .D(net3950),
    .Q_N(_14919_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[5][5] ));
 sg13g2_dfrbp_1 _35709_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net546),
    .D(_02301_),
    .Q_N(_14918_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[5][6] ));
 sg13g2_dfrbp_1 _35710_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net544),
    .D(_02302_),
    .Q_N(_14917_),
    .Q(\soc_I.rx_uart_i.fifo_i.ram[5][7] ));
 sg13g2_dfrbp_1 _35711_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net542),
    .D(_02303_),
    .Q_N(_14916_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][0] ));
 sg13g2_dfrbp_1 _35712_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net540),
    .D(_02304_),
    .Q_N(_14915_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][1] ));
 sg13g2_dfrbp_1 _35713_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net538),
    .D(_02305_),
    .Q_N(_14914_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][2] ));
 sg13g2_dfrbp_1 _35714_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net536),
    .D(_02306_),
    .Q_N(_14913_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][3] ));
 sg13g2_dfrbp_1 _35715_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net534),
    .D(_02307_),
    .Q_N(_14912_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][4] ));
 sg13g2_dfrbp_1 _35716_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net532),
    .D(_02308_),
    .Q_N(_14911_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][5] ));
 sg13g2_dfrbp_1 _35717_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net530),
    .D(_02309_),
    .Q_N(_14910_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][6] ));
 sg13g2_dfrbp_1 _35718_ (.CLK(clknet_leaf_319_clk),
    .RESET_B(net528),
    .D(_02310_),
    .Q_N(_14909_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][7] ));
 sg13g2_dfrbp_1 _35719_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net526),
    .D(_02311_),
    .Q_N(_14908_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][8] ));
 sg13g2_dfrbp_1 _35720_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net524),
    .D(_02312_),
    .Q_N(_14907_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][9] ));
 sg13g2_dfrbp_1 _35721_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net522),
    .D(_02313_),
    .Q_N(_14906_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][10] ));
 sg13g2_dfrbp_1 _35722_ (.CLK(clknet_leaf_318_clk),
    .RESET_B(net520),
    .D(_02314_),
    .Q_N(_14905_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][11] ));
 sg13g2_dfrbp_1 _35723_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net518),
    .D(_02315_),
    .Q_N(_14904_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][12] ));
 sg13g2_dfrbp_1 _35724_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net516),
    .D(_02316_),
    .Q_N(_14903_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][13] ));
 sg13g2_dfrbp_1 _35725_ (.CLK(clknet_leaf_301_clk),
    .RESET_B(net514),
    .D(_02317_),
    .Q_N(_14902_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][14] ));
 sg13g2_dfrbp_1 _35726_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net512),
    .D(_02318_),
    .Q_N(_14901_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][15] ));
 sg13g2_dfrbp_1 _35727_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net510),
    .D(_02319_),
    .Q_N(_14900_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][16] ));
 sg13g2_dfrbp_1 _35728_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net508),
    .D(_02320_),
    .Q_N(_14899_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][17] ));
 sg13g2_dfrbp_1 _35729_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net506),
    .D(_02321_),
    .Q_N(_14898_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][18] ));
 sg13g2_dfrbp_1 _35730_ (.CLK(clknet_leaf_289_clk),
    .RESET_B(net504),
    .D(_02322_),
    .Q_N(_14897_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][19] ));
 sg13g2_dfrbp_1 _35731_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net502),
    .D(_02323_),
    .Q_N(_14896_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][20] ));
 sg13g2_dfrbp_1 _35732_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net500),
    .D(_02324_),
    .Q_N(_14895_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][21] ));
 sg13g2_dfrbp_1 _35733_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net498),
    .D(_02325_),
    .Q_N(_14894_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][22] ));
 sg13g2_dfrbp_1 _35734_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net496),
    .D(_02326_),
    .Q_N(_14893_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][23] ));
 sg13g2_dfrbp_1 _35735_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net494),
    .D(_02327_),
    .Q_N(_14892_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][24] ));
 sg13g2_dfrbp_1 _35736_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net492),
    .D(_02328_),
    .Q_N(_14891_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][25] ));
 sg13g2_dfrbp_1 _35737_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net490),
    .D(_02329_),
    .Q_N(_14890_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][26] ));
 sg13g2_dfrbp_1 _35738_ (.CLK(clknet_leaf_295_clk),
    .RESET_B(net488),
    .D(_02330_),
    .Q_N(_14889_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][27] ));
 sg13g2_dfrbp_1 _35739_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net486),
    .D(_02331_),
    .Q_N(_14888_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][28] ));
 sg13g2_dfrbp_1 _35740_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net484),
    .D(_02332_),
    .Q_N(_14887_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][29] ));
 sg13g2_dfrbp_1 _35741_ (.CLK(clknet_leaf_277_clk),
    .RESET_B(net482),
    .D(_02333_),
    .Q_N(_14886_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][30] ));
 sg13g2_dfrbp_1 _35742_ (.CLK(clknet_leaf_286_clk),
    .RESET_B(net480),
    .D(_02334_),
    .Q_N(_14885_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][31] ));
 sg13g2_dfrbp_1 _35743_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net478),
    .D(_02335_),
    .Q_N(_14884_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][0] ));
 sg13g2_dfrbp_1 _35744_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net476),
    .D(_02336_),
    .Q_N(_14883_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][1] ));
 sg13g2_dfrbp_1 _35745_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net474),
    .D(_02337_),
    .Q_N(_14882_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][2] ));
 sg13g2_dfrbp_1 _35746_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net472),
    .D(_02338_),
    .Q_N(_14881_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][3] ));
 sg13g2_dfrbp_1 _35747_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net470),
    .D(_02339_),
    .Q_N(_14880_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][4] ));
 sg13g2_dfrbp_1 _35748_ (.CLK(clknet_leaf_264_clk),
    .RESET_B(net468),
    .D(_02340_),
    .Q_N(_14879_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][5] ));
 sg13g2_dfrbp_1 _35749_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net466),
    .D(_02341_),
    .Q_N(_14878_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][6] ));
 sg13g2_dfrbp_1 _35750_ (.CLK(clknet_leaf_305_clk),
    .RESET_B(net464),
    .D(_02342_),
    .Q_N(_14877_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][7] ));
 sg13g2_dfrbp_1 _35751_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net462),
    .D(_02343_),
    .Q_N(_14876_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][8] ));
 sg13g2_dfrbp_1 _35752_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net460),
    .D(_02344_),
    .Q_N(_14875_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][9] ));
 sg13g2_dfrbp_1 _35753_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net458),
    .D(_02345_),
    .Q_N(_14874_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][10] ));
 sg13g2_dfrbp_1 _35754_ (.CLK(clknet_leaf_317_clk),
    .RESET_B(net456),
    .D(_02346_),
    .Q_N(_14873_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][11] ));
 sg13g2_dfrbp_1 _35755_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net454),
    .D(_02347_),
    .Q_N(_14872_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][12] ));
 sg13g2_dfrbp_1 _35756_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net452),
    .D(_02348_),
    .Q_N(_14871_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][13] ));
 sg13g2_dfrbp_1 _35757_ (.CLK(clknet_leaf_289_clk),
    .RESET_B(net450),
    .D(_02349_),
    .Q_N(_14870_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][14] ));
 sg13g2_dfrbp_1 _35758_ (.CLK(clknet_leaf_310_clk),
    .RESET_B(net448),
    .D(_02350_),
    .Q_N(_14869_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][15] ));
 sg13g2_dfrbp_1 _35759_ (.CLK(clknet_leaf_314_clk),
    .RESET_B(net446),
    .D(_02351_),
    .Q_N(_14868_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][16] ));
 sg13g2_dfrbp_1 _35760_ (.CLK(clknet_leaf_311_clk),
    .RESET_B(net444),
    .D(net3778),
    .Q_N(_14867_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][17] ));
 sg13g2_dfrbp_1 _35761_ (.CLK(clknet_leaf_302_clk),
    .RESET_B(net442),
    .D(_02353_),
    .Q_N(_14866_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][18] ));
 sg13g2_dfrbp_1 _35762_ (.CLK(clknet_leaf_301_clk),
    .RESET_B(net440),
    .D(_02354_),
    .Q_N(_14865_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][19] ));
 sg13g2_dfrbp_1 _35763_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net438),
    .D(_02355_),
    .Q_N(_14864_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][20] ));
 sg13g2_dfrbp_1 _35764_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net436),
    .D(_02356_),
    .Q_N(_14863_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][21] ));
 sg13g2_dfrbp_1 _35765_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net434),
    .D(_02357_),
    .Q_N(_14862_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][22] ));
 sg13g2_dfrbp_1 _35766_ (.CLK(clknet_leaf_307_clk),
    .RESET_B(net432),
    .D(_02358_),
    .Q_N(_14861_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][23] ));
 sg13g2_dfrbp_1 _35767_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net430),
    .D(_02359_),
    .Q_N(_14860_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][24] ));
 sg13g2_dfrbp_1 _35768_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net428),
    .D(_02360_),
    .Q_N(_14859_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][25] ));
 sg13g2_dfrbp_1 _35769_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net426),
    .D(_02361_),
    .Q_N(_14858_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][26] ));
 sg13g2_dfrbp_1 _35770_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net424),
    .D(_02362_),
    .Q_N(_14857_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][27] ));
 sg13g2_dfrbp_1 _35771_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net422),
    .D(_02363_),
    .Q_N(_14856_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][28] ));
 sg13g2_dfrbp_1 _35772_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net420),
    .D(_02364_),
    .Q_N(_14855_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][29] ));
 sg13g2_dfrbp_1 _35773_ (.CLK(clknet_leaf_291_clk),
    .RESET_B(net418),
    .D(_02365_),
    .Q_N(_14854_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][30] ));
 sg13g2_dfrbp_1 _35774_ (.CLK(clknet_leaf_306_clk),
    .RESET_B(net416),
    .D(_02366_),
    .Q_N(_14853_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][31] ));
 sg13g2_dfrbp_1 _35775_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net414),
    .D(_02367_),
    .Q_N(_14852_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][0] ));
 sg13g2_dfrbp_1 _35776_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net412),
    .D(_02368_),
    .Q_N(_14851_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][1] ));
 sg13g2_dfrbp_1 _35777_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net410),
    .D(_02369_),
    .Q_N(_14850_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][2] ));
 sg13g2_dfrbp_1 _35778_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net408),
    .D(_02370_),
    .Q_N(_14849_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][3] ));
 sg13g2_dfrbp_1 _35779_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net406),
    .D(_02371_),
    .Q_N(_14848_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][4] ));
 sg13g2_dfrbp_1 _35780_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net404),
    .D(_02372_),
    .Q_N(_14847_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][5] ));
 sg13g2_dfrbp_1 _35781_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net402),
    .D(_02373_),
    .Q_N(_14846_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][6] ));
 sg13g2_dfrbp_1 _35782_ (.CLK(clknet_leaf_306_clk),
    .RESET_B(net400),
    .D(_02374_),
    .Q_N(_14845_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][7] ));
 sg13g2_dfrbp_1 _35783_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net398),
    .D(_02375_),
    .Q_N(_14844_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][8] ));
 sg13g2_dfrbp_1 _35784_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net396),
    .D(_02376_),
    .Q_N(_14843_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][9] ));
 sg13g2_dfrbp_1 _35785_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net394),
    .D(_02377_),
    .Q_N(_14842_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][10] ));
 sg13g2_dfrbp_1 _35786_ (.CLK(clknet_leaf_315_clk),
    .RESET_B(net392),
    .D(_02378_),
    .Q_N(_14841_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][11] ));
 sg13g2_dfrbp_1 _35787_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net390),
    .D(_02379_),
    .Q_N(_14840_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][12] ));
 sg13g2_dfrbp_1 _35788_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net388),
    .D(_02380_),
    .Q_N(_14839_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][13] ));
 sg13g2_dfrbp_1 _35789_ (.CLK(clknet_leaf_294_clk),
    .RESET_B(net386),
    .D(_02381_),
    .Q_N(_14838_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][14] ));
 sg13g2_dfrbp_1 _35790_ (.CLK(clknet_leaf_309_clk),
    .RESET_B(net384),
    .D(_02382_),
    .Q_N(_14837_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][15] ));
 sg13g2_dfrbp_1 _35791_ (.CLK(clknet_leaf_314_clk),
    .RESET_B(net382),
    .D(_02383_),
    .Q_N(_14836_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][16] ));
 sg13g2_dfrbp_1 _35792_ (.CLK(clknet_leaf_312_clk),
    .RESET_B(net380),
    .D(_02384_),
    .Q_N(_14835_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][17] ));
 sg13g2_dfrbp_1 _35793_ (.CLK(clknet_leaf_308_clk),
    .RESET_B(net378),
    .D(_02385_),
    .Q_N(_14834_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][18] ));
 sg13g2_dfrbp_1 _35794_ (.CLK(clknet_leaf_288_clk),
    .RESET_B(net376),
    .D(_02386_),
    .Q_N(_14833_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][19] ));
 sg13g2_dfrbp_1 _35795_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net374),
    .D(_02387_),
    .Q_N(_14832_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][20] ));
 sg13g2_dfrbp_1 _35796_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net372),
    .D(_02388_),
    .Q_N(_14831_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][21] ));
 sg13g2_dfrbp_1 _35797_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net370),
    .D(_02389_),
    .Q_N(_14830_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][22] ));
 sg13g2_dfrbp_1 _35798_ (.CLK(clknet_leaf_306_clk),
    .RESET_B(net368),
    .D(_02390_),
    .Q_N(_14829_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][23] ));
 sg13g2_dfrbp_1 _35799_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net366),
    .D(_02391_),
    .Q_N(_14828_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][24] ));
 sg13g2_dfrbp_1 _35800_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net364),
    .D(_02392_),
    .Q_N(_14827_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][25] ));
 sg13g2_dfrbp_1 _35801_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net362),
    .D(_02393_),
    .Q_N(_14826_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][26] ));
 sg13g2_dfrbp_1 _35802_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net360),
    .D(_02394_),
    .Q_N(_14825_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][27] ));
 sg13g2_dfrbp_1 _35803_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net358),
    .D(_02395_),
    .Q_N(_14824_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][28] ));
 sg13g2_dfrbp_1 _35804_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net356),
    .D(_02396_),
    .Q_N(_14823_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][29] ));
 sg13g2_dfrbp_1 _35805_ (.CLK(clknet_leaf_291_clk),
    .RESET_B(net354),
    .D(_02397_),
    .Q_N(_14822_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][30] ));
 sg13g2_dfrbp_1 _35806_ (.CLK(clknet_leaf_307_clk),
    .RESET_B(net352),
    .D(_02398_),
    .Q_N(_14821_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][31] ));
 sg13g2_dfrbp_1 _35807_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net350),
    .D(_02399_),
    .Q_N(_14820_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][0] ));
 sg13g2_dfrbp_1 _35808_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net348),
    .D(_02400_),
    .Q_N(_14819_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][1] ));
 sg13g2_dfrbp_1 _35809_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net346),
    .D(_02401_),
    .Q_N(_14818_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][2] ));
 sg13g2_dfrbp_1 _35810_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net344),
    .D(_02402_),
    .Q_N(_14817_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][3] ));
 sg13g2_dfrbp_1 _35811_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net342),
    .D(_02403_),
    .Q_N(_14816_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][4] ));
 sg13g2_dfrbp_1 _35812_ (.CLK(clknet_leaf_263_clk),
    .RESET_B(net340),
    .D(_02404_),
    .Q_N(_14815_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][5] ));
 sg13g2_dfrbp_1 _35813_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net338),
    .D(_02405_),
    .Q_N(_14814_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][6] ));
 sg13g2_dfrbp_1 _35814_ (.CLK(clknet_leaf_323_clk),
    .RESET_B(net285),
    .D(_02406_),
    .Q_N(_14813_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][7] ));
 sg13g2_dfrbp_1 _35815_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net283),
    .D(_02407_),
    .Q_N(_14812_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][8] ));
 sg13g2_dfrbp_1 _35816_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net281),
    .D(_02408_),
    .Q_N(_14811_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][9] ));
 sg13g2_dfrbp_1 _35817_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net279),
    .D(_02409_),
    .Q_N(_14810_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][10] ));
 sg13g2_dfrbp_1 _35818_ (.CLK(clknet_leaf_322_clk),
    .RESET_B(net277),
    .D(_02410_),
    .Q_N(_14809_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][11] ));
 sg13g2_dfrbp_1 _35819_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net275),
    .D(_02411_),
    .Q_N(_14808_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][12] ));
 sg13g2_dfrbp_1 _35820_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net273),
    .D(_02412_),
    .Q_N(_14807_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][13] ));
 sg13g2_dfrbp_1 _35821_ (.CLK(clknet_leaf_278_clk),
    .RESET_B(net271),
    .D(_02413_),
    .Q_N(_14806_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][14] ));
 sg13g2_dfrbp_1 _35822_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net269),
    .D(_02414_),
    .Q_N(_14805_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][15] ));
 sg13g2_dfrbp_1 _35823_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net263),
    .D(_02415_),
    .Q_N(_14804_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][16] ));
 sg13g2_dfrbp_1 _35824_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net261),
    .D(_02416_),
    .Q_N(_14803_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][17] ));
 sg13g2_dfrbp_1 _35825_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net259),
    .D(_02417_),
    .Q_N(_14802_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][18] ));
 sg13g2_dfrbp_1 _35826_ (.CLK(clknet_leaf_300_clk),
    .RESET_B(net257),
    .D(_02418_),
    .Q_N(_14801_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][19] ));
 sg13g2_dfrbp_1 _35827_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net255),
    .D(_02419_),
    .Q_N(_14800_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][20] ));
 sg13g2_dfrbp_1 _35828_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net253),
    .D(_02420_),
    .Q_N(_14799_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][21] ));
 sg13g2_dfrbp_1 _35829_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net251),
    .D(_02421_),
    .Q_N(_14798_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][22] ));
 sg13g2_dfrbp_1 _35830_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net249),
    .D(_02422_),
    .Q_N(_14797_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][23] ));
 sg13g2_dfrbp_1 _35831_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net247),
    .D(_02423_),
    .Q_N(_14796_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][24] ));
 sg13g2_dfrbp_1 _35832_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net245),
    .D(_02424_),
    .Q_N(_14795_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][25] ));
 sg13g2_dfrbp_1 _35833_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net243),
    .D(_02425_),
    .Q_N(_14794_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][26] ));
 sg13g2_dfrbp_1 _35834_ (.CLK(clknet_leaf_296_clk),
    .RESET_B(net241),
    .D(_02426_),
    .Q_N(_14793_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][27] ));
 sg13g2_dfrbp_1 _35835_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net239),
    .D(_02427_),
    .Q_N(_14792_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][28] ));
 sg13g2_dfrbp_1 _35836_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net237),
    .D(_02428_),
    .Q_N(_14791_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][29] ));
 sg13g2_dfrbp_1 _35837_ (.CLK(clknet_leaf_296_clk),
    .RESET_B(net235),
    .D(_02429_),
    .Q_N(_14790_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][30] ));
 sg13g2_dfrbp_1 _35838_ (.CLK(clknet_leaf_308_clk),
    .RESET_B(net233),
    .D(_02430_),
    .Q_N(_14789_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][31] ));
 sg13g2_dfrbp_1 _35839_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net231),
    .D(_02431_),
    .Q_N(_14788_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][0] ));
 sg13g2_dfrbp_1 _35840_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net229),
    .D(_02432_),
    .Q_N(_14787_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][1] ));
 sg13g2_dfrbp_1 _35841_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net227),
    .D(_02433_),
    .Q_N(_14786_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][2] ));
 sg13g2_dfrbp_1 _35842_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net225),
    .D(_02434_),
    .Q_N(_14785_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][3] ));
 sg13g2_dfrbp_1 _35843_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net223),
    .D(_02435_),
    .Q_N(_14784_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][4] ));
 sg13g2_dfrbp_1 _35844_ (.CLK(clknet_leaf_264_clk),
    .RESET_B(net221),
    .D(_02436_),
    .Q_N(_14783_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][5] ));
 sg13g2_dfrbp_1 _35845_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net219),
    .D(_02437_),
    .Q_N(_14782_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][6] ));
 sg13g2_dfrbp_1 _35846_ (.CLK(clknet_leaf_321_clk),
    .RESET_B(net217),
    .D(_02438_),
    .Q_N(_14781_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][7] ));
 sg13g2_dfrbp_1 _35847_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net215),
    .D(_02439_),
    .Q_N(_14780_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][8] ));
 sg13g2_dfrbp_1 _35848_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net213),
    .D(_02440_),
    .Q_N(_14779_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][9] ));
 sg13g2_dfrbp_1 _35849_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net211),
    .D(_02441_),
    .Q_N(_14778_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][10] ));
 sg13g2_dfrbp_1 _35850_ (.CLK(clknet_leaf_322_clk),
    .RESET_B(net209),
    .D(_02442_),
    .Q_N(_14777_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][11] ));
 sg13g2_dfrbp_1 _35851_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net207),
    .D(_02443_),
    .Q_N(_14776_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][12] ));
 sg13g2_dfrbp_1 _35852_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net205),
    .D(_02444_),
    .Q_N(_14775_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][13] ));
 sg13g2_dfrbp_1 _35853_ (.CLK(clknet_leaf_295_clk),
    .RESET_B(net203),
    .D(_02445_),
    .Q_N(_14774_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][14] ));
 sg13g2_dfrbp_1 _35854_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net201),
    .D(_02446_),
    .Q_N(_14773_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][15] ));
 sg13g2_dfrbp_1 _35855_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net199),
    .D(_02447_),
    .Q_N(_14772_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][16] ));
 sg13g2_dfrbp_1 _35856_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net197),
    .D(_02448_),
    .Q_N(_14771_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][17] ));
 sg13g2_dfrbp_1 _35857_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net195),
    .D(_02449_),
    .Q_N(_14770_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][18] ));
 sg13g2_dfrbp_1 _35858_ (.CLK(clknet_leaf_299_clk),
    .RESET_B(net193),
    .D(_02450_),
    .Q_N(_14769_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][19] ));
 sg13g2_dfrbp_1 _35859_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net191),
    .D(_02451_),
    .Q_N(_14768_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][20] ));
 sg13g2_dfrbp_1 _35860_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net189),
    .D(_02452_),
    .Q_N(_14767_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][21] ));
 sg13g2_dfrbp_1 _35861_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net187),
    .D(_02453_),
    .Q_N(_14766_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][22] ));
 sg13g2_dfrbp_1 _35862_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net185),
    .D(_02454_),
    .Q_N(_14765_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][23] ));
 sg13g2_dfrbp_1 _35863_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net183),
    .D(_02455_),
    .Q_N(_14764_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][24] ));
 sg13g2_dfrbp_1 _35864_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net181),
    .D(_02456_),
    .Q_N(_14763_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][25] ));
 sg13g2_dfrbp_1 _35865_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net179),
    .D(_02457_),
    .Q_N(_14762_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][26] ));
 sg13g2_dfrbp_1 _35866_ (.CLK(clknet_leaf_296_clk),
    .RESET_B(net177),
    .D(_02458_),
    .Q_N(_14761_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][27] ));
 sg13g2_dfrbp_1 _35867_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net175),
    .D(_02459_),
    .Q_N(_14760_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][28] ));
 sg13g2_dfrbp_1 _35868_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net173),
    .D(_02460_),
    .Q_N(_14759_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][29] ));
 sg13g2_dfrbp_1 _35869_ (.CLK(clknet_leaf_298_clk),
    .RESET_B(net171),
    .D(_02461_),
    .Q_N(_14758_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][30] ));
 sg13g2_dfrbp_1 _35870_ (.CLK(clknet_leaf_309_clk),
    .RESET_B(net169),
    .D(_02462_),
    .Q_N(_14757_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][31] ));
 sg13g2_dfrbp_1 _35871_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net167),
    .D(_02463_),
    .Q_N(_14756_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][0] ));
 sg13g2_dfrbp_1 _35872_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net165),
    .D(_02464_),
    .Q_N(_14755_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][1] ));
 sg13g2_dfrbp_1 _35873_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net163),
    .D(_02465_),
    .Q_N(_14754_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][2] ));
 sg13g2_dfrbp_1 _35874_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net161),
    .D(_02466_),
    .Q_N(_14753_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][3] ));
 sg13g2_dfrbp_1 _35875_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net159),
    .D(_02467_),
    .Q_N(_14752_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][4] ));
 sg13g2_dfrbp_1 _35876_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net157),
    .D(_02468_),
    .Q_N(_14751_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][5] ));
 sg13g2_dfrbp_1 _35877_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net155),
    .D(_02469_),
    .Q_N(_14750_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][6] ));
 sg13g2_dfrbp_1 _35878_ (.CLK(clknet_leaf_320_clk),
    .RESET_B(net153),
    .D(_02470_),
    .Q_N(_14749_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][7] ));
 sg13g2_dfrbp_1 _35879_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net151),
    .D(_02471_),
    .Q_N(_14748_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][8] ));
 sg13g2_dfrbp_1 _35880_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net149),
    .D(_02472_),
    .Q_N(_14747_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][9] ));
 sg13g2_dfrbp_1 _35881_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net147),
    .D(_02473_),
    .Q_N(_14746_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][10] ));
 sg13g2_dfrbp_1 _35882_ (.CLK(clknet_leaf_322_clk),
    .RESET_B(net145),
    .D(_02474_),
    .Q_N(_14745_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][11] ));
 sg13g2_dfrbp_1 _35883_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net143),
    .D(_02475_),
    .Q_N(_14744_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][12] ));
 sg13g2_dfrbp_1 _35884_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net141),
    .D(_02476_),
    .Q_N(_14743_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][13] ));
 sg13g2_dfrbp_1 _35885_ (.CLK(clknet_leaf_293_clk),
    .RESET_B(net139),
    .D(_02477_),
    .Q_N(_14742_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][14] ));
 sg13g2_dfrbp_1 _35886_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net137),
    .D(_02478_),
    .Q_N(_14741_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][15] ));
 sg13g2_dfrbp_1 _35887_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net135),
    .D(_02479_),
    .Q_N(_14740_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][16] ));
 sg13g2_dfrbp_1 _35888_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net133),
    .D(_02480_),
    .Q_N(_14739_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][17] ));
 sg13g2_dfrbp_1 _35889_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net131),
    .D(_02481_),
    .Q_N(_14738_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][18] ));
 sg13g2_dfrbp_1 _35890_ (.CLK(clknet_leaf_303_clk),
    .RESET_B(net129),
    .D(_02482_),
    .Q_N(_14737_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][19] ));
 sg13g2_dfrbp_1 _35891_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net127),
    .D(_02483_),
    .Q_N(_14736_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][20] ));
 sg13g2_dfrbp_1 _35892_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net125),
    .D(_02484_),
    .Q_N(_14735_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][21] ));
 sg13g2_dfrbp_1 _35893_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net123),
    .D(_02485_),
    .Q_N(_14734_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][22] ));
 sg13g2_dfrbp_1 _35894_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net121),
    .D(_02486_),
    .Q_N(_14733_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][23] ));
 sg13g2_dfrbp_1 _35895_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net118),
    .D(_02487_),
    .Q_N(_14732_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][24] ));
 sg13g2_dfrbp_1 _35896_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net116),
    .D(_02488_),
    .Q_N(_14731_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][25] ));
 sg13g2_dfrbp_1 _35897_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net114),
    .D(_02489_),
    .Q_N(_14730_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][26] ));
 sg13g2_dfrbp_1 _35898_ (.CLK(clknet_leaf_297_clk),
    .RESET_B(net112),
    .D(_02490_),
    .Q_N(_14729_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][27] ));
 sg13g2_dfrbp_1 _35899_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net110),
    .D(_02491_),
    .Q_N(_14728_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][28] ));
 sg13g2_dfrbp_1 _35900_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net108),
    .D(_02492_),
    .Q_N(_14727_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][29] ));
 sg13g2_dfrbp_1 _35901_ (.CLK(clknet_leaf_297_clk),
    .RESET_B(net106),
    .D(_02493_),
    .Q_N(_14726_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][30] ));
 sg13g2_dfrbp_1 _35902_ (.CLK(clknet_leaf_286_clk),
    .RESET_B(net104),
    .D(_02494_),
    .Q_N(_14725_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][31] ));
 sg13g2_dfrbp_1 _35903_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net70),
    .D(_02495_),
    .Q_N(_14724_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][0] ));
 sg13g2_dfrbp_1 _35904_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net68),
    .D(_02496_),
    .Q_N(_14723_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][1] ));
 sg13g2_dfrbp_1 _35905_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net66),
    .D(_02497_),
    .Q_N(_14722_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][2] ));
 sg13g2_dfrbp_1 _35906_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net64),
    .D(_02498_),
    .Q_N(_14721_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][3] ));
 sg13g2_dfrbp_1 _35907_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net62),
    .D(_02499_),
    .Q_N(_14720_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][4] ));
 sg13g2_dfrbp_1 _35908_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net60),
    .D(_02500_),
    .Q_N(_14719_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][5] ));
 sg13g2_dfrbp_1 _35909_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net58),
    .D(_02501_),
    .Q_N(_14718_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][6] ));
 sg13g2_dfrbp_1 _35910_ (.CLK(clknet_leaf_308_clk),
    .RESET_B(net56),
    .D(_02502_),
    .Q_N(_14717_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][7] ));
 sg13g2_dfrbp_1 _35911_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net54),
    .D(_02503_),
    .Q_N(_14716_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][8] ));
 sg13g2_dfrbp_1 _35912_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net52),
    .D(_02504_),
    .Q_N(_14715_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][9] ));
 sg13g2_dfrbp_1 _35913_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net50),
    .D(_02505_),
    .Q_N(_14714_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][10] ));
 sg13g2_dfrbp_1 _35914_ (.CLK(clknet_leaf_316_clk),
    .RESET_B(net48),
    .D(_02506_),
    .Q_N(_14713_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][11] ));
 sg13g2_dfrbp_1 _35915_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net46),
    .D(_02507_),
    .Q_N(_14712_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][12] ));
 sg13g2_dfrbp_1 _35916_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net44),
    .D(_02508_),
    .Q_N(_14711_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][13] ));
 sg13g2_dfrbp_1 _35917_ (.CLK(clknet_leaf_299_clk),
    .RESET_B(net42),
    .D(_02509_),
    .Q_N(_14710_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][14] ));
 sg13g2_dfrbp_1 _35918_ (.CLK(clknet_leaf_310_clk),
    .RESET_B(net40),
    .D(_02510_),
    .Q_N(_14709_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][15] ));
 sg13g2_dfrbp_1 _35919_ (.CLK(clknet_leaf_316_clk),
    .RESET_B(net38),
    .D(_02511_),
    .Q_N(_14708_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][16] ));
 sg13g2_dfrbp_1 _35920_ (.CLK(clknet_leaf_314_clk),
    .RESET_B(net36),
    .D(_02512_),
    .Q_N(_14707_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][17] ));
 sg13g2_dfrbp_1 _35921_ (.CLK(clknet_leaf_303_clk),
    .RESET_B(net34),
    .D(_02513_),
    .Q_N(_14706_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][18] ));
 sg13g2_dfrbp_1 _35922_ (.CLK(clknet_leaf_303_clk),
    .RESET_B(net32),
    .D(_02514_),
    .Q_N(_14705_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][19] ));
 sg13g2_dfrbp_1 _35923_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net30),
    .D(_02515_),
    .Q_N(_14704_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][20] ));
 sg13g2_dfrbp_1 _35924_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net28),
    .D(_02516_),
    .Q_N(_14703_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][21] ));
 sg13g2_dfrbp_1 _35925_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net26),
    .D(_02517_),
    .Q_N(_14702_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][22] ));
 sg13g2_dfrbp_1 _35926_ (.CLK(clknet_leaf_309_clk),
    .RESET_B(net24),
    .D(_02518_),
    .Q_N(_14701_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][23] ));
 sg13g2_dfrbp_1 _35927_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net22),
    .D(_02519_),
    .Q_N(_14700_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][24] ));
 sg13g2_dfrbp_1 _35928_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net20),
    .D(_02520_),
    .Q_N(_14699_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][25] ));
 sg13g2_dfrbp_1 _35929_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net18),
    .D(_02521_),
    .Q_N(_14698_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][26] ));
 sg13g2_dfrbp_1 _35930_ (.CLK(clknet_leaf_296_clk),
    .RESET_B(net16),
    .D(_02522_),
    .Q_N(_14697_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][27] ));
 sg13g2_dfrbp_1 _35931_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net14),
    .D(_02523_),
    .Q_N(_14696_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][28] ));
 sg13g2_dfrbp_1 _35932_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net2592),
    .D(_02524_),
    .Q_N(_14695_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][29] ));
 sg13g2_dfrbp_1 _35933_ (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2590),
    .D(_02525_),
    .Q_N(_14694_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][30] ));
 sg13g2_dfrbp_1 _35934_ (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2334),
    .D(_02526_),
    .Q_N(_16753_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][31] ));
 sg13g2_dfrbp_1 _35935_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2335),
    .D(_00004_),
    .Q_N(_00243_),
    .Q(\soc_I.qqspi_I.state[0] ));
 sg13g2_dfrbp_1 _35936_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2336),
    .D(_00005_),
    .Q_N(_16754_),
    .Q(\soc_I.qqspi_I.state[1] ));
 sg13g2_dfrbp_1 _35937_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2337),
    .D(_00006_),
    .Q_N(_16755_),
    .Q(\soc_I.qqspi_I.state[2] ));
 sg13g2_dfrbp_1 _35938_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2338),
    .D(_00007_),
    .Q_N(_16756_),
    .Q(\soc_I.qqspi_I.state[3] ));
 sg13g2_dfrbp_1 _35939_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2339),
    .D(net3106),
    .Q_N(_00150_),
    .Q(\soc_I.qqspi_I.state[4] ));
 sg13g2_dfrbp_1 _35940_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2447),
    .D(_00009_),
    .Q_N(_00291_),
    .Q(\soc_I.qqspi_I.state[5] ));
 sg13g2_dfrbp_1 _35941_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net2588),
    .D(_00010_),
    .Q_N(_00242_),
    .Q(\soc_I.qqspi_I.state[6] ));
 sg13g2_dfrbp_1 _35942_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net2586),
    .D(_02527_),
    .Q_N(_14693_),
    .Q(\soc_I.tx_uart_i.state[0] ));
 sg13g2_dfrbp_1 _35943_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net2582),
    .D(_02528_),
    .Q_N(_14692_),
    .Q(\soc_I.tx_uart_i.state[1] ));
 sg13g2_dfrbp_1 _35944_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net2578),
    .D(_02529_),
    .Q_N(_14691_),
    .Q(\soc_I.qqspi_I.spi_buf[8] ));
 sg13g2_dfrbp_1 _35945_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net2569),
    .D(_02530_),
    .Q_N(_14690_),
    .Q(\soc_I.qqspi_I.spi_buf[9] ));
 sg13g2_dfrbp_1 _35946_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2565),
    .D(_02531_),
    .Q_N(_14689_),
    .Q(\soc_I.qqspi_I.spi_buf[10] ));
 sg13g2_dfrbp_1 _35947_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net2561),
    .D(_02532_),
    .Q_N(_14688_),
    .Q(\soc_I.qqspi_I.spi_buf[11] ));
 sg13g2_dfrbp_1 _35948_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2557),
    .D(_02533_),
    .Q_N(_14687_),
    .Q(\soc_I.qqspi_I.spi_buf[12] ));
 sg13g2_dfrbp_1 _35949_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net2521),
    .D(_02534_),
    .Q_N(_14686_),
    .Q(\soc_I.qqspi_I.spi_buf[13] ));
 sg13g2_dfrbp_1 _35950_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net2517),
    .D(_02535_),
    .Q_N(_14685_),
    .Q(\soc_I.qqspi_I.spi_buf[14] ));
 sg13g2_dfrbp_1 _35951_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2513),
    .D(_02536_),
    .Q_N(_14684_),
    .Q(\soc_I.qqspi_I.spi_buf[15] ));
 sg13g2_dfrbp_1 _35952_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2509),
    .D(_02537_),
    .Q_N(_14683_),
    .Q(\soc_I.qqspi_I.spi_buf[16] ));
 sg13g2_dfrbp_1 _35953_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2505),
    .D(_02538_),
    .Q_N(_14682_),
    .Q(\soc_I.qqspi_I.spi_buf[17] ));
 sg13g2_dfrbp_1 _35954_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2501),
    .D(_02539_),
    .Q_N(_14681_),
    .Q(\soc_I.qqspi_I.spi_buf[18] ));
 sg13g2_dfrbp_1 _35955_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2497),
    .D(_02540_),
    .Q_N(_14680_),
    .Q(\soc_I.qqspi_I.spi_buf[19] ));
 sg13g2_dfrbp_1 _35956_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2493),
    .D(_02541_),
    .Q_N(_14679_),
    .Q(\soc_I.qqspi_I.spi_buf[20] ));
 sg13g2_dfrbp_1 _35957_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net2489),
    .D(_02542_),
    .Q_N(_14678_),
    .Q(\soc_I.qqspi_I.spi_buf[21] ));
 sg13g2_dfrbp_1 _35958_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net2485),
    .D(_02543_),
    .Q_N(_14677_),
    .Q(\soc_I.qqspi_I.spi_buf[22] ));
 sg13g2_dfrbp_1 _35959_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2481),
    .D(_02544_),
    .Q_N(_14676_),
    .Q(\soc_I.qqspi_I.spi_buf[23] ));
 sg13g2_dfrbp_1 _35960_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2477),
    .D(_02545_),
    .Q_N(_14675_),
    .Q(\soc_I.qqspi_I.spi_buf[0] ));
 sg13g2_dfrbp_1 _35961_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net2473),
    .D(_02546_),
    .Q_N(_14674_),
    .Q(\soc_I.qqspi_I.spi_buf[1] ));
 sg13g2_dfrbp_1 _35962_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net2469),
    .D(_02547_),
    .Q_N(_14673_),
    .Q(\soc_I.qqspi_I.spi_buf[2] ));
 sg13g2_dfrbp_1 _35963_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net2465),
    .D(_02548_),
    .Q_N(_14672_),
    .Q(\soc_I.qqspi_I.spi_buf[3] ));
 sg13g2_dfrbp_1 _35964_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net2461),
    .D(_02549_),
    .Q_N(_14671_),
    .Q(\soc_I.qqspi_I.spi_buf[4] ));
 sg13g2_dfrbp_1 _35965_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net2457),
    .D(_02550_),
    .Q_N(_14670_),
    .Q(\soc_I.qqspi_I.spi_buf[5] ));
 sg13g2_dfrbp_1 _35966_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net2453),
    .D(_02551_),
    .Q_N(_14669_),
    .Q(\soc_I.qqspi_I.spi_buf[6] ));
 sg13g2_dfrbp_1 _35967_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2449),
    .D(net5349),
    .Q_N(_14668_),
    .Q(\soc_I.qqspi_I.spi_buf[7] ));
 sg13g2_dfrbp_1 _35968_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2445),
    .D(_02553_),
    .Q_N(_14667_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][0] ));
 sg13g2_dfrbp_1 _35969_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2440),
    .D(_02554_),
    .Q_N(_14666_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][1] ));
 sg13g2_dfrbp_1 _35970_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2438),
    .D(_02555_),
    .Q_N(_14665_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][2] ));
 sg13g2_dfrbp_1 _35971_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2435),
    .D(_02556_),
    .Q_N(_14664_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][3] ));
 sg13g2_dfrbp_1 _35972_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2433),
    .D(_02557_),
    .Q_N(_14663_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][4] ));
 sg13g2_dfrbp_1 _35973_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2431),
    .D(_02558_),
    .Q_N(_14662_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][5] ));
 sg13g2_dfrbp_1 _35974_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2429),
    .D(_02559_),
    .Q_N(_14661_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][6] ));
 sg13g2_dfrbp_1 _35975_ (.CLK(clknet_leaf_304_clk),
    .RESET_B(net2427),
    .D(_02560_),
    .Q_N(_14660_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][7] ));
 sg13g2_dfrbp_1 _35976_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2425),
    .D(_02561_),
    .Q_N(_14659_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][8] ));
 sg13g2_dfrbp_1 _35977_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2423),
    .D(_02562_),
    .Q_N(_14658_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][9] ));
 sg13g2_dfrbp_1 _35978_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2421),
    .D(_02563_),
    .Q_N(_14657_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][10] ));
 sg13g2_dfrbp_1 _35979_ (.CLK(clknet_leaf_313_clk),
    .RESET_B(net2419),
    .D(_02564_),
    .Q_N(_14656_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][11] ));
 sg13g2_dfrbp_1 _35980_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2417),
    .D(_02565_),
    .Q_N(_14655_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][12] ));
 sg13g2_dfrbp_1 _35981_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2415),
    .D(_02566_),
    .Q_N(_14654_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][13] ));
 sg13g2_dfrbp_1 _35982_ (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2317),
    .D(_02567_),
    .Q_N(_14653_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][14] ));
 sg13g2_dfrbp_1 _35983_ (.CLK(clknet_leaf_309_clk),
    .RESET_B(net2313),
    .D(_02568_),
    .Q_N(_14652_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][15] ));
 sg13g2_dfrbp_1 _35984_ (.CLK(clknet_leaf_319_clk),
    .RESET_B(net2309),
    .D(_02569_),
    .Q_N(_14651_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][16] ));
 sg13g2_dfrbp_1 _35985_ (.CLK(clknet_leaf_313_clk),
    .RESET_B(net2305),
    .D(_02570_),
    .Q_N(_14650_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][17] ));
 sg13g2_dfrbp_1 _35986_ (.CLK(clknet_leaf_304_clk),
    .RESET_B(net2301),
    .D(_02571_),
    .Q_N(_14649_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][18] ));
 sg13g2_dfrbp_1 _35987_ (.CLK(clknet_leaf_303_clk),
    .RESET_B(net2297),
    .D(_02572_),
    .Q_N(_14648_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][19] ));
 sg13g2_dfrbp_1 _35988_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2293),
    .D(_02573_),
    .Q_N(_14647_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][20] ));
 sg13g2_dfrbp_1 _35989_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net2289),
    .D(_02574_),
    .Q_N(_14646_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][21] ));
 sg13g2_dfrbp_1 _35990_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2285),
    .D(_02575_),
    .Q_N(_14645_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][22] ));
 sg13g2_dfrbp_1 _35991_ (.CLK(clknet_leaf_306_clk),
    .RESET_B(net2281),
    .D(_02576_),
    .Q_N(_14644_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][23] ));
 sg13g2_dfrbp_1 _35992_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2277),
    .D(_02577_),
    .Q_N(_14643_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][24] ));
 sg13g2_dfrbp_1 _35993_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2137),
    .D(_02578_),
    .Q_N(_14642_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][25] ));
 sg13g2_dfrbp_1 _35994_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2133),
    .D(_02579_),
    .Q_N(_14641_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][26] ));
 sg13g2_dfrbp_1 _35995_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2001),
    .D(_02580_),
    .Q_N(_14640_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][27] ));
 sg13g2_dfrbp_1 _35996_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1725),
    .D(_02581_),
    .Q_N(_14639_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][28] ));
 sg13g2_dfrbp_1 _35997_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1721),
    .D(_02582_),
    .Q_N(_14638_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][29] ));
 sg13g2_dfrbp_1 _35998_ (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1717),
    .D(_02583_),
    .Q_N(_14637_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][30] ));
 sg13g2_dfrbp_1 _35999_ (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1713),
    .D(_02584_),
    .Q_N(_14636_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][31] ));
 sg13g2_dfrbp_1 _36000_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1709),
    .D(_02585_),
    .Q_N(_14635_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][0] ));
 sg13g2_dfrbp_1 _36001_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1705),
    .D(_02586_),
    .Q_N(_14634_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][1] ));
 sg13g2_dfrbp_1 _36002_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1701),
    .D(_02587_),
    .Q_N(_14633_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][2] ));
 sg13g2_dfrbp_1 _36003_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1697),
    .D(_02588_),
    .Q_N(_14632_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][3] ));
 sg13g2_dfrbp_1 _36004_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1693),
    .D(_02589_),
    .Q_N(_14631_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][4] ));
 sg13g2_dfrbp_1 _36005_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1689),
    .D(_02590_),
    .Q_N(_14630_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][5] ));
 sg13g2_dfrbp_1 _36006_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1685),
    .D(_02591_),
    .Q_N(_14629_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][6] ));
 sg13g2_dfrbp_1 _36007_ (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1681),
    .D(_02592_),
    .Q_N(_14628_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][7] ));
 sg13g2_dfrbp_1 _36008_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1677),
    .D(_02593_),
    .Q_N(_14627_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][8] ));
 sg13g2_dfrbp_1 _36009_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1673),
    .D(_02594_),
    .Q_N(_14626_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][9] ));
 sg13g2_dfrbp_1 _36010_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1665),
    .D(_02595_),
    .Q_N(_14625_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][10] ));
 sg13g2_dfrbp_1 _36011_ (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1661),
    .D(_02596_),
    .Q_N(_14624_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][11] ));
 sg13g2_dfrbp_1 _36012_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1657),
    .D(_02597_),
    .Q_N(_14623_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][12] ));
 sg13g2_dfrbp_1 _36013_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1653),
    .D(_02598_),
    .Q_N(_14622_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][13] ));
 sg13g2_dfrbp_1 _36014_ (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1649),
    .D(_02599_),
    .Q_N(_14621_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][14] ));
 sg13g2_dfrbp_1 _36015_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1645),
    .D(_02600_),
    .Q_N(_14620_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][15] ));
 sg13g2_dfrbp_1 _36016_ (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1641),
    .D(_02601_),
    .Q_N(_14619_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][16] ));
 sg13g2_dfrbp_1 _36017_ (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1637),
    .D(_02602_),
    .Q_N(_14618_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][17] ));
 sg13g2_dfrbp_1 _36018_ (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1633),
    .D(_02603_),
    .Q_N(_14617_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][18] ));
 sg13g2_dfrbp_1 _36019_ (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1629),
    .D(_02604_),
    .Q_N(_14616_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][19] ));
 sg13g2_dfrbp_1 _36020_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1625),
    .D(_02605_),
    .Q_N(_14615_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][20] ));
 sg13g2_dfrbp_1 _36021_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1621),
    .D(_02606_),
    .Q_N(_14614_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][21] ));
 sg13g2_dfrbp_1 _36022_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1617),
    .D(_02607_),
    .Q_N(_14613_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][22] ));
 sg13g2_dfrbp_1 _36023_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1613),
    .D(_02608_),
    .Q_N(_14612_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][23] ));
 sg13g2_dfrbp_1 _36024_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1609),
    .D(_02609_),
    .Q_N(_14611_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][24] ));
 sg13g2_dfrbp_1 _36025_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1605),
    .D(_02610_),
    .Q_N(_14610_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][25] ));
 sg13g2_dfrbp_1 _36026_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1601),
    .D(_02611_),
    .Q_N(_14609_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][26] ));
 sg13g2_dfrbp_1 _36027_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1597),
    .D(_02612_),
    .Q_N(_14608_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][27] ));
 sg13g2_dfrbp_1 _36028_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1593),
    .D(_02613_),
    .Q_N(_14607_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][28] ));
 sg13g2_dfrbp_1 _36029_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1589),
    .D(_02614_),
    .Q_N(_14606_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][29] ));
 sg13g2_dfrbp_1 _36030_ (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1585),
    .D(_02615_),
    .Q_N(_14605_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][30] ));
 sg13g2_dfrbp_1 _36031_ (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1581),
    .D(_02616_),
    .Q_N(_14604_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][31] ));
 sg13g2_dfrbp_1 _36032_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1577),
    .D(_02617_),
    .Q_N(_14603_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][0] ));
 sg13g2_dfrbp_1 _36033_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1573),
    .D(_02618_),
    .Q_N(_14602_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][1] ));
 sg13g2_dfrbp_1 _36034_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1569),
    .D(_02619_),
    .Q_N(_14601_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][2] ));
 sg13g2_dfrbp_1 _36035_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1565),
    .D(_02620_),
    .Q_N(_14600_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][3] ));
 sg13g2_dfrbp_1 _36036_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1561),
    .D(_02621_),
    .Q_N(_14599_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][4] ));
 sg13g2_dfrbp_1 _36037_ (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1557),
    .D(_02622_),
    .Q_N(_14598_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][5] ));
 sg13g2_dfrbp_1 _36038_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1553),
    .D(_02623_),
    .Q_N(_14597_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][6] ));
 sg13g2_dfrbp_1 _36039_ (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1549),
    .D(_02624_),
    .Q_N(_14596_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][7] ));
 sg13g2_dfrbp_1 _36040_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1545),
    .D(_02625_),
    .Q_N(_14595_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][8] ));
 sg13g2_dfrbp_1 _36041_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1541),
    .D(_02626_),
    .Q_N(_14594_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][9] ));
 sg13g2_dfrbp_1 _36042_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1535),
    .D(_02627_),
    .Q_N(_14593_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][10] ));
 sg13g2_dfrbp_1 _36043_ (.CLK(clknet_leaf_319_clk),
    .RESET_B(net1531),
    .D(_02628_),
    .Q_N(_14592_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][11] ));
 sg13g2_dfrbp_1 _36044_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1527),
    .D(_02629_),
    .Q_N(_14591_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][12] ));
 sg13g2_dfrbp_1 _36045_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1523),
    .D(_02630_),
    .Q_N(_14590_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][13] ));
 sg13g2_dfrbp_1 _36046_ (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1519),
    .D(_02631_),
    .Q_N(_14589_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][14] ));
 sg13g2_dfrbp_1 _36047_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1515),
    .D(_02632_),
    .Q_N(_14588_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][15] ));
 sg13g2_dfrbp_1 _36048_ (.CLK(clknet_leaf_320_clk),
    .RESET_B(net1511),
    .D(_02633_),
    .Q_N(_14587_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][16] ));
 sg13g2_dfrbp_1 _36049_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1507),
    .D(_02634_),
    .Q_N(_14586_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][17] ));
 sg13g2_dfrbp_1 _36050_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1503),
    .D(_02635_),
    .Q_N(_14585_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][18] ));
 sg13g2_dfrbp_1 _36051_ (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1499),
    .D(_02636_),
    .Q_N(_14584_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][19] ));
 sg13g2_dfrbp_1 _36052_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1495),
    .D(_02637_),
    .Q_N(_14583_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][20] ));
 sg13g2_dfrbp_1 _36053_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1491),
    .D(_02638_),
    .Q_N(_14582_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][21] ));
 sg13g2_dfrbp_1 _36054_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1487),
    .D(_02639_),
    .Q_N(_14581_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][22] ));
 sg13g2_dfrbp_1 _36055_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1483),
    .D(_02640_),
    .Q_N(_14580_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][23] ));
 sg13g2_dfrbp_1 _36056_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1479),
    .D(_02641_),
    .Q_N(_14579_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][24] ));
 sg13g2_dfrbp_1 _36057_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1475),
    .D(_02642_),
    .Q_N(_14578_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][25] ));
 sg13g2_dfrbp_1 _36058_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1471),
    .D(_02643_),
    .Q_N(_14577_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][26] ));
 sg13g2_dfrbp_1 _36059_ (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1467),
    .D(_02644_),
    .Q_N(_14576_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][27] ));
 sg13g2_dfrbp_1 _36060_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1463),
    .D(_02645_),
    .Q_N(_14575_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][28] ));
 sg13g2_dfrbp_1 _36061_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1459),
    .D(_02646_),
    .Q_N(_14574_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][29] ));
 sg13g2_dfrbp_1 _36062_ (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1455),
    .D(_02647_),
    .Q_N(_14573_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][30] ));
 sg13g2_dfrbp_1 _36063_ (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1451),
    .D(_02648_),
    .Q_N(_14572_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][31] ));
 sg13g2_dfrbp_1 _36064_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1447),
    .D(_02649_),
    .Q_N(_14571_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][0] ));
 sg13g2_dfrbp_1 _36065_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1443),
    .D(_02650_),
    .Q_N(_14570_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][1] ));
 sg13g2_dfrbp_1 _36066_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1439),
    .D(_02651_),
    .Q_N(_14569_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][2] ));
 sg13g2_dfrbp_1 _36067_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1435),
    .D(_02652_),
    .Q_N(_14568_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][3] ));
 sg13g2_dfrbp_1 _36068_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1431),
    .D(_02653_),
    .Q_N(_14567_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][4] ));
 sg13g2_dfrbp_1 _36069_ (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1427),
    .D(_02654_),
    .Q_N(_14566_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][5] ));
 sg13g2_dfrbp_1 _36070_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1423),
    .D(_02655_),
    .Q_N(_14565_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][6] ));
 sg13g2_dfrbp_1 _36071_ (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1419),
    .D(_02656_),
    .Q_N(_14564_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][7] ));
 sg13g2_dfrbp_1 _36072_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1415),
    .D(_02657_),
    .Q_N(_14563_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][8] ));
 sg13g2_dfrbp_1 _36073_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1411),
    .D(_02658_),
    .Q_N(_14562_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][9] ));
 sg13g2_dfrbp_1 _36074_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1286),
    .D(_02659_),
    .Q_N(_14561_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][10] ));
 sg13g2_dfrbp_1 _36075_ (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1282),
    .D(_02660_),
    .Q_N(_14560_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][11] ));
 sg13g2_dfrbp_1 _36076_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1278),
    .D(_02661_),
    .Q_N(_14559_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][12] ));
 sg13g2_dfrbp_1 _36077_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1274),
    .D(_02662_),
    .Q_N(_14558_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][13] ));
 sg13g2_dfrbp_1 _36078_ (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1270),
    .D(_02663_),
    .Q_N(_14557_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][14] ));
 sg13g2_dfrbp_1 _36079_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1266),
    .D(_02664_),
    .Q_N(_14556_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][15] ));
 sg13g2_dfrbp_1 _36080_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1262),
    .D(_02665_),
    .Q_N(_14555_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][16] ));
 sg13g2_dfrbp_1 _36081_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1258),
    .D(_02666_),
    .Q_N(_14554_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][17] ));
 sg13g2_dfrbp_1 _36082_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1254),
    .D(_02667_),
    .Q_N(_14553_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][18] ));
 sg13g2_dfrbp_1 _36083_ (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1250),
    .D(_02668_),
    .Q_N(_14552_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][19] ));
 sg13g2_dfrbp_1 _36084_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1246),
    .D(_02669_),
    .Q_N(_14551_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][20] ));
 sg13g2_dfrbp_1 _36085_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1242),
    .D(_02670_),
    .Q_N(_14550_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][21] ));
 sg13g2_dfrbp_1 _36086_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1238),
    .D(_02671_),
    .Q_N(_14549_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][22] ));
 sg13g2_dfrbp_1 _36087_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1234),
    .D(_02672_),
    .Q_N(_14548_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][23] ));
 sg13g2_dfrbp_1 _36088_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1230),
    .D(_02673_),
    .Q_N(_14547_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][24] ));
 sg13g2_dfrbp_1 _36089_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1226),
    .D(_02674_),
    .Q_N(_14546_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][25] ));
 sg13g2_dfrbp_1 _36090_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1222),
    .D(_02675_),
    .Q_N(_14545_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][26] ));
 sg13g2_dfrbp_1 _36091_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1218),
    .D(_02676_),
    .Q_N(_14544_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][27] ));
 sg13g2_dfrbp_1 _36092_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1214),
    .D(_02677_),
    .Q_N(_14543_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][28] ));
 sg13g2_dfrbp_1 _36093_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1210),
    .D(_02678_),
    .Q_N(_14542_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][29] ));
 sg13g2_dfrbp_1 _36094_ (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1206),
    .D(_02679_),
    .Q_N(_14541_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][30] ));
 sg13g2_dfrbp_1 _36095_ (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1202),
    .D(_02680_),
    .Q_N(_14540_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][31] ));
 sg13g2_dfrbp_1 _36096_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1198),
    .D(_02681_),
    .Q_N(_00209_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[0] ));
 sg13g2_dfrbp_1 _36097_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1194),
    .D(_02682_),
    .Q_N(_00205_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[1] ));
 sg13g2_dfrbp_1 _36098_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1190),
    .D(_02683_),
    .Q_N(_00201_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[2] ));
 sg13g2_dfrbp_1 _36099_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1186),
    .D(_02684_),
    .Q_N(_00237_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[3] ));
 sg13g2_dfrbp_1 _36100_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1182),
    .D(_02685_),
    .Q_N(_00197_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[4] ));
 sg13g2_dfrbp_1 _36101_ (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1178),
    .D(_02686_),
    .Q_N(_00193_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[5] ));
 sg13g2_dfrbp_1 _36102_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1174),
    .D(_02687_),
    .Q_N(_00187_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[6] ));
 sg13g2_dfrbp_1 _36103_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1170),
    .D(_02688_),
    .Q_N(_00235_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[7] ));
 sg13g2_dfrbp_1 _36104_ (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1166),
    .D(_02689_),
    .Q_N(_00211_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[8] ));
 sg13g2_dfrbp_1 _36105_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1098),
    .D(_02690_),
    .Q_N(_00207_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[9] ));
 sg13g2_dfrbp_1 _36106_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1094),
    .D(_02691_),
    .Q_N(_00203_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[10] ));
 sg13g2_dfrbp_1 _36107_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1082),
    .D(_02692_),
    .Q_N(_00234_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[11] ));
 sg13g2_dfrbp_1 _36108_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1078),
    .D(_02693_),
    .Q_N(_00199_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[12] ));
 sg13g2_dfrbp_1 _36109_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1074),
    .D(_02694_),
    .Q_N(_00195_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[13] ));
 sg13g2_dfrbp_1 _36110_ (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1070),
    .D(_02695_),
    .Q_N(_00191_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[14] ));
 sg13g2_dfrbp_1 _36111_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1066),
    .D(_02696_),
    .Q_N(_00233_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[15] ));
 sg13g2_dfrbp_1 _36112_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1062),
    .D(_02697_),
    .Q_N(_00232_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[16] ));
 sg13g2_dfrbp_1 _36113_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1058),
    .D(_02698_),
    .Q_N(_00231_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[17] ));
 sg13g2_dfrbp_1 _36114_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1054),
    .D(_02699_),
    .Q_N(_00230_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[18] ));
 sg13g2_dfrbp_1 _36115_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1050),
    .D(_02700_),
    .Q_N(_00229_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[19] ));
 sg13g2_dfrbp_1 _36116_ (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1046),
    .D(_02701_),
    .Q_N(_00228_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[20] ));
 sg13g2_dfrbp_1 _36117_ (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1042),
    .D(_02702_),
    .Q_N(_00227_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[21] ));
 sg13g2_dfrbp_1 _36118_ (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1038),
    .D(_02703_),
    .Q_N(_00226_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[22] ));
 sg13g2_dfrbp_1 _36119_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1034),
    .D(_02704_),
    .Q_N(_00225_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[23] ));
 sg13g2_dfrbp_1 _36120_ (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1030),
    .D(_02705_),
    .Q_N(_00224_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[24] ));
 sg13g2_dfrbp_1 _36121_ (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1026),
    .D(_02706_),
    .Q_N(_00223_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[25] ));
 sg13g2_dfrbp_1 _36122_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1022),
    .D(_02707_),
    .Q_N(_00222_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[26] ));
 sg13g2_dfrbp_1 _36123_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1018),
    .D(_02708_),
    .Q_N(_00221_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[27] ));
 sg13g2_dfrbp_1 _36124_ (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1014),
    .D(_02709_),
    .Q_N(_00220_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[28] ));
 sg13g2_dfrbp_1 _36125_ (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1010),
    .D(_02710_),
    .Q_N(_00219_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[29] ));
 sg13g2_dfrbp_1 _36126_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1006),
    .D(_02711_),
    .Q_N(_00218_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[30] ));
 sg13g2_dfrbp_1 _36127_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1002),
    .D(_02712_),
    .Q_N(_00217_),
    .Q(\soc_I.kianv_I.datapath_unit_I.A2[31] ));
 sg13g2_dfrbp_1 _36128_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net998),
    .D(_02713_),
    .Q_N(_14539_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][0] ));
 sg13g2_dfrbp_1 _36129_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net994),
    .D(_02714_),
    .Q_N(_14538_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][1] ));
 sg13g2_dfrbp_1 _36130_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net990),
    .D(_02715_),
    .Q_N(_14537_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][2] ));
 sg13g2_dfrbp_1 _36131_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net986),
    .D(_02716_),
    .Q_N(_14536_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][3] ));
 sg13g2_dfrbp_1 _36132_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net982),
    .D(_02717_),
    .Q_N(_14535_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][4] ));
 sg13g2_dfrbp_1 _36133_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net978),
    .D(_02718_),
    .Q_N(_14534_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][5] ));
 sg13g2_dfrbp_1 _36134_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net974),
    .D(_02719_),
    .Q_N(_14533_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][6] ));
 sg13g2_dfrbp_1 _36135_ (.CLK(clknet_leaf_304_clk),
    .RESET_B(net970),
    .D(_02720_),
    .Q_N(_14532_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][7] ));
 sg13g2_dfrbp_1 _36136_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net966),
    .D(_02721_),
    .Q_N(_14531_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][8] ));
 sg13g2_dfrbp_1 _36137_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net962),
    .D(_02722_),
    .Q_N(_14530_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][9] ));
 sg13g2_dfrbp_1 _36138_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net958),
    .D(_02723_),
    .Q_N(_14529_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][10] ));
 sg13g2_dfrbp_1 _36139_ (.CLK(clknet_leaf_315_clk),
    .RESET_B(net954),
    .D(_02724_),
    .Q_N(_14528_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][11] ));
 sg13g2_dfrbp_1 _36140_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net950),
    .D(_02725_),
    .Q_N(_14527_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][12] ));
 sg13g2_dfrbp_1 _36141_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net946),
    .D(_02726_),
    .Q_N(_14526_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][13] ));
 sg13g2_dfrbp_1 _36142_ (.CLK(clknet_leaf_299_clk),
    .RESET_B(net942),
    .D(_02727_),
    .Q_N(_14525_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][14] ));
 sg13g2_dfrbp_1 _36143_ (.CLK(clknet_leaf_310_clk),
    .RESET_B(net938),
    .D(_02728_),
    .Q_N(_14524_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][15] ));
 sg13g2_dfrbp_1 _36144_ (.CLK(clknet_leaf_316_clk),
    .RESET_B(net934),
    .D(_02729_),
    .Q_N(_14523_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][16] ));
 sg13g2_dfrbp_1 _36145_ (.CLK(clknet_leaf_311_clk),
    .RESET_B(net930),
    .D(net2898),
    .Q_N(_14522_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][17] ));
 sg13g2_dfrbp_1 _36146_ (.CLK(clknet_leaf_303_clk),
    .RESET_B(net926),
    .D(_02731_),
    .Q_N(_14521_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][18] ));
 sg13g2_dfrbp_1 _36147_ (.CLK(clknet_leaf_300_clk),
    .RESET_B(net922),
    .D(_02732_),
    .Q_N(_14520_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][19] ));
 sg13g2_dfrbp_1 _36148_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net918),
    .D(_02733_),
    .Q_N(_14519_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][20] ));
 sg13g2_dfrbp_1 _36149_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net914),
    .D(_02734_),
    .Q_N(_14518_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][21] ));
 sg13g2_dfrbp_1 _36150_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net910),
    .D(_02735_),
    .Q_N(_14517_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][22] ));
 sg13g2_dfrbp_1 _36151_ (.CLK(clknet_leaf_310_clk),
    .RESET_B(net906),
    .D(_02736_),
    .Q_N(_14516_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][23] ));
 sg13g2_dfrbp_1 _36152_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net902),
    .D(_02737_),
    .Q_N(_14515_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][24] ));
 sg13g2_dfrbp_1 _36153_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net898),
    .D(_02738_),
    .Q_N(_14514_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][25] ));
 sg13g2_dfrbp_1 _36154_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net894),
    .D(_02739_),
    .Q_N(_14513_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][26] ));
 sg13g2_dfrbp_1 _36155_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net890),
    .D(_02740_),
    .Q_N(_14512_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][27] ));
 sg13g2_dfrbp_1 _36156_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net886),
    .D(_02741_),
    .Q_N(_14511_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][28] ));
 sg13g2_dfrbp_1 _36157_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net882),
    .D(_02742_),
    .Q_N(_14510_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][29] ));
 sg13g2_dfrbp_1 _36158_ (.CLK(clknet_leaf_296_clk),
    .RESET_B(net878),
    .D(_02743_),
    .Q_N(_14509_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][30] ));
 sg13g2_dfrbp_1 _36159_ (.CLK(clknet_leaf_286_clk),
    .RESET_B(net874),
    .D(_02744_),
    .Q_N(_14508_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][31] ));
 sg13g2_dfrbp_1 _36160_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net870),
    .D(_02745_),
    .Q_N(_14507_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][0] ));
 sg13g2_dfrbp_1 _36161_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net866),
    .D(_02746_),
    .Q_N(_14506_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][1] ));
 sg13g2_dfrbp_1 _36162_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net862),
    .D(_02747_),
    .Q_N(_14505_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][2] ));
 sg13g2_dfrbp_1 _36163_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net858),
    .D(_02748_),
    .Q_N(_14504_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][3] ));
 sg13g2_dfrbp_1 _36164_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net854),
    .D(_02749_),
    .Q_N(_14503_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][4] ));
 sg13g2_dfrbp_1 _36165_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net850),
    .D(_02750_),
    .Q_N(_14502_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][5] ));
 sg13g2_dfrbp_1 _36166_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net846),
    .D(_02751_),
    .Q_N(_14501_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][6] ));
 sg13g2_dfrbp_1 _36167_ (.CLK(clknet_leaf_285_clk),
    .RESET_B(net778),
    .D(_02752_),
    .Q_N(_14500_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][7] ));
 sg13g2_dfrbp_1 _36168_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net774),
    .D(_02753_),
    .Q_N(_14499_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][8] ));
 sg13g2_dfrbp_1 _36169_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net770),
    .D(_02754_),
    .Q_N(_14498_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][9] ));
 sg13g2_dfrbp_1 _36170_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net733),
    .D(_02755_),
    .Q_N(_14497_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][10] ));
 sg13g2_dfrbp_1 _36171_ (.CLK(clknet_leaf_317_clk),
    .RESET_B(net2584),
    .D(_02756_),
    .Q_N(_14496_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][11] ));
 sg13g2_dfrbp_1 _36172_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2580),
    .D(_02757_),
    .Q_N(_14495_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][12] ));
 sg13g2_dfrbp_1 _36173_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2571),
    .D(_02758_),
    .Q_N(_14494_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][13] ));
 sg13g2_dfrbp_1 _36174_ (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2567),
    .D(_02759_),
    .Q_N(_14493_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][14] ));
 sg13g2_dfrbp_1 _36175_ (.CLK(clknet_leaf_310_clk),
    .RESET_B(net2563),
    .D(_02760_),
    .Q_N(_14492_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][15] ));
 sg13g2_dfrbp_1 _36176_ (.CLK(clknet_leaf_317_clk),
    .RESET_B(net2559),
    .D(_02761_),
    .Q_N(_14491_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][16] ));
 sg13g2_dfrbp_1 _36177_ (.CLK(clknet_leaf_311_clk),
    .RESET_B(net2555),
    .D(_02762_),
    .Q_N(_14490_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][17] ));
 sg13g2_dfrbp_1 _36178_ (.CLK(clknet_leaf_302_clk),
    .RESET_B(net2519),
    .D(_02763_),
    .Q_N(_14489_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][18] ));
 sg13g2_dfrbp_1 _36179_ (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2515),
    .D(_02764_),
    .Q_N(_14488_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][19] ));
 sg13g2_dfrbp_1 _36180_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2511),
    .D(_02765_),
    .Q_N(_14487_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][20] ));
 sg13g2_dfrbp_1 _36181_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2507),
    .D(_02766_),
    .Q_N(_14486_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][21] ));
 sg13g2_dfrbp_1 _36182_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2503),
    .D(_02767_),
    .Q_N(_14485_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][22] ));
 sg13g2_dfrbp_1 _36183_ (.CLK(clknet_leaf_311_clk),
    .RESET_B(net2499),
    .D(_02768_),
    .Q_N(_14484_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][23] ));
 sg13g2_dfrbp_1 _36184_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2495),
    .D(_02769_),
    .Q_N(_14483_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][24] ));
 sg13g2_dfrbp_1 _36185_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2491),
    .D(_02770_),
    .Q_N(_14482_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][25] ));
 sg13g2_dfrbp_1 _36186_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2487),
    .D(_02771_),
    .Q_N(_14481_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][26] ));
 sg13g2_dfrbp_1 _36187_ (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2483),
    .D(_02772_),
    .Q_N(_14480_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][27] ));
 sg13g2_dfrbp_1 _36188_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2479),
    .D(_02773_),
    .Q_N(_14479_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][28] ));
 sg13g2_dfrbp_1 _36189_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net2475),
    .D(_02774_),
    .Q_N(_14478_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][29] ));
 sg13g2_dfrbp_1 _36190_ (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2471),
    .D(_02775_),
    .Q_N(_14477_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][30] ));
 sg13g2_dfrbp_1 _36191_ (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2467),
    .D(_02776_),
    .Q_N(_14476_),
    .Q(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][31] ));
 sg13g2_dfrbp_1 _36192_ (.CLK(clknet_leaf_325_clk),
    .RESET_B(net2463),
    .D(_02777_),
    .Q_N(_14475_),
    .Q(_00000_));
 sg13g2_dfrbp_1 _36193_ (.CLK(clknet_leaf_325_clk),
    .RESET_B(net2459),
    .D(_02778_),
    .Q_N(_14474_),
    .Q(_00001_));
 sg13g2_dfrbp_1 _36194_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net2455),
    .D(_02779_),
    .Q_N(_14473_),
    .Q(_00002_));
 sg13g2_dfrbp_1 _36195_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net2451),
    .D(net3148),
    .Q_N(_14472_),
    .Q(_00003_));
 sg13g2_tiehi _35181__15 (.L_HI(net15));
 sg13g2_tiehi _35930__16 (.L_HI(net16));
 sg13g2_tiehi _35180__17 (.L_HI(net17));
 sg13g2_tiehi _35929__18 (.L_HI(net18));
 sg13g2_tiehi _35179__19 (.L_HI(net19));
 sg13g2_tiehi _35928__20 (.L_HI(net20));
 sg13g2_tiehi _35178__21 (.L_HI(net21));
 sg13g2_tiehi _35927__22 (.L_HI(net22));
 sg13g2_tiehi _35177__23 (.L_HI(net23));
 sg13g2_tiehi _35926__24 (.L_HI(net24));
 sg13g2_tiehi _35176__25 (.L_HI(net25));
 sg13g2_tiehi _35925__26 (.L_HI(net26));
 sg13g2_tiehi _35175__27 (.L_HI(net27));
 sg13g2_tiehi _35924__28 (.L_HI(net28));
 sg13g2_tiehi _35174__29 (.L_HI(net29));
 sg13g2_tiehi _35923__30 (.L_HI(net30));
 sg13g2_tiehi _35173__31 (.L_HI(net31));
 sg13g2_tiehi _35922__32 (.L_HI(net32));
 sg13g2_tiehi _35172__33 (.L_HI(net33));
 sg13g2_tiehi _35921__34 (.L_HI(net34));
 sg13g2_tiehi _35171__35 (.L_HI(net35));
 sg13g2_tiehi _35920__36 (.L_HI(net36));
 sg13g2_tiehi _35170__37 (.L_HI(net37));
 sg13g2_tiehi _35919__38 (.L_HI(net38));
 sg13g2_tiehi _35169__39 (.L_HI(net39));
 sg13g2_tiehi _35918__40 (.L_HI(net40));
 sg13g2_tiehi _35168__41 (.L_HI(net41));
 sg13g2_tiehi _35917__42 (.L_HI(net42));
 sg13g2_tiehi _35167__43 (.L_HI(net43));
 sg13g2_tiehi _35916__44 (.L_HI(net44));
 sg13g2_tiehi _35166__45 (.L_HI(net45));
 sg13g2_tiehi _35915__46 (.L_HI(net46));
 sg13g2_tiehi _35165__47 (.L_HI(net47));
 sg13g2_tiehi _35914__48 (.L_HI(net48));
 sg13g2_tiehi _35164__49 (.L_HI(net49));
 sg13g2_tiehi _35913__50 (.L_HI(net50));
 sg13g2_tiehi _35163__51 (.L_HI(net51));
 sg13g2_tiehi _35912__52 (.L_HI(net52));
 sg13g2_tiehi _35162__53 (.L_HI(net53));
 sg13g2_tiehi _35911__54 (.L_HI(net54));
 sg13g2_tiehi _35161__55 (.L_HI(net55));
 sg13g2_tiehi _35910__56 (.L_HI(net56));
 sg13g2_tiehi _35160__57 (.L_HI(net57));
 sg13g2_tiehi _35909__58 (.L_HI(net58));
 sg13g2_tiehi _35159__59 (.L_HI(net59));
 sg13g2_tiehi _35908__60 (.L_HI(net60));
 sg13g2_tiehi _35158__61 (.L_HI(net61));
 sg13g2_tiehi _35907__62 (.L_HI(net62));
 sg13g2_tiehi _35157__63 (.L_HI(net63));
 sg13g2_tiehi _35906__64 (.L_HI(net64));
 sg13g2_tiehi _35156__65 (.L_HI(net65));
 sg13g2_tiehi _35905__66 (.L_HI(net66));
 sg13g2_tiehi _35155__67 (.L_HI(net67));
 sg13g2_tiehi _35904__68 (.L_HI(net68));
 sg13g2_tiehi _35154__69 (.L_HI(net69));
 sg13g2_tiehi _35903__70 (.L_HI(net70));
 sg13g2_tiehi _35153__71 (.L_HI(net71));
 sg13g2_tiehi _35152__72 (.L_HI(net72));
 sg13g2_tiehi _35151__73 (.L_HI(net73));
 sg13g2_tiehi _35150__74 (.L_HI(net74));
 sg13g2_tiehi _35149__75 (.L_HI(net75));
 sg13g2_tiehi _35148__76 (.L_HI(net76));
 sg13g2_tiehi _35147__77 (.L_HI(net77));
 sg13g2_tiehi _35146__78 (.L_HI(net78));
 sg13g2_tiehi _35145__79 (.L_HI(net79));
 sg13g2_tiehi _35144__80 (.L_HI(net80));
 sg13g2_tiehi _35143__81 (.L_HI(net81));
 sg13g2_tiehi _35142__82 (.L_HI(net82));
 sg13g2_tiehi _35141__83 (.L_HI(net83));
 sg13g2_tiehi _35140__84 (.L_HI(net84));
 sg13g2_tiehi _35139__85 (.L_HI(net85));
 sg13g2_tiehi _35138__86 (.L_HI(net86));
 sg13g2_tiehi _35137__87 (.L_HI(net87));
 sg13g2_tiehi _35136__88 (.L_HI(net88));
 sg13g2_tiehi _35135__89 (.L_HI(net89));
 sg13g2_tiehi _35134__90 (.L_HI(net90));
 sg13g2_tiehi _35133__91 (.L_HI(net91));
 sg13g2_tiehi _35132__92 (.L_HI(net92));
 sg13g2_tiehi _35131__93 (.L_HI(net93));
 sg13g2_tiehi _35130__94 (.L_HI(net94));
 sg13g2_tiehi _35129__95 (.L_HI(net95));
 sg13g2_tiehi _35128__96 (.L_HI(net96));
 sg13g2_tiehi _35127__97 (.L_HI(net97));
 sg13g2_tiehi _35126__98 (.L_HI(net98));
 sg13g2_tiehi _35125__99 (.L_HI(net99));
 sg13g2_tiehi _35124__100 (.L_HI(net100));
 sg13g2_tiehi _35123__101 (.L_HI(net101));
 sg13g2_tiehi _35122__102 (.L_HI(net102));
 sg13g2_tiehi _35121__103 (.L_HI(net103));
 sg13g2_tiehi _35902__104 (.L_HI(net104));
 sg13g2_tiehi _35120__105 (.L_HI(net105));
 sg13g2_tiehi _35901__106 (.L_HI(net106));
 sg13g2_tiehi _35119__107 (.L_HI(net107));
 sg13g2_tiehi _35900__108 (.L_HI(net108));
 sg13g2_tiehi _35118__109 (.L_HI(net109));
 sg13g2_tiehi _35899__110 (.L_HI(net110));
 sg13g2_tiehi _35117__111 (.L_HI(net111));
 sg13g2_tiehi _35898__112 (.L_HI(net112));
 sg13g2_tiehi _35116__113 (.L_HI(net113));
 sg13g2_tiehi _35897__114 (.L_HI(net114));
 sg13g2_tiehi _35115__115 (.L_HI(net115));
 sg13g2_tiehi _35896__116 (.L_HI(net116));
 sg13g2_tiehi _35114__117 (.L_HI(net117));
 sg13g2_tiehi _35895__118 (.L_HI(net118));
 sg13g2_tiehi _35113__119 (.L_HI(net119));
 sg13g2_tiehi _35112__120 (.L_HI(net120));
 sg13g2_tiehi _35894__121 (.L_HI(net121));
 sg13g2_tiehi _35111__122 (.L_HI(net122));
 sg13g2_tiehi _35893__123 (.L_HI(net123));
 sg13g2_tiehi _35110__124 (.L_HI(net124));
 sg13g2_tiehi _35892__125 (.L_HI(net125));
 sg13g2_tiehi _35109__126 (.L_HI(net126));
 sg13g2_tiehi _35891__127 (.L_HI(net127));
 sg13g2_tiehi _35108__128 (.L_HI(net128));
 sg13g2_tiehi _35890__129 (.L_HI(net129));
 sg13g2_tiehi _35107__130 (.L_HI(net130));
 sg13g2_tiehi _35889__131 (.L_HI(net131));
 sg13g2_tiehi _35106__132 (.L_HI(net132));
 sg13g2_tiehi _35888__133 (.L_HI(net133));
 sg13g2_tiehi _35105__134 (.L_HI(net134));
 sg13g2_tiehi _35887__135 (.L_HI(net135));
 sg13g2_tiehi _35104__136 (.L_HI(net136));
 sg13g2_tiehi _35886__137 (.L_HI(net137));
 sg13g2_tiehi _35103__138 (.L_HI(net138));
 sg13g2_tiehi _35885__139 (.L_HI(net139));
 sg13g2_tiehi _35102__140 (.L_HI(net140));
 sg13g2_tiehi _35884__141 (.L_HI(net141));
 sg13g2_tiehi _35101__142 (.L_HI(net142));
 sg13g2_tiehi _35883__143 (.L_HI(net143));
 sg13g2_tiehi _35100__144 (.L_HI(net144));
 sg13g2_tiehi _35882__145 (.L_HI(net145));
 sg13g2_tiehi _35099__146 (.L_HI(net146));
 sg13g2_tiehi _35881__147 (.L_HI(net147));
 sg13g2_tiehi _35098__148 (.L_HI(net148));
 sg13g2_tiehi _35880__149 (.L_HI(net149));
 sg13g2_tiehi _35097__150 (.L_HI(net150));
 sg13g2_tiehi _35879__151 (.L_HI(net151));
 sg13g2_tiehi _35096__152 (.L_HI(net152));
 sg13g2_tiehi _35878__153 (.L_HI(net153));
 sg13g2_tiehi _35095__154 (.L_HI(net154));
 sg13g2_tiehi _35877__155 (.L_HI(net155));
 sg13g2_tiehi _35094__156 (.L_HI(net156));
 sg13g2_tiehi _35876__157 (.L_HI(net157));
 sg13g2_tiehi _35093__158 (.L_HI(net158));
 sg13g2_tiehi _35875__159 (.L_HI(net159));
 sg13g2_tiehi _35092__160 (.L_HI(net160));
 sg13g2_tiehi _35874__161 (.L_HI(net161));
 sg13g2_tiehi _35091__162 (.L_HI(net162));
 sg13g2_tiehi _35873__163 (.L_HI(net163));
 sg13g2_tiehi _35090__164 (.L_HI(net164));
 sg13g2_tiehi _35872__165 (.L_HI(net165));
 sg13g2_tiehi _35089__166 (.L_HI(net166));
 sg13g2_tiehi _35871__167 (.L_HI(net167));
 sg13g2_tiehi _35088__168 (.L_HI(net168));
 sg13g2_tiehi _35870__169 (.L_HI(net169));
 sg13g2_tiehi _35087__170 (.L_HI(net170));
 sg13g2_tiehi _35869__171 (.L_HI(net171));
 sg13g2_tiehi _35086__172 (.L_HI(net172));
 sg13g2_tiehi _35868__173 (.L_HI(net173));
 sg13g2_tiehi _35085__174 (.L_HI(net174));
 sg13g2_tiehi _35867__175 (.L_HI(net175));
 sg13g2_tiehi _35084__176 (.L_HI(net176));
 sg13g2_tiehi _35866__177 (.L_HI(net177));
 sg13g2_tiehi _35083__178 (.L_HI(net178));
 sg13g2_tiehi _35865__179 (.L_HI(net179));
 sg13g2_tiehi _35082__180 (.L_HI(net180));
 sg13g2_tiehi _35864__181 (.L_HI(net181));
 sg13g2_tiehi _35081__182 (.L_HI(net182));
 sg13g2_tiehi _35863__183 (.L_HI(net183));
 sg13g2_tiehi _35080__184 (.L_HI(net184));
 sg13g2_tiehi _35862__185 (.L_HI(net185));
 sg13g2_tiehi _35079__186 (.L_HI(net186));
 sg13g2_tiehi _35861__187 (.L_HI(net187));
 sg13g2_tiehi _35078__188 (.L_HI(net188));
 sg13g2_tiehi _35860__189 (.L_HI(net189));
 sg13g2_tiehi _35077__190 (.L_HI(net190));
 sg13g2_tiehi _35859__191 (.L_HI(net191));
 sg13g2_tiehi _35076__192 (.L_HI(net192));
 sg13g2_tiehi _35858__193 (.L_HI(net193));
 sg13g2_tiehi _35075__194 (.L_HI(net194));
 sg13g2_tiehi _35857__195 (.L_HI(net195));
 sg13g2_tiehi _35074__196 (.L_HI(net196));
 sg13g2_tiehi _35856__197 (.L_HI(net197));
 sg13g2_tiehi _35073__198 (.L_HI(net198));
 sg13g2_tiehi _35855__199 (.L_HI(net199));
 sg13g2_tiehi _35072__200 (.L_HI(net200));
 sg13g2_tiehi _35854__201 (.L_HI(net201));
 sg13g2_tiehi _35071__202 (.L_HI(net202));
 sg13g2_tiehi _35853__203 (.L_HI(net203));
 sg13g2_tiehi _35070__204 (.L_HI(net204));
 sg13g2_tiehi _35852__205 (.L_HI(net205));
 sg13g2_tiehi _35069__206 (.L_HI(net206));
 sg13g2_tiehi _35851__207 (.L_HI(net207));
 sg13g2_tiehi _35068__208 (.L_HI(net208));
 sg13g2_tiehi _35850__209 (.L_HI(net209));
 sg13g2_tiehi _35067__210 (.L_HI(net210));
 sg13g2_tiehi _35849__211 (.L_HI(net211));
 sg13g2_tiehi _35066__212 (.L_HI(net212));
 sg13g2_tiehi _35848__213 (.L_HI(net213));
 sg13g2_tiehi _35065__214 (.L_HI(net214));
 sg13g2_tiehi _35847__215 (.L_HI(net215));
 sg13g2_tiehi _35064__216 (.L_HI(net216));
 sg13g2_tiehi _35846__217 (.L_HI(net217));
 sg13g2_tiehi _35063__218 (.L_HI(net218));
 sg13g2_tiehi _35845__219 (.L_HI(net219));
 sg13g2_tiehi _35062__220 (.L_HI(net220));
 sg13g2_tiehi _35844__221 (.L_HI(net221));
 sg13g2_tiehi _35061__222 (.L_HI(net222));
 sg13g2_tiehi _35843__223 (.L_HI(net223));
 sg13g2_tiehi _35060__224 (.L_HI(net224));
 sg13g2_tiehi _35842__225 (.L_HI(net225));
 sg13g2_tiehi _35059__226 (.L_HI(net226));
 sg13g2_tiehi _35841__227 (.L_HI(net227));
 sg13g2_tiehi _35058__228 (.L_HI(net228));
 sg13g2_tiehi _35840__229 (.L_HI(net229));
 sg13g2_tiehi _35057__230 (.L_HI(net230));
 sg13g2_tiehi _35839__231 (.L_HI(net231));
 sg13g2_tiehi _35056__232 (.L_HI(net232));
 sg13g2_tiehi _35838__233 (.L_HI(net233));
 sg13g2_tiehi _35055__234 (.L_HI(net234));
 sg13g2_tiehi _35837__235 (.L_HI(net235));
 sg13g2_tiehi _35054__236 (.L_HI(net236));
 sg13g2_tiehi _35836__237 (.L_HI(net237));
 sg13g2_tiehi _35053__238 (.L_HI(net238));
 sg13g2_tiehi _35835__239 (.L_HI(net239));
 sg13g2_tiehi _35052__240 (.L_HI(net240));
 sg13g2_tiehi _35834__241 (.L_HI(net241));
 sg13g2_tiehi _35051__242 (.L_HI(net242));
 sg13g2_tiehi _35833__243 (.L_HI(net243));
 sg13g2_tiehi _35050__244 (.L_HI(net244));
 sg13g2_tiehi _35832__245 (.L_HI(net245));
 sg13g2_tiehi _35049__246 (.L_HI(net246));
 sg13g2_tiehi _35831__247 (.L_HI(net247));
 sg13g2_tiehi _35048__248 (.L_HI(net248));
 sg13g2_tiehi _35830__249 (.L_HI(net249));
 sg13g2_tiehi _35047__250 (.L_HI(net250));
 sg13g2_tiehi _35829__251 (.L_HI(net251));
 sg13g2_tiehi _35046__252 (.L_HI(net252));
 sg13g2_tiehi _35828__253 (.L_HI(net253));
 sg13g2_tiehi _35045__254 (.L_HI(net254));
 sg13g2_tiehi _35827__255 (.L_HI(net255));
 sg13g2_tiehi _35044__256 (.L_HI(net256));
 sg13g2_tiehi _35826__257 (.L_HI(net257));
 sg13g2_tiehi _35043__258 (.L_HI(net258));
 sg13g2_tiehi _35825__259 (.L_HI(net259));
 sg13g2_tiehi _35042__260 (.L_HI(net260));
 sg13g2_tiehi _35824__261 (.L_HI(net261));
 sg13g2_tiehi _35041__262 (.L_HI(net262));
 sg13g2_tiehi _35823__263 (.L_HI(net263));
 sg13g2_tiehi _35040__264 (.L_HI(net264));
 sg13g2_tiehi _35039__265 (.L_HI(net265));
 sg13g2_tiehi _35038__266 (.L_HI(net266));
 sg13g2_tiehi _35037__267 (.L_HI(net267));
 sg13g2_tiehi _35036__268 (.L_HI(net268));
 sg13g2_tiehi _35822__269 (.L_HI(net269));
 sg13g2_tiehi _35035__270 (.L_HI(net270));
 sg13g2_tiehi _35821__271 (.L_HI(net271));
 sg13g2_tiehi _35034__272 (.L_HI(net272));
 sg13g2_tiehi _35820__273 (.L_HI(net273));
 sg13g2_tiehi _35033__274 (.L_HI(net274));
 sg13g2_tiehi _35819__275 (.L_HI(net275));
 sg13g2_tiehi _35032__276 (.L_HI(net276));
 sg13g2_tiehi _35818__277 (.L_HI(net277));
 sg13g2_tiehi _35031__278 (.L_HI(net278));
 sg13g2_tiehi _35817__279 (.L_HI(net279));
 sg13g2_tiehi _35030__280 (.L_HI(net280));
 sg13g2_tiehi _35816__281 (.L_HI(net281));
 sg13g2_tiehi _35029__282 (.L_HI(net282));
 sg13g2_tiehi _35815__283 (.L_HI(net283));
 sg13g2_tiehi _35028__284 (.L_HI(net284));
 sg13g2_tiehi _35814__285 (.L_HI(net285));
 sg13g2_tiehi _35027__286 (.L_HI(net286));
 sg13g2_tiehi _35026__287 (.L_HI(net287));
 sg13g2_tiehi _35025__288 (.L_HI(net288));
 sg13g2_tiehi _35024__289 (.L_HI(net289));
 sg13g2_tiehi _35023__290 (.L_HI(net290));
 sg13g2_tiehi _35022__291 (.L_HI(net291));
 sg13g2_tiehi _35021__292 (.L_HI(net292));
 sg13g2_tiehi _35020__293 (.L_HI(net293));
 sg13g2_tiehi _35019__294 (.L_HI(net294));
 sg13g2_tiehi _35018__295 (.L_HI(net295));
 sg13g2_tiehi _35017__296 (.L_HI(net296));
 sg13g2_tiehi _35016__297 (.L_HI(net297));
 sg13g2_tiehi _35015__298 (.L_HI(net298));
 sg13g2_tiehi _35014__299 (.L_HI(net299));
 sg13g2_tiehi _35013__300 (.L_HI(net300));
 sg13g2_tiehi _35012__301 (.L_HI(net301));
 sg13g2_tiehi _35011__302 (.L_HI(net302));
 sg13g2_tiehi _35010__303 (.L_HI(net303));
 sg13g2_tiehi _35009__304 (.L_HI(net304));
 sg13g2_tiehi _35008__305 (.L_HI(net305));
 sg13g2_tiehi _35005__306 (.L_HI(net306));
 sg13g2_tiehi _34908__307 (.L_HI(net307));
 sg13g2_tiehi _34907__308 (.L_HI(net308));
 sg13g2_tiehi _34906__309 (.L_HI(net309));
 sg13g2_tiehi _34905__310 (.L_HI(net310));
 sg13g2_tiehi _34904__311 (.L_HI(net311));
 sg13g2_tiehi _34903__312 (.L_HI(net312));
 sg13g2_tiehi _34902__313 (.L_HI(net313));
 sg13g2_tiehi _34901__314 (.L_HI(net314));
 sg13g2_tiehi _34900__315 (.L_HI(net315));
 sg13g2_tiehi _34899__316 (.L_HI(net316));
 sg13g2_tiehi _34898__317 (.L_HI(net317));
 sg13g2_tiehi _34897__318 (.L_HI(net318));
 sg13g2_tiehi _34896__319 (.L_HI(net319));
 sg13g2_tiehi _34895__320 (.L_HI(net320));
 sg13g2_tiehi _34894__321 (.L_HI(net321));
 sg13g2_tiehi _34893__322 (.L_HI(net322));
 sg13g2_tiehi _34892__323 (.L_HI(net323));
 sg13g2_tiehi _34891__324 (.L_HI(net324));
 sg13g2_tiehi _34890__325 (.L_HI(net325));
 sg13g2_tiehi _34889__326 (.L_HI(net326));
 sg13g2_tiehi _34888__327 (.L_HI(net327));
 sg13g2_tiehi _34887__328 (.L_HI(net328));
 sg13g2_tiehi _34886__329 (.L_HI(net329));
 sg13g2_tiehi _34885__330 (.L_HI(net330));
 sg13g2_tiehi _34884__331 (.L_HI(net331));
 sg13g2_tiehi _34883__332 (.L_HI(net332));
 sg13g2_tiehi _34882__333 (.L_HI(net333));
 sg13g2_tiehi _34881__334 (.L_HI(net334));
 sg13g2_tiehi _34880__335 (.L_HI(net335));
 sg13g2_tiehi _34879__336 (.L_HI(net336));
 sg13g2_tiehi _34878__337 (.L_HI(net337));
 sg13g2_tiehi _35813__338 (.L_HI(net338));
 sg13g2_tiehi _34877__339 (.L_HI(net339));
 sg13g2_tiehi _35812__340 (.L_HI(net340));
 sg13g2_tiehi _34876__341 (.L_HI(net341));
 sg13g2_tiehi _35811__342 (.L_HI(net342));
 sg13g2_tiehi _34875__343 (.L_HI(net343));
 sg13g2_tiehi _35810__344 (.L_HI(net344));
 sg13g2_tiehi _34874__345 (.L_HI(net345));
 sg13g2_tiehi _35809__346 (.L_HI(net346));
 sg13g2_tiehi _34873__347 (.L_HI(net347));
 sg13g2_tiehi _35808__348 (.L_HI(net348));
 sg13g2_tiehi _34872__349 (.L_HI(net349));
 sg13g2_tiehi _35807__350 (.L_HI(net350));
 sg13g2_tiehi _34871__351 (.L_HI(net351));
 sg13g2_tiehi _35806__352 (.L_HI(net352));
 sg13g2_tiehi _34870__353 (.L_HI(net353));
 sg13g2_tiehi _35805__354 (.L_HI(net354));
 sg13g2_tiehi _34869__355 (.L_HI(net355));
 sg13g2_tiehi _35804__356 (.L_HI(net356));
 sg13g2_tiehi _34868__357 (.L_HI(net357));
 sg13g2_tiehi _35803__358 (.L_HI(net358));
 sg13g2_tiehi _34867__359 (.L_HI(net359));
 sg13g2_tiehi _35802__360 (.L_HI(net360));
 sg13g2_tiehi _34866__361 (.L_HI(net361));
 sg13g2_tiehi _35801__362 (.L_HI(net362));
 sg13g2_tiehi _34865__363 (.L_HI(net363));
 sg13g2_tiehi _35800__364 (.L_HI(net364));
 sg13g2_tiehi _34864__365 (.L_HI(net365));
 sg13g2_tiehi _35799__366 (.L_HI(net366));
 sg13g2_tiehi _34863__367 (.L_HI(net367));
 sg13g2_tiehi _35798__368 (.L_HI(net368));
 sg13g2_tiehi _34862__369 (.L_HI(net369));
 sg13g2_tiehi _35797__370 (.L_HI(net370));
 sg13g2_tiehi _34861__371 (.L_HI(net371));
 sg13g2_tiehi _35796__372 (.L_HI(net372));
 sg13g2_tiehi _34860__373 (.L_HI(net373));
 sg13g2_tiehi _35795__374 (.L_HI(net374));
 sg13g2_tiehi _34859__375 (.L_HI(net375));
 sg13g2_tiehi _35794__376 (.L_HI(net376));
 sg13g2_tiehi _34858__377 (.L_HI(net377));
 sg13g2_tiehi _35793__378 (.L_HI(net378));
 sg13g2_tiehi _34857__379 (.L_HI(net379));
 sg13g2_tiehi _35792__380 (.L_HI(net380));
 sg13g2_tiehi _34856__381 (.L_HI(net381));
 sg13g2_tiehi _35791__382 (.L_HI(net382));
 sg13g2_tiehi _34855__383 (.L_HI(net383));
 sg13g2_tiehi _35790__384 (.L_HI(net384));
 sg13g2_tiehi _34854__385 (.L_HI(net385));
 sg13g2_tiehi _35789__386 (.L_HI(net386));
 sg13g2_tiehi _34853__387 (.L_HI(net387));
 sg13g2_tiehi _35788__388 (.L_HI(net388));
 sg13g2_tiehi _34852__389 (.L_HI(net389));
 sg13g2_tiehi _35787__390 (.L_HI(net390));
 sg13g2_tiehi _34851__391 (.L_HI(net391));
 sg13g2_tiehi _35786__392 (.L_HI(net392));
 sg13g2_tiehi _34850__393 (.L_HI(net393));
 sg13g2_tiehi _35785__394 (.L_HI(net394));
 sg13g2_tiehi _34849__395 (.L_HI(net395));
 sg13g2_tiehi _35784__396 (.L_HI(net396));
 sg13g2_tiehi _34848__397 (.L_HI(net397));
 sg13g2_tiehi _35783__398 (.L_HI(net398));
 sg13g2_tiehi _34847__399 (.L_HI(net399));
 sg13g2_tiehi _35782__400 (.L_HI(net400));
 sg13g2_tiehi _34846__401 (.L_HI(net401));
 sg13g2_tiehi _35781__402 (.L_HI(net402));
 sg13g2_tiehi _34845__403 (.L_HI(net403));
 sg13g2_tiehi _35780__404 (.L_HI(net404));
 sg13g2_tiehi _34844__405 (.L_HI(net405));
 sg13g2_tiehi _35779__406 (.L_HI(net406));
 sg13g2_tiehi _34843__407 (.L_HI(net407));
 sg13g2_tiehi _35778__408 (.L_HI(net408));
 sg13g2_tiehi _34842__409 (.L_HI(net409));
 sg13g2_tiehi _35777__410 (.L_HI(net410));
 sg13g2_tiehi _34841__411 (.L_HI(net411));
 sg13g2_tiehi _35776__412 (.L_HI(net412));
 sg13g2_tiehi _34840__413 (.L_HI(net413));
 sg13g2_tiehi _35775__414 (.L_HI(net414));
 sg13g2_tiehi _34839__415 (.L_HI(net415));
 sg13g2_tiehi _35774__416 (.L_HI(net416));
 sg13g2_tiehi _34838__417 (.L_HI(net417));
 sg13g2_tiehi _35773__418 (.L_HI(net418));
 sg13g2_tiehi _34837__419 (.L_HI(net419));
 sg13g2_tiehi _35772__420 (.L_HI(net420));
 sg13g2_tiehi _34836__421 (.L_HI(net421));
 sg13g2_tiehi _35771__422 (.L_HI(net422));
 sg13g2_tiehi _34835__423 (.L_HI(net423));
 sg13g2_tiehi _35770__424 (.L_HI(net424));
 sg13g2_tiehi _34834__425 (.L_HI(net425));
 sg13g2_tiehi _35769__426 (.L_HI(net426));
 sg13g2_tiehi _34833__427 (.L_HI(net427));
 sg13g2_tiehi _35768__428 (.L_HI(net428));
 sg13g2_tiehi _34832__429 (.L_HI(net429));
 sg13g2_tiehi _35767__430 (.L_HI(net430));
 sg13g2_tiehi _34831__431 (.L_HI(net431));
 sg13g2_tiehi _35766__432 (.L_HI(net432));
 sg13g2_tiehi _34830__433 (.L_HI(net433));
 sg13g2_tiehi _35765__434 (.L_HI(net434));
 sg13g2_tiehi _34829__435 (.L_HI(net435));
 sg13g2_tiehi _35764__436 (.L_HI(net436));
 sg13g2_tiehi _34828__437 (.L_HI(net437));
 sg13g2_tiehi _35763__438 (.L_HI(net438));
 sg13g2_tiehi _34827__439 (.L_HI(net439));
 sg13g2_tiehi _35762__440 (.L_HI(net440));
 sg13g2_tiehi _34826__441 (.L_HI(net441));
 sg13g2_tiehi _35761__442 (.L_HI(net442));
 sg13g2_tiehi _34825__443 (.L_HI(net443));
 sg13g2_tiehi _35760__444 (.L_HI(net444));
 sg13g2_tiehi _34824__445 (.L_HI(net445));
 sg13g2_tiehi _35759__446 (.L_HI(net446));
 sg13g2_tiehi _34823__447 (.L_HI(net447));
 sg13g2_tiehi _35758__448 (.L_HI(net448));
 sg13g2_tiehi _34822__449 (.L_HI(net449));
 sg13g2_tiehi _35757__450 (.L_HI(net450));
 sg13g2_tiehi _34821__451 (.L_HI(net451));
 sg13g2_tiehi _35756__452 (.L_HI(net452));
 sg13g2_tiehi _34820__453 (.L_HI(net453));
 sg13g2_tiehi _35755__454 (.L_HI(net454));
 sg13g2_tiehi _34819__455 (.L_HI(net455));
 sg13g2_tiehi _35754__456 (.L_HI(net456));
 sg13g2_tiehi _34818__457 (.L_HI(net457));
 sg13g2_tiehi _35753__458 (.L_HI(net458));
 sg13g2_tiehi _34817__459 (.L_HI(net459));
 sg13g2_tiehi _35752__460 (.L_HI(net460));
 sg13g2_tiehi _34816__461 (.L_HI(net461));
 sg13g2_tiehi _35751__462 (.L_HI(net462));
 sg13g2_tiehi _34815__463 (.L_HI(net463));
 sg13g2_tiehi _35750__464 (.L_HI(net464));
 sg13g2_tiehi _34814__465 (.L_HI(net465));
 sg13g2_tiehi _35749__466 (.L_HI(net466));
 sg13g2_tiehi _34813__467 (.L_HI(net467));
 sg13g2_tiehi _35748__468 (.L_HI(net468));
 sg13g2_tiehi _34812__469 (.L_HI(net469));
 sg13g2_tiehi _35747__470 (.L_HI(net470));
 sg13g2_tiehi _34811__471 (.L_HI(net471));
 sg13g2_tiehi _35746__472 (.L_HI(net472));
 sg13g2_tiehi _34810__473 (.L_HI(net473));
 sg13g2_tiehi _35745__474 (.L_HI(net474));
 sg13g2_tiehi _34809__475 (.L_HI(net475));
 sg13g2_tiehi _35744__476 (.L_HI(net476));
 sg13g2_tiehi _34808__477 (.L_HI(net477));
 sg13g2_tiehi _35743__478 (.L_HI(net478));
 sg13g2_tiehi _34807__479 (.L_HI(net479));
 sg13g2_tiehi _35742__480 (.L_HI(net480));
 sg13g2_tiehi _34806__481 (.L_HI(net481));
 sg13g2_tiehi _35741__482 (.L_HI(net482));
 sg13g2_tiehi _34805__483 (.L_HI(net483));
 sg13g2_tiehi _35740__484 (.L_HI(net484));
 sg13g2_tiehi _34804__485 (.L_HI(net485));
 sg13g2_tiehi _35739__486 (.L_HI(net486));
 sg13g2_tiehi _34803__487 (.L_HI(net487));
 sg13g2_tiehi _35738__488 (.L_HI(net488));
 sg13g2_tiehi _34802__489 (.L_HI(net489));
 sg13g2_tiehi _35737__490 (.L_HI(net490));
 sg13g2_tiehi _34801__491 (.L_HI(net491));
 sg13g2_tiehi _35736__492 (.L_HI(net492));
 sg13g2_tiehi _34800__493 (.L_HI(net493));
 sg13g2_tiehi _35735__494 (.L_HI(net494));
 sg13g2_tiehi _34799__495 (.L_HI(net495));
 sg13g2_tiehi _35734__496 (.L_HI(net496));
 sg13g2_tiehi _34798__497 (.L_HI(net497));
 sg13g2_tiehi _35733__498 (.L_HI(net498));
 sg13g2_tiehi _34797__499 (.L_HI(net499));
 sg13g2_tiehi _35732__500 (.L_HI(net500));
 sg13g2_tiehi _34796__501 (.L_HI(net501));
 sg13g2_tiehi _35731__502 (.L_HI(net502));
 sg13g2_tiehi _34795__503 (.L_HI(net503));
 sg13g2_tiehi _35730__504 (.L_HI(net504));
 sg13g2_tiehi _34794__505 (.L_HI(net505));
 sg13g2_tiehi _35729__506 (.L_HI(net506));
 sg13g2_tiehi _34793__507 (.L_HI(net507));
 sg13g2_tiehi _35728__508 (.L_HI(net508));
 sg13g2_tiehi _34792__509 (.L_HI(net509));
 sg13g2_tiehi _35727__510 (.L_HI(net510));
 sg13g2_tiehi _34791__511 (.L_HI(net511));
 sg13g2_tiehi _35726__512 (.L_HI(net512));
 sg13g2_tiehi _34790__513 (.L_HI(net513));
 sg13g2_tiehi _35725__514 (.L_HI(net514));
 sg13g2_tiehi _34789__515 (.L_HI(net515));
 sg13g2_tiehi _35724__516 (.L_HI(net516));
 sg13g2_tiehi _34788__517 (.L_HI(net517));
 sg13g2_tiehi _35723__518 (.L_HI(net518));
 sg13g2_tiehi _34787__519 (.L_HI(net519));
 sg13g2_tiehi _35722__520 (.L_HI(net520));
 sg13g2_tiehi _34786__521 (.L_HI(net521));
 sg13g2_tiehi _35721__522 (.L_HI(net522));
 sg13g2_tiehi _34785__523 (.L_HI(net523));
 sg13g2_tiehi _35720__524 (.L_HI(net524));
 sg13g2_tiehi _34784__525 (.L_HI(net525));
 sg13g2_tiehi _35719__526 (.L_HI(net526));
 sg13g2_tiehi _34783__527 (.L_HI(net527));
 sg13g2_tiehi _35718__528 (.L_HI(net528));
 sg13g2_tiehi _34782__529 (.L_HI(net529));
 sg13g2_tiehi _35717__530 (.L_HI(net530));
 sg13g2_tiehi _34781__531 (.L_HI(net531));
 sg13g2_tiehi _35716__532 (.L_HI(net532));
 sg13g2_tiehi _34780__533 (.L_HI(net533));
 sg13g2_tiehi _35715__534 (.L_HI(net534));
 sg13g2_tiehi _34779__535 (.L_HI(net535));
 sg13g2_tiehi _35714__536 (.L_HI(net536));
 sg13g2_tiehi _34778__537 (.L_HI(net537));
 sg13g2_tiehi _35713__538 (.L_HI(net538));
 sg13g2_tiehi _34777__539 (.L_HI(net539));
 sg13g2_tiehi _35712__540 (.L_HI(net540));
 sg13g2_tiehi _34776__541 (.L_HI(net541));
 sg13g2_tiehi _35711__542 (.L_HI(net542));
 sg13g2_tiehi _34775__543 (.L_HI(net543));
 sg13g2_tiehi _35710__544 (.L_HI(net544));
 sg13g2_tiehi _34774__545 (.L_HI(net545));
 sg13g2_tiehi _35709__546 (.L_HI(net546));
 sg13g2_tiehi _34773__547 (.L_HI(net547));
 sg13g2_tiehi _35708__548 (.L_HI(net548));
 sg13g2_tiehi _34772__549 (.L_HI(net549));
 sg13g2_tiehi _35707__550 (.L_HI(net550));
 sg13g2_tiehi _34771__551 (.L_HI(net551));
 sg13g2_tiehi _35706__552 (.L_HI(net552));
 sg13g2_tiehi _34770__553 (.L_HI(net553));
 sg13g2_tiehi _35705__554 (.L_HI(net554));
 sg13g2_tiehi _34769__555 (.L_HI(net555));
 sg13g2_tiehi _35704__556 (.L_HI(net556));
 sg13g2_tiehi _34768__557 (.L_HI(net557));
 sg13g2_tiehi _35703__558 (.L_HI(net558));
 sg13g2_tiehi _34767__559 (.L_HI(net559));
 sg13g2_tiehi _35702__560 (.L_HI(net560));
 sg13g2_tiehi _34766__561 (.L_HI(net561));
 sg13g2_tiehi _35701__562 (.L_HI(net562));
 sg13g2_tiehi _34765__563 (.L_HI(net563));
 sg13g2_tiehi _35700__564 (.L_HI(net564));
 sg13g2_tiehi _34764__565 (.L_HI(net565));
 sg13g2_tiehi _35699__566 (.L_HI(net566));
 sg13g2_tiehi _34763__567 (.L_HI(net567));
 sg13g2_tiehi _35698__568 (.L_HI(net568));
 sg13g2_tiehi _34762__569 (.L_HI(net569));
 sg13g2_tiehi _35697__570 (.L_HI(net570));
 sg13g2_tiehi _34761__571 (.L_HI(net571));
 sg13g2_tiehi _35696__572 (.L_HI(net572));
 sg13g2_tiehi _34760__573 (.L_HI(net573));
 sg13g2_tiehi _35695__574 (.L_HI(net574));
 sg13g2_tiehi _34759__575 (.L_HI(net575));
 sg13g2_tiehi _35694__576 (.L_HI(net576));
 sg13g2_tiehi _34758__577 (.L_HI(net577));
 sg13g2_tiehi _35693__578 (.L_HI(net578));
 sg13g2_tiehi _34757__579 (.L_HI(net579));
 sg13g2_tiehi _35692__580 (.L_HI(net580));
 sg13g2_tiehi _34756__581 (.L_HI(net581));
 sg13g2_tiehi _35691__582 (.L_HI(net582));
 sg13g2_tiehi _34755__583 (.L_HI(net583));
 sg13g2_tiehi _35690__584 (.L_HI(net584));
 sg13g2_tiehi _34754__585 (.L_HI(net585));
 sg13g2_tiehi _35689__586 (.L_HI(net586));
 sg13g2_tiehi _34753__587 (.L_HI(net587));
 sg13g2_tiehi _35688__588 (.L_HI(net588));
 sg13g2_tiehi _34752__589 (.L_HI(net589));
 sg13g2_tiehi _35687__590 (.L_HI(net590));
 sg13g2_tiehi _34751__591 (.L_HI(net591));
 sg13g2_tiehi _35686__592 (.L_HI(net592));
 sg13g2_tiehi _34750__593 (.L_HI(net593));
 sg13g2_tiehi _35685__594 (.L_HI(net594));
 sg13g2_tiehi _34749__595 (.L_HI(net595));
 sg13g2_tiehi _35684__596 (.L_HI(net596));
 sg13g2_tiehi _34748__597 (.L_HI(net597));
 sg13g2_tiehi _35683__598 (.L_HI(net598));
 sg13g2_tiehi _34747__599 (.L_HI(net599));
 sg13g2_tiehi _35682__600 (.L_HI(net600));
 sg13g2_tiehi _34746__601 (.L_HI(net601));
 sg13g2_tiehi _35681__602 (.L_HI(net602));
 sg13g2_tiehi _34745__603 (.L_HI(net603));
 sg13g2_tiehi _35680__604 (.L_HI(net604));
 sg13g2_tiehi _34744__605 (.L_HI(net605));
 sg13g2_tiehi _35679__606 (.L_HI(net606));
 sg13g2_tiehi _34743__607 (.L_HI(net607));
 sg13g2_tiehi _35678__608 (.L_HI(net608));
 sg13g2_tiehi _34742__609 (.L_HI(net609));
 sg13g2_tiehi _35677__610 (.L_HI(net610));
 sg13g2_tiehi _34741__611 (.L_HI(net611));
 sg13g2_tiehi _35676__612 (.L_HI(net612));
 sg13g2_tiehi _34740__613 (.L_HI(net613));
 sg13g2_tiehi _35675__614 (.L_HI(net614));
 sg13g2_tiehi _34739__615 (.L_HI(net615));
 sg13g2_tiehi _35674__616 (.L_HI(net616));
 sg13g2_tiehi _34738__617 (.L_HI(net617));
 sg13g2_tiehi _35673__618 (.L_HI(net618));
 sg13g2_tiehi _34737__619 (.L_HI(net619));
 sg13g2_tiehi _35672__620 (.L_HI(net620));
 sg13g2_tiehi _34736__621 (.L_HI(net621));
 sg13g2_tiehi _35671__622 (.L_HI(net622));
 sg13g2_tiehi _34735__623 (.L_HI(net623));
 sg13g2_tiehi _35670__624 (.L_HI(net624));
 sg13g2_tiehi _34734__625 (.L_HI(net625));
 sg13g2_tiehi _35669__626 (.L_HI(net626));
 sg13g2_tiehi _34733__627 (.L_HI(net627));
 sg13g2_tiehi _35668__628 (.L_HI(net628));
 sg13g2_tiehi _34732__629 (.L_HI(net629));
 sg13g2_tiehi _35667__630 (.L_HI(net630));
 sg13g2_tiehi _34731__631 (.L_HI(net631));
 sg13g2_tiehi _35666__632 (.L_HI(net632));
 sg13g2_tiehi _34730__633 (.L_HI(net633));
 sg13g2_tiehi _35665__634 (.L_HI(net634));
 sg13g2_tiehi _34729__635 (.L_HI(net635));
 sg13g2_tiehi _35664__636 (.L_HI(net636));
 sg13g2_tiehi _34728__637 (.L_HI(net637));
 sg13g2_tiehi _35663__638 (.L_HI(net638));
 sg13g2_tiehi _34727__639 (.L_HI(net639));
 sg13g2_tiehi _35662__640 (.L_HI(net640));
 sg13g2_tiehi _34726__641 (.L_HI(net641));
 sg13g2_tiehi _35661__642 (.L_HI(net642));
 sg13g2_tiehi _34725__643 (.L_HI(net643));
 sg13g2_tiehi _35660__644 (.L_HI(net644));
 sg13g2_tiehi _34724__645 (.L_HI(net645));
 sg13g2_tiehi _35659__646 (.L_HI(net646));
 sg13g2_tiehi _34723__647 (.L_HI(net647));
 sg13g2_tiehi _35658__648 (.L_HI(net648));
 sg13g2_tiehi _34722__649 (.L_HI(net649));
 sg13g2_tiehi _35657__650 (.L_HI(net650));
 sg13g2_tiehi _34721__651 (.L_HI(net651));
 sg13g2_tiehi _35656__652 (.L_HI(net652));
 sg13g2_tiehi _34720__653 (.L_HI(net653));
 sg13g2_tiehi _35655__654 (.L_HI(net654));
 sg13g2_tiehi _34719__655 (.L_HI(net655));
 sg13g2_tiehi _35654__656 (.L_HI(net656));
 sg13g2_tiehi _34718__657 (.L_HI(net657));
 sg13g2_tiehi _35653__658 (.L_HI(net658));
 sg13g2_tiehi _34717__659 (.L_HI(net659));
 sg13g2_tiehi _35652__660 (.L_HI(net660));
 sg13g2_tiehi _34716__661 (.L_HI(net661));
 sg13g2_tiehi _35651__662 (.L_HI(net662));
 sg13g2_tiehi _34715__663 (.L_HI(net663));
 sg13g2_tiehi _35650__664 (.L_HI(net664));
 sg13g2_tiehi _34714__665 (.L_HI(net665));
 sg13g2_tiehi _35649__666 (.L_HI(net666));
 sg13g2_tiehi _34713__667 (.L_HI(net667));
 sg13g2_tiehi _35648__668 (.L_HI(net668));
 sg13g2_tiehi _34712__669 (.L_HI(net669));
 sg13g2_tiehi _35647__670 (.L_HI(net670));
 sg13g2_tiehi _34711__671 (.L_HI(net671));
 sg13g2_tiehi _35646__672 (.L_HI(net672));
 sg13g2_tiehi _34710__673 (.L_HI(net673));
 sg13g2_tiehi _35645__674 (.L_HI(net674));
 sg13g2_tiehi _34709__675 (.L_HI(net675));
 sg13g2_tiehi _35644__676 (.L_HI(net676));
 sg13g2_tiehi _34708__677 (.L_HI(net677));
 sg13g2_tiehi _35643__678 (.L_HI(net678));
 sg13g2_tiehi _34707__679 (.L_HI(net679));
 sg13g2_tiehi _35642__680 (.L_HI(net680));
 sg13g2_tiehi _34706__681 (.L_HI(net681));
 sg13g2_tiehi _35641__682 (.L_HI(net682));
 sg13g2_tiehi _34705__683 (.L_HI(net683));
 sg13g2_tiehi _35640__684 (.L_HI(net684));
 sg13g2_tiehi _34704__685 (.L_HI(net685));
 sg13g2_tiehi _35639__686 (.L_HI(net686));
 sg13g2_tiehi _34703__687 (.L_HI(net687));
 sg13g2_tiehi _35638__688 (.L_HI(net688));
 sg13g2_tiehi _34702__689 (.L_HI(net689));
 sg13g2_tiehi _35637__690 (.L_HI(net690));
 sg13g2_tiehi _34701__691 (.L_HI(net691));
 sg13g2_tiehi _35636__692 (.L_HI(net692));
 sg13g2_tiehi _34700__693 (.L_HI(net693));
 sg13g2_tiehi _35635__694 (.L_HI(net694));
 sg13g2_tiehi _34699__695 (.L_HI(net695));
 sg13g2_tiehi _35634__696 (.L_HI(net696));
 sg13g2_tiehi _34698__697 (.L_HI(net697));
 sg13g2_tiehi _35633__698 (.L_HI(net698));
 sg13g2_tiehi _34697__699 (.L_HI(net699));
 sg13g2_tiehi _35632__700 (.L_HI(net700));
 sg13g2_tiehi _34696__701 (.L_HI(net701));
 sg13g2_tiehi _35631__702 (.L_HI(net702));
 sg13g2_tiehi _34695__703 (.L_HI(net703));
 sg13g2_tiehi _35630__704 (.L_HI(net704));
 sg13g2_tiehi _34694__705 (.L_HI(net705));
 sg13g2_tiehi _35629__706 (.L_HI(net706));
 sg13g2_tiehi _34693__707 (.L_HI(net707));
 sg13g2_tiehi _35628__708 (.L_HI(net708));
 sg13g2_tiehi _34692__709 (.L_HI(net709));
 sg13g2_tiehi _35627__710 (.L_HI(net710));
 sg13g2_tiehi _34691__711 (.L_HI(net711));
 sg13g2_tiehi _35626__712 (.L_HI(net712));
 sg13g2_tiehi _34690__713 (.L_HI(net713));
 sg13g2_tiehi _35625__714 (.L_HI(net714));
 sg13g2_tiehi _34689__715 (.L_HI(net715));
 sg13g2_tiehi _35624__716 (.L_HI(net716));
 sg13g2_tiehi _34688__717 (.L_HI(net717));
 sg13g2_tiehi _35623__718 (.L_HI(net718));
 sg13g2_tiehi _34687__719 (.L_HI(net719));
 sg13g2_tiehi _35622__720 (.L_HI(net720));
 sg13g2_tiehi _34686__721 (.L_HI(net721));
 sg13g2_tiehi _35621__722 (.L_HI(net722));
 sg13g2_tiehi _34685__723 (.L_HI(net723));
 sg13g2_tiehi _35620__724 (.L_HI(net724));
 sg13g2_tiehi _34684__725 (.L_HI(net725));
 sg13g2_tiehi _34683__726 (.L_HI(net726));
 sg13g2_tiehi _35619__727 (.L_HI(net727));
 sg13g2_tiehi _34682__728 (.L_HI(net728));
 sg13g2_tiehi _35618__729 (.L_HI(net729));
 sg13g2_tiehi _34681__730 (.L_HI(net730));
 sg13g2_tiehi _35617__731 (.L_HI(net731));
 sg13g2_tiehi _34680__732 (.L_HI(net732));
 sg13g2_tiehi _36170__733 (.L_HI(net733));
 sg13g2_tiehi _34679__734 (.L_HI(net734));
 sg13g2_tiehi _35616__735 (.L_HI(net735));
 sg13g2_tiehi _34678__736 (.L_HI(net736));
 sg13g2_tiehi _34677__737 (.L_HI(net737));
 sg13g2_tiehi _34676__738 (.L_HI(net738));
 sg13g2_tiehi _34675__739 (.L_HI(net739));
 sg13g2_tiehi _34674__740 (.L_HI(net740));
 sg13g2_tiehi _34673__741 (.L_HI(net741));
 sg13g2_tiehi _34672__742 (.L_HI(net742));
 sg13g2_tiehi _34671__743 (.L_HI(net743));
 sg13g2_tiehi _34670__744 (.L_HI(net744));
 sg13g2_tiehi _34669__745 (.L_HI(net745));
 sg13g2_tiehi _34668__746 (.L_HI(net746));
 sg13g2_tiehi _34667__747 (.L_HI(net747));
 sg13g2_tiehi _34666__748 (.L_HI(net748));
 sg13g2_tiehi _34665__749 (.L_HI(net749));
 sg13g2_tiehi _34664__750 (.L_HI(net750));
 sg13g2_tiehi _34663__751 (.L_HI(net751));
 sg13g2_tiehi _34662__752 (.L_HI(net752));
 sg13g2_tiehi _34661__753 (.L_HI(net753));
 sg13g2_tiehi _34660__754 (.L_HI(net754));
 sg13g2_tiehi _34659__755 (.L_HI(net755));
 sg13g2_tiehi _34658__756 (.L_HI(net756));
 sg13g2_tiehi _34657__757 (.L_HI(net757));
 sg13g2_tiehi _34656__758 (.L_HI(net758));
 sg13g2_tiehi _34655__759 (.L_HI(net759));
 sg13g2_tiehi _34654__760 (.L_HI(net760));
 sg13g2_tiehi _34653__761 (.L_HI(net761));
 sg13g2_tiehi _34652__762 (.L_HI(net762));
 sg13g2_tiehi _34651__763 (.L_HI(net763));
 sg13g2_tiehi _34650__764 (.L_HI(net764));
 sg13g2_tiehi _34649__765 (.L_HI(net765));
 sg13g2_tiehi _34648__766 (.L_HI(net766));
 sg13g2_tiehi _34647__767 (.L_HI(net767));
 sg13g2_tiehi _34646__768 (.L_HI(net768));
 sg13g2_tiehi _34645__769 (.L_HI(net769));
 sg13g2_tiehi _36169__770 (.L_HI(net770));
 sg13g2_tiehi _34644__771 (.L_HI(net771));
 sg13g2_tiehi _35615__772 (.L_HI(net772));
 sg13g2_tiehi _34643__773 (.L_HI(net773));
 sg13g2_tiehi _36168__774 (.L_HI(net774));
 sg13g2_tiehi _34642__775 (.L_HI(net775));
 sg13g2_tiehi _35614__776 (.L_HI(net776));
 sg13g2_tiehi _34641__777 (.L_HI(net777));
 sg13g2_tiehi _36167__778 (.L_HI(net778));
 sg13g2_tiehi _34640__779 (.L_HI(net779));
 sg13g2_tiehi _35613__780 (.L_HI(net780));
 sg13g2_tiehi _34639__781 (.L_HI(net781));
 sg13g2_tiehi _34638__782 (.L_HI(net782));
 sg13g2_tiehi _34637__783 (.L_HI(net783));
 sg13g2_tiehi _34636__784 (.L_HI(net784));
 sg13g2_tiehi _34635__785 (.L_HI(net785));
 sg13g2_tiehi _34634__786 (.L_HI(net786));
 sg13g2_tiehi _34633__787 (.L_HI(net787));
 sg13g2_tiehi _34632__788 (.L_HI(net788));
 sg13g2_tiehi _34631__789 (.L_HI(net789));
 sg13g2_tiehi _34630__790 (.L_HI(net790));
 sg13g2_tiehi _34629__791 (.L_HI(net791));
 sg13g2_tiehi _34628__792 (.L_HI(net792));
 sg13g2_tiehi _34627__793 (.L_HI(net793));
 sg13g2_tiehi _34626__794 (.L_HI(net794));
 sg13g2_tiehi _34625__795 (.L_HI(net795));
 sg13g2_tiehi _34624__796 (.L_HI(net796));
 sg13g2_tiehi _34623__797 (.L_HI(net797));
 sg13g2_tiehi _34622__798 (.L_HI(net798));
 sg13g2_tiehi _34621__799 (.L_HI(net799));
 sg13g2_tiehi _34620__800 (.L_HI(net800));
 sg13g2_tiehi _34619__801 (.L_HI(net801));
 sg13g2_tiehi _34618__802 (.L_HI(net802));
 sg13g2_tiehi _34617__803 (.L_HI(net803));
 sg13g2_tiehi _34616__804 (.L_HI(net804));
 sg13g2_tiehi _34615__805 (.L_HI(net805));
 sg13g2_tiehi _34614__806 (.L_HI(net806));
 sg13g2_tiehi _34613__807 (.L_HI(net807));
 sg13g2_tiehi _34612__808 (.L_HI(net808));
 sg13g2_tiehi _34611__809 (.L_HI(net809));
 sg13g2_tiehi _34610__810 (.L_HI(net810));
 sg13g2_tiehi _34609__811 (.L_HI(net811));
 sg13g2_tiehi _34608__812 (.L_HI(net812));
 sg13g2_tiehi _34607__813 (.L_HI(net813));
 sg13g2_tiehi _34606__814 (.L_HI(net814));
 sg13g2_tiehi _34605__815 (.L_HI(net815));
 sg13g2_tiehi _34604__816 (.L_HI(net816));
 sg13g2_tiehi _34603__817 (.L_HI(net817));
 sg13g2_tiehi _34602__818 (.L_HI(net818));
 sg13g2_tiehi _34601__819 (.L_HI(net819));
 sg13g2_tiehi _34600__820 (.L_HI(net820));
 sg13g2_tiehi _34599__821 (.L_HI(net821));
 sg13g2_tiehi _34598__822 (.L_HI(net822));
 sg13g2_tiehi _34597__823 (.L_HI(net823));
 sg13g2_tiehi _34596__824 (.L_HI(net824));
 sg13g2_tiehi _34595__825 (.L_HI(net825));
 sg13g2_tiehi _34594__826 (.L_HI(net826));
 sg13g2_tiehi _34593__827 (.L_HI(net827));
 sg13g2_tiehi _34592__828 (.L_HI(net828));
 sg13g2_tiehi _34591__829 (.L_HI(net829));
 sg13g2_tiehi _34590__830 (.L_HI(net830));
 sg13g2_tiehi _34589__831 (.L_HI(net831));
 sg13g2_tiehi _34588__832 (.L_HI(net832));
 sg13g2_tiehi _34587__833 (.L_HI(net833));
 sg13g2_tiehi _34586__834 (.L_HI(net834));
 sg13g2_tiehi _34585__835 (.L_HI(net835));
 sg13g2_tiehi _34584__836 (.L_HI(net836));
 sg13g2_tiehi _34583__837 (.L_HI(net837));
 sg13g2_tiehi _34582__838 (.L_HI(net838));
 sg13g2_tiehi _34581__839 (.L_HI(net839));
 sg13g2_tiehi _34580__840 (.L_HI(net840));
 sg13g2_tiehi _34579__841 (.L_HI(net841));
 sg13g2_tiehi _34578__842 (.L_HI(net842));
 sg13g2_tiehi _34577__843 (.L_HI(net843));
 sg13g2_tiehi _34576__844 (.L_HI(net844));
 sg13g2_tiehi _34575__845 (.L_HI(net845));
 sg13g2_tiehi _36166__846 (.L_HI(net846));
 sg13g2_tiehi _34574__847 (.L_HI(net847));
 sg13g2_tiehi _35612__848 (.L_HI(net848));
 sg13g2_tiehi _34573__849 (.L_HI(net849));
 sg13g2_tiehi _36165__850 (.L_HI(net850));
 sg13g2_tiehi _34572__851 (.L_HI(net851));
 sg13g2_tiehi _35611__852 (.L_HI(net852));
 sg13g2_tiehi _34571__853 (.L_HI(net853));
 sg13g2_tiehi _36164__854 (.L_HI(net854));
 sg13g2_tiehi _34570__855 (.L_HI(net855));
 sg13g2_tiehi _35610__856 (.L_HI(net856));
 sg13g2_tiehi _34569__857 (.L_HI(net857));
 sg13g2_tiehi _36163__858 (.L_HI(net858));
 sg13g2_tiehi _34568__859 (.L_HI(net859));
 sg13g2_tiehi _35609__860 (.L_HI(net860));
 sg13g2_tiehi _34567__861 (.L_HI(net861));
 sg13g2_tiehi _36162__862 (.L_HI(net862));
 sg13g2_tiehi _34566__863 (.L_HI(net863));
 sg13g2_tiehi _35608__864 (.L_HI(net864));
 sg13g2_tiehi _34565__865 (.L_HI(net865));
 sg13g2_tiehi _36161__866 (.L_HI(net866));
 sg13g2_tiehi _34564__867 (.L_HI(net867));
 sg13g2_tiehi _35607__868 (.L_HI(net868));
 sg13g2_tiehi _34563__869 (.L_HI(net869));
 sg13g2_tiehi _36160__870 (.L_HI(net870));
 sg13g2_tiehi _34562__871 (.L_HI(net871));
 sg13g2_tiehi _35606__872 (.L_HI(net872));
 sg13g2_tiehi _34561__873 (.L_HI(net873));
 sg13g2_tiehi _36159__874 (.L_HI(net874));
 sg13g2_tiehi _34560__875 (.L_HI(net875));
 sg13g2_tiehi _35605__876 (.L_HI(net876));
 sg13g2_tiehi _34559__877 (.L_HI(net877));
 sg13g2_tiehi _36158__878 (.L_HI(net878));
 sg13g2_tiehi _34558__879 (.L_HI(net879));
 sg13g2_tiehi _35604__880 (.L_HI(net880));
 sg13g2_tiehi _34557__881 (.L_HI(net881));
 sg13g2_tiehi _36157__882 (.L_HI(net882));
 sg13g2_tiehi _34556__883 (.L_HI(net883));
 sg13g2_tiehi _35603__884 (.L_HI(net884));
 sg13g2_tiehi _34555__885 (.L_HI(net885));
 sg13g2_tiehi _36156__886 (.L_HI(net886));
 sg13g2_tiehi _34554__887 (.L_HI(net887));
 sg13g2_tiehi _35602__888 (.L_HI(net888));
 sg13g2_tiehi _34553__889 (.L_HI(net889));
 sg13g2_tiehi _36155__890 (.L_HI(net890));
 sg13g2_tiehi _34552__891 (.L_HI(net891));
 sg13g2_tiehi _35601__892 (.L_HI(net892));
 sg13g2_tiehi _34551__893 (.L_HI(net893));
 sg13g2_tiehi _36154__894 (.L_HI(net894));
 sg13g2_tiehi _34550__895 (.L_HI(net895));
 sg13g2_tiehi _35600__896 (.L_HI(net896));
 sg13g2_tiehi _34549__897 (.L_HI(net897));
 sg13g2_tiehi _36153__898 (.L_HI(net898));
 sg13g2_tiehi _34548__899 (.L_HI(net899));
 sg13g2_tiehi _35599__900 (.L_HI(net900));
 sg13g2_tiehi _34547__901 (.L_HI(net901));
 sg13g2_tiehi _36152__902 (.L_HI(net902));
 sg13g2_tiehi _34546__903 (.L_HI(net903));
 sg13g2_tiehi _35598__904 (.L_HI(net904));
 sg13g2_tiehi _34545__905 (.L_HI(net905));
 sg13g2_tiehi _36151__906 (.L_HI(net906));
 sg13g2_tiehi _34544__907 (.L_HI(net907));
 sg13g2_tiehi _35597__908 (.L_HI(net908));
 sg13g2_tiehi _34543__909 (.L_HI(net909));
 sg13g2_tiehi _36150__910 (.L_HI(net910));
 sg13g2_tiehi _34542__911 (.L_HI(net911));
 sg13g2_tiehi _35596__912 (.L_HI(net912));
 sg13g2_tiehi _34541__913 (.L_HI(net913));
 sg13g2_tiehi _36149__914 (.L_HI(net914));
 sg13g2_tiehi _34540__915 (.L_HI(net915));
 sg13g2_tiehi _35595__916 (.L_HI(net916));
 sg13g2_tiehi _34539__917 (.L_HI(net917));
 sg13g2_tiehi _36148__918 (.L_HI(net918));
 sg13g2_tiehi _34538__919 (.L_HI(net919));
 sg13g2_tiehi _35594__920 (.L_HI(net920));
 sg13g2_tiehi _34537__921 (.L_HI(net921));
 sg13g2_tiehi _36147__922 (.L_HI(net922));
 sg13g2_tiehi _34536__923 (.L_HI(net923));
 sg13g2_tiehi _35593__924 (.L_HI(net924));
 sg13g2_tiehi _34535__925 (.L_HI(net925));
 sg13g2_tiehi _36146__926 (.L_HI(net926));
 sg13g2_tiehi _34534__927 (.L_HI(net927));
 sg13g2_tiehi _35592__928 (.L_HI(net928));
 sg13g2_tiehi _34533__929 (.L_HI(net929));
 sg13g2_tiehi _36145__930 (.L_HI(net930));
 sg13g2_tiehi _34532__931 (.L_HI(net931));
 sg13g2_tiehi _35591__932 (.L_HI(net932));
 sg13g2_tiehi _34531__933 (.L_HI(net933));
 sg13g2_tiehi _36144__934 (.L_HI(net934));
 sg13g2_tiehi _34530__935 (.L_HI(net935));
 sg13g2_tiehi _35590__936 (.L_HI(net936));
 sg13g2_tiehi _34529__937 (.L_HI(net937));
 sg13g2_tiehi _36143__938 (.L_HI(net938));
 sg13g2_tiehi _34528__939 (.L_HI(net939));
 sg13g2_tiehi _35589__940 (.L_HI(net940));
 sg13g2_tiehi _34527__941 (.L_HI(net941));
 sg13g2_tiehi _36142__942 (.L_HI(net942));
 sg13g2_tiehi _34526__943 (.L_HI(net943));
 sg13g2_tiehi _35588__944 (.L_HI(net944));
 sg13g2_tiehi _34525__945 (.L_HI(net945));
 sg13g2_tiehi _36141__946 (.L_HI(net946));
 sg13g2_tiehi _34524__947 (.L_HI(net947));
 sg13g2_tiehi _35587__948 (.L_HI(net948));
 sg13g2_tiehi _34523__949 (.L_HI(net949));
 sg13g2_tiehi _36140__950 (.L_HI(net950));
 sg13g2_tiehi _34522__951 (.L_HI(net951));
 sg13g2_tiehi _35586__952 (.L_HI(net952));
 sg13g2_tiehi _34521__953 (.L_HI(net953));
 sg13g2_tiehi _36139__954 (.L_HI(net954));
 sg13g2_tiehi _34520__955 (.L_HI(net955));
 sg13g2_tiehi _35585__956 (.L_HI(net956));
 sg13g2_tiehi _34519__957 (.L_HI(net957));
 sg13g2_tiehi _36138__958 (.L_HI(net958));
 sg13g2_tiehi _34518__959 (.L_HI(net959));
 sg13g2_tiehi _35584__960 (.L_HI(net960));
 sg13g2_tiehi _34517__961 (.L_HI(net961));
 sg13g2_tiehi _36137__962 (.L_HI(net962));
 sg13g2_tiehi _34516__963 (.L_HI(net963));
 sg13g2_tiehi _35583__964 (.L_HI(net964));
 sg13g2_tiehi _34515__965 (.L_HI(net965));
 sg13g2_tiehi _36136__966 (.L_HI(net966));
 sg13g2_tiehi _34514__967 (.L_HI(net967));
 sg13g2_tiehi _35582__968 (.L_HI(net968));
 sg13g2_tiehi _34513__969 (.L_HI(net969));
 sg13g2_tiehi _36135__970 (.L_HI(net970));
 sg13g2_tiehi _34512__971 (.L_HI(net971));
 sg13g2_tiehi _35581__972 (.L_HI(net972));
 sg13g2_tiehi _34511__973 (.L_HI(net973));
 sg13g2_tiehi _36134__974 (.L_HI(net974));
 sg13g2_tiehi _34510__975 (.L_HI(net975));
 sg13g2_tiehi _35580__976 (.L_HI(net976));
 sg13g2_tiehi _34509__977 (.L_HI(net977));
 sg13g2_tiehi _36133__978 (.L_HI(net978));
 sg13g2_tiehi _34508__979 (.L_HI(net979));
 sg13g2_tiehi _35579__980 (.L_HI(net980));
 sg13g2_tiehi _34507__981 (.L_HI(net981));
 sg13g2_tiehi _36132__982 (.L_HI(net982));
 sg13g2_tiehi _34506__983 (.L_HI(net983));
 sg13g2_tiehi _35578__984 (.L_HI(net984));
 sg13g2_tiehi _34505__985 (.L_HI(net985));
 sg13g2_tiehi _36131__986 (.L_HI(net986));
 sg13g2_tiehi _34504__987 (.L_HI(net987));
 sg13g2_tiehi _35577__988 (.L_HI(net988));
 sg13g2_tiehi _34503__989 (.L_HI(net989));
 sg13g2_tiehi _36130__990 (.L_HI(net990));
 sg13g2_tiehi _34502__991 (.L_HI(net991));
 sg13g2_tiehi _35576__992 (.L_HI(net992));
 sg13g2_tiehi _34501__993 (.L_HI(net993));
 sg13g2_tiehi _36129__994 (.L_HI(net994));
 sg13g2_tiehi _34500__995 (.L_HI(net995));
 sg13g2_tiehi _35575__996 (.L_HI(net996));
 sg13g2_tiehi _34499__997 (.L_HI(net997));
 sg13g2_tiehi _36128__998 (.L_HI(net998));
 sg13g2_tiehi _34498__999 (.L_HI(net999));
 sg13g2_tiehi _35574__1000 (.L_HI(net1000));
 sg13g2_tiehi _34497__1001 (.L_HI(net1001));
 sg13g2_tiehi _36127__1002 (.L_HI(net1002));
 sg13g2_tiehi _34496__1003 (.L_HI(net1003));
 sg13g2_tiehi _35573__1004 (.L_HI(net1004));
 sg13g2_tiehi _34495__1005 (.L_HI(net1005));
 sg13g2_tiehi _36126__1006 (.L_HI(net1006));
 sg13g2_tiehi _34494__1007 (.L_HI(net1007));
 sg13g2_tiehi _35572__1008 (.L_HI(net1008));
 sg13g2_tiehi _34493__1009 (.L_HI(net1009));
 sg13g2_tiehi _36125__1010 (.L_HI(net1010));
 sg13g2_tiehi _34492__1011 (.L_HI(net1011));
 sg13g2_tiehi _35571__1012 (.L_HI(net1012));
 sg13g2_tiehi _34491__1013 (.L_HI(net1013));
 sg13g2_tiehi _36124__1014 (.L_HI(net1014));
 sg13g2_tiehi _34490__1015 (.L_HI(net1015));
 sg13g2_tiehi _35570__1016 (.L_HI(net1016));
 sg13g2_tiehi _34489__1017 (.L_HI(net1017));
 sg13g2_tiehi _36123__1018 (.L_HI(net1018));
 sg13g2_tiehi _34488__1019 (.L_HI(net1019));
 sg13g2_tiehi _35569__1020 (.L_HI(net1020));
 sg13g2_tiehi _34487__1021 (.L_HI(net1021));
 sg13g2_tiehi _36122__1022 (.L_HI(net1022));
 sg13g2_tiehi _34486__1023 (.L_HI(net1023));
 sg13g2_tiehi _35568__1024 (.L_HI(net1024));
 sg13g2_tiehi _34485__1025 (.L_HI(net1025));
 sg13g2_tiehi _36121__1026 (.L_HI(net1026));
 sg13g2_tiehi _34484__1027 (.L_HI(net1027));
 sg13g2_tiehi _35567__1028 (.L_HI(net1028));
 sg13g2_tiehi _34483__1029 (.L_HI(net1029));
 sg13g2_tiehi _36120__1030 (.L_HI(net1030));
 sg13g2_tiehi _34482__1031 (.L_HI(net1031));
 sg13g2_tiehi _35566__1032 (.L_HI(net1032));
 sg13g2_tiehi _34481__1033 (.L_HI(net1033));
 sg13g2_tiehi _36119__1034 (.L_HI(net1034));
 sg13g2_tiehi _34480__1035 (.L_HI(net1035));
 sg13g2_tiehi _35565__1036 (.L_HI(net1036));
 sg13g2_tiehi _34479__1037 (.L_HI(net1037));
 sg13g2_tiehi _36118__1038 (.L_HI(net1038));
 sg13g2_tiehi _34478__1039 (.L_HI(net1039));
 sg13g2_tiehi _35564__1040 (.L_HI(net1040));
 sg13g2_tiehi _34477__1041 (.L_HI(net1041));
 sg13g2_tiehi _36117__1042 (.L_HI(net1042));
 sg13g2_tiehi _34476__1043 (.L_HI(net1043));
 sg13g2_tiehi _35563__1044 (.L_HI(net1044));
 sg13g2_tiehi _34475__1045 (.L_HI(net1045));
 sg13g2_tiehi _36116__1046 (.L_HI(net1046));
 sg13g2_tiehi _34474__1047 (.L_HI(net1047));
 sg13g2_tiehi _35562__1048 (.L_HI(net1048));
 sg13g2_tiehi _34473__1049 (.L_HI(net1049));
 sg13g2_tiehi _36115__1050 (.L_HI(net1050));
 sg13g2_tiehi _34472__1051 (.L_HI(net1051));
 sg13g2_tiehi _35561__1052 (.L_HI(net1052));
 sg13g2_tiehi _34471__1053 (.L_HI(net1053));
 sg13g2_tiehi _36114__1054 (.L_HI(net1054));
 sg13g2_tiehi _34470__1055 (.L_HI(net1055));
 sg13g2_tiehi _35560__1056 (.L_HI(net1056));
 sg13g2_tiehi _34469__1057 (.L_HI(net1057));
 sg13g2_tiehi _36113__1058 (.L_HI(net1058));
 sg13g2_tiehi _34468__1059 (.L_HI(net1059));
 sg13g2_tiehi _35559__1060 (.L_HI(net1060));
 sg13g2_tiehi _34467__1061 (.L_HI(net1061));
 sg13g2_tiehi _36112__1062 (.L_HI(net1062));
 sg13g2_tiehi _34466__1063 (.L_HI(net1063));
 sg13g2_tiehi _35558__1064 (.L_HI(net1064));
 sg13g2_tiehi _34465__1065 (.L_HI(net1065));
 sg13g2_tiehi _36111__1066 (.L_HI(net1066));
 sg13g2_tiehi _34464__1067 (.L_HI(net1067));
 sg13g2_tiehi _35557__1068 (.L_HI(net1068));
 sg13g2_tiehi _34463__1069 (.L_HI(net1069));
 sg13g2_tiehi _36110__1070 (.L_HI(net1070));
 sg13g2_tiehi _34462__1071 (.L_HI(net1071));
 sg13g2_tiehi _35556__1072 (.L_HI(net1072));
 sg13g2_tiehi _34461__1073 (.L_HI(net1073));
 sg13g2_tiehi _36109__1074 (.L_HI(net1074));
 sg13g2_tiehi _34460__1075 (.L_HI(net1075));
 sg13g2_tiehi _35555__1076 (.L_HI(net1076));
 sg13g2_tiehi _34459__1077 (.L_HI(net1077));
 sg13g2_tiehi _36108__1078 (.L_HI(net1078));
 sg13g2_tiehi _34458__1079 (.L_HI(net1079));
 sg13g2_tiehi _35554__1080 (.L_HI(net1080));
 sg13g2_tiehi _34457__1081 (.L_HI(net1081));
 sg13g2_tiehi _36107__1082 (.L_HI(net1082));
 sg13g2_tiehi _34456__1083 (.L_HI(net1083));
 sg13g2_tiehi _35553__1084 (.L_HI(net1084));
 sg13g2_tiehi _34455__1085 (.L_HI(net1085));
 sg13g2_tiehi _35552__1086 (.L_HI(net1086));
 sg13g2_tiehi _34454__1087 (.L_HI(net1087));
 sg13g2_tiehi _35551__1088 (.L_HI(net1088));
 sg13g2_tiehi _34453__1089 (.L_HI(net1089));
 sg13g2_tiehi _35550__1090 (.L_HI(net1090));
 sg13g2_tiehi _34452__1091 (.L_HI(net1091));
 sg13g2_tiehi _35549__1092 (.L_HI(net1092));
 sg13g2_tiehi _34451__1093 (.L_HI(net1093));
 sg13g2_tiehi _36106__1094 (.L_HI(net1094));
 sg13g2_tiehi _34450__1095 (.L_HI(net1095));
 sg13g2_tiehi _35548__1096 (.L_HI(net1096));
 sg13g2_tiehi _34449__1097 (.L_HI(net1097));
 sg13g2_tiehi _36105__1098 (.L_HI(net1098));
 sg13g2_tiehi _34448__1099 (.L_HI(net1099));
 sg13g2_tiehi _35547__1100 (.L_HI(net1100));
 sg13g2_tiehi _34447__1101 (.L_HI(net1101));
 sg13g2_tiehi _34446__1102 (.L_HI(net1102));
 sg13g2_tiehi _34445__1103 (.L_HI(net1103));
 sg13g2_tiehi _34444__1104 (.L_HI(net1104));
 sg13g2_tiehi _34443__1105 (.L_HI(net1105));
 sg13g2_tiehi _34442__1106 (.L_HI(net1106));
 sg13g2_tiehi _34441__1107 (.L_HI(net1107));
 sg13g2_tiehi _34440__1108 (.L_HI(net1108));
 sg13g2_tiehi _34439__1109 (.L_HI(net1109));
 sg13g2_tiehi _34438__1110 (.L_HI(net1110));
 sg13g2_tiehi _34437__1111 (.L_HI(net1111));
 sg13g2_tiehi _34436__1112 (.L_HI(net1112));
 sg13g2_tiehi _34435__1113 (.L_HI(net1113));
 sg13g2_tiehi _34434__1114 (.L_HI(net1114));
 sg13g2_tiehi _34433__1115 (.L_HI(net1115));
 sg13g2_tiehi _34432__1116 (.L_HI(net1116));
 sg13g2_tiehi _34431__1117 (.L_HI(net1117));
 sg13g2_tiehi _34430__1118 (.L_HI(net1118));
 sg13g2_tiehi _34429__1119 (.L_HI(net1119));
 sg13g2_tiehi _34428__1120 (.L_HI(net1120));
 sg13g2_tiehi _34427__1121 (.L_HI(net1121));
 sg13g2_tiehi _34426__1122 (.L_HI(net1122));
 sg13g2_tiehi _34425__1123 (.L_HI(net1123));
 sg13g2_tiehi _34424__1124 (.L_HI(net1124));
 sg13g2_tiehi _34423__1125 (.L_HI(net1125));
 sg13g2_tiehi _34422__1126 (.L_HI(net1126));
 sg13g2_tiehi _34421__1127 (.L_HI(net1127));
 sg13g2_tiehi _34420__1128 (.L_HI(net1128));
 sg13g2_tiehi _34419__1129 (.L_HI(net1129));
 sg13g2_tiehi _34418__1130 (.L_HI(net1130));
 sg13g2_tiehi _34417__1131 (.L_HI(net1131));
 sg13g2_tiehi _34416__1132 (.L_HI(net1132));
 sg13g2_tiehi _34415__1133 (.L_HI(net1133));
 sg13g2_tiehi _34414__1134 (.L_HI(net1134));
 sg13g2_tiehi _34413__1135 (.L_HI(net1135));
 sg13g2_tiehi _34412__1136 (.L_HI(net1136));
 sg13g2_tiehi _34411__1137 (.L_HI(net1137));
 sg13g2_tiehi _34410__1138 (.L_HI(net1138));
 sg13g2_tiehi _34409__1139 (.L_HI(net1139));
 sg13g2_tiehi _34408__1140 (.L_HI(net1140));
 sg13g2_tiehi _34407__1141 (.L_HI(net1141));
 sg13g2_tiehi _34406__1142 (.L_HI(net1142));
 sg13g2_tiehi _34405__1143 (.L_HI(net1143));
 sg13g2_tiehi _34404__1144 (.L_HI(net1144));
 sg13g2_tiehi _34403__1145 (.L_HI(net1145));
 sg13g2_tiehi _34402__1146 (.L_HI(net1146));
 sg13g2_tiehi _34401__1147 (.L_HI(net1147));
 sg13g2_tiehi _34400__1148 (.L_HI(net1148));
 sg13g2_tiehi _34399__1149 (.L_HI(net1149));
 sg13g2_tiehi _34398__1150 (.L_HI(net1150));
 sg13g2_tiehi _34397__1151 (.L_HI(net1151));
 sg13g2_tiehi _34396__1152 (.L_HI(net1152));
 sg13g2_tiehi _34395__1153 (.L_HI(net1153));
 sg13g2_tiehi _34394__1154 (.L_HI(net1154));
 sg13g2_tiehi _34393__1155 (.L_HI(net1155));
 sg13g2_tiehi _34392__1156 (.L_HI(net1156));
 sg13g2_tiehi _34391__1157 (.L_HI(net1157));
 sg13g2_tiehi _34390__1158 (.L_HI(net1158));
 sg13g2_tiehi _34389__1159 (.L_HI(net1159));
 sg13g2_tiehi _34388__1160 (.L_HI(net1160));
 sg13g2_tiehi _34387__1161 (.L_HI(net1161));
 sg13g2_tiehi _34386__1162 (.L_HI(net1162));
 sg13g2_tiehi _34385__1163 (.L_HI(net1163));
 sg13g2_tiehi _34384__1164 (.L_HI(net1164));
 sg13g2_tiehi _34383__1165 (.L_HI(net1165));
 sg13g2_tiehi _36104__1166 (.L_HI(net1166));
 sg13g2_tiehi _34382__1167 (.L_HI(net1167));
 sg13g2_tiehi _35546__1168 (.L_HI(net1168));
 sg13g2_tiehi _34381__1169 (.L_HI(net1169));
 sg13g2_tiehi _36103__1170 (.L_HI(net1170));
 sg13g2_tiehi _34380__1171 (.L_HI(net1171));
 sg13g2_tiehi _35545__1172 (.L_HI(net1172));
 sg13g2_tiehi _34379__1173 (.L_HI(net1173));
 sg13g2_tiehi _36102__1174 (.L_HI(net1174));
 sg13g2_tiehi _34378__1175 (.L_HI(net1175));
 sg13g2_tiehi _35544__1176 (.L_HI(net1176));
 sg13g2_tiehi _34377__1177 (.L_HI(net1177));
 sg13g2_tiehi _36101__1178 (.L_HI(net1178));
 sg13g2_tiehi _34376__1179 (.L_HI(net1179));
 sg13g2_tiehi _35543__1180 (.L_HI(net1180));
 sg13g2_tiehi _34375__1181 (.L_HI(net1181));
 sg13g2_tiehi _36100__1182 (.L_HI(net1182));
 sg13g2_tiehi _34374__1183 (.L_HI(net1183));
 sg13g2_tiehi _35542__1184 (.L_HI(net1184));
 sg13g2_tiehi _34373__1185 (.L_HI(net1185));
 sg13g2_tiehi _36099__1186 (.L_HI(net1186));
 sg13g2_tiehi _34372__1187 (.L_HI(net1187));
 sg13g2_tiehi _35541__1188 (.L_HI(net1188));
 sg13g2_tiehi _34371__1189 (.L_HI(net1189));
 sg13g2_tiehi _36098__1190 (.L_HI(net1190));
 sg13g2_tiehi _34370__1191 (.L_HI(net1191));
 sg13g2_tiehi _35540__1192 (.L_HI(net1192));
 sg13g2_tiehi _34369__1193 (.L_HI(net1193));
 sg13g2_tiehi _36097__1194 (.L_HI(net1194));
 sg13g2_tiehi _34368__1195 (.L_HI(net1195));
 sg13g2_tiehi _35539__1196 (.L_HI(net1196));
 sg13g2_tiehi _34367__1197 (.L_HI(net1197));
 sg13g2_tiehi _36096__1198 (.L_HI(net1198));
 sg13g2_tiehi _34366__1199 (.L_HI(net1199));
 sg13g2_tiehi _35538__1200 (.L_HI(net1200));
 sg13g2_tiehi _34365__1201 (.L_HI(net1201));
 sg13g2_tiehi _36095__1202 (.L_HI(net1202));
 sg13g2_tiehi _34364__1203 (.L_HI(net1203));
 sg13g2_tiehi _35537__1204 (.L_HI(net1204));
 sg13g2_tiehi _34363__1205 (.L_HI(net1205));
 sg13g2_tiehi _36094__1206 (.L_HI(net1206));
 sg13g2_tiehi _34362__1207 (.L_HI(net1207));
 sg13g2_tiehi _35536__1208 (.L_HI(net1208));
 sg13g2_tiehi _34361__1209 (.L_HI(net1209));
 sg13g2_tiehi _36093__1210 (.L_HI(net1210));
 sg13g2_tiehi _34360__1211 (.L_HI(net1211));
 sg13g2_tiehi _35535__1212 (.L_HI(net1212));
 sg13g2_tiehi _34359__1213 (.L_HI(net1213));
 sg13g2_tiehi _36092__1214 (.L_HI(net1214));
 sg13g2_tiehi _34358__1215 (.L_HI(net1215));
 sg13g2_tiehi _35534__1216 (.L_HI(net1216));
 sg13g2_tiehi _34357__1217 (.L_HI(net1217));
 sg13g2_tiehi _36091__1218 (.L_HI(net1218));
 sg13g2_tiehi _34356__1219 (.L_HI(net1219));
 sg13g2_tiehi _35533__1220 (.L_HI(net1220));
 sg13g2_tiehi _34355__1221 (.L_HI(net1221));
 sg13g2_tiehi _36090__1222 (.L_HI(net1222));
 sg13g2_tiehi _34354__1223 (.L_HI(net1223));
 sg13g2_tiehi _35532__1224 (.L_HI(net1224));
 sg13g2_tiehi _34353__1225 (.L_HI(net1225));
 sg13g2_tiehi _36089__1226 (.L_HI(net1226));
 sg13g2_tiehi _34352__1227 (.L_HI(net1227));
 sg13g2_tiehi _35531__1228 (.L_HI(net1228));
 sg13g2_tiehi _34351__1229 (.L_HI(net1229));
 sg13g2_tiehi _36088__1230 (.L_HI(net1230));
 sg13g2_tiehi _34350__1231 (.L_HI(net1231));
 sg13g2_tiehi _35530__1232 (.L_HI(net1232));
 sg13g2_tiehi _34349__1233 (.L_HI(net1233));
 sg13g2_tiehi _36087__1234 (.L_HI(net1234));
 sg13g2_tiehi _34348__1235 (.L_HI(net1235));
 sg13g2_tiehi _35529__1236 (.L_HI(net1236));
 sg13g2_tiehi _34347__1237 (.L_HI(net1237));
 sg13g2_tiehi _36086__1238 (.L_HI(net1238));
 sg13g2_tiehi _34346__1239 (.L_HI(net1239));
 sg13g2_tiehi _35528__1240 (.L_HI(net1240));
 sg13g2_tiehi _34345__1241 (.L_HI(net1241));
 sg13g2_tiehi _36085__1242 (.L_HI(net1242));
 sg13g2_tiehi _34344__1243 (.L_HI(net1243));
 sg13g2_tiehi _35527__1244 (.L_HI(net1244));
 sg13g2_tiehi _34343__1245 (.L_HI(net1245));
 sg13g2_tiehi _36084__1246 (.L_HI(net1246));
 sg13g2_tiehi _34342__1247 (.L_HI(net1247));
 sg13g2_tiehi _35526__1248 (.L_HI(net1248));
 sg13g2_tiehi _34341__1249 (.L_HI(net1249));
 sg13g2_tiehi _36083__1250 (.L_HI(net1250));
 sg13g2_tiehi _34340__1251 (.L_HI(net1251));
 sg13g2_tiehi _35525__1252 (.L_HI(net1252));
 sg13g2_tiehi _34339__1253 (.L_HI(net1253));
 sg13g2_tiehi _36082__1254 (.L_HI(net1254));
 sg13g2_tiehi _34338__1255 (.L_HI(net1255));
 sg13g2_tiehi _35524__1256 (.L_HI(net1256));
 sg13g2_tiehi _34337__1257 (.L_HI(net1257));
 sg13g2_tiehi _36081__1258 (.L_HI(net1258));
 sg13g2_tiehi _34336__1259 (.L_HI(net1259));
 sg13g2_tiehi _35523__1260 (.L_HI(net1260));
 sg13g2_tiehi _34335__1261 (.L_HI(net1261));
 sg13g2_tiehi _36080__1262 (.L_HI(net1262));
 sg13g2_tiehi _34334__1263 (.L_HI(net1263));
 sg13g2_tiehi _35522__1264 (.L_HI(net1264));
 sg13g2_tiehi _34333__1265 (.L_HI(net1265));
 sg13g2_tiehi _36079__1266 (.L_HI(net1266));
 sg13g2_tiehi _34332__1267 (.L_HI(net1267));
 sg13g2_tiehi _35521__1268 (.L_HI(net1268));
 sg13g2_tiehi _34331__1269 (.L_HI(net1269));
 sg13g2_tiehi _36078__1270 (.L_HI(net1270));
 sg13g2_tiehi _34330__1271 (.L_HI(net1271));
 sg13g2_tiehi _35520__1272 (.L_HI(net1272));
 sg13g2_tiehi _34329__1273 (.L_HI(net1273));
 sg13g2_tiehi _36077__1274 (.L_HI(net1274));
 sg13g2_tiehi _34328__1275 (.L_HI(net1275));
 sg13g2_tiehi _35519__1276 (.L_HI(net1276));
 sg13g2_tiehi _34327__1277 (.L_HI(net1277));
 sg13g2_tiehi _36076__1278 (.L_HI(net1278));
 sg13g2_tiehi _34326__1279 (.L_HI(net1279));
 sg13g2_tiehi _35518__1280 (.L_HI(net1280));
 sg13g2_tiehi _34325__1281 (.L_HI(net1281));
 sg13g2_tiehi _36075__1282 (.L_HI(net1282));
 sg13g2_tiehi _34324__1283 (.L_HI(net1283));
 sg13g2_tiehi _35517__1284 (.L_HI(net1284));
 sg13g2_tiehi _34323__1285 (.L_HI(net1285));
 sg13g2_tiehi _36074__1286 (.L_HI(net1286));
 sg13g2_tiehi _34322__1287 (.L_HI(net1287));
 sg13g2_tiehi _35516__1288 (.L_HI(net1288));
 sg13g2_tiehi _34321__1289 (.L_HI(net1289));
 sg13g2_tiehi _35515__1290 (.L_HI(net1290));
 sg13g2_tiehi _34320__1291 (.L_HI(net1291));
 sg13g2_tiehi _35514__1292 (.L_HI(net1292));
 sg13g2_tiehi _34319__1293 (.L_HI(net1293));
 sg13g2_tiehi _35513__1294 (.L_HI(net1294));
 sg13g2_tiehi _34318__1295 (.L_HI(net1295));
 sg13g2_tiehi _35512__1296 (.L_HI(net1296));
 sg13g2_tiehi _34317__1297 (.L_HI(net1297));
 sg13g2_tiehi _35511__1298 (.L_HI(net1298));
 sg13g2_tiehi _34316__1299 (.L_HI(net1299));
 sg13g2_tiehi _35510__1300 (.L_HI(net1300));
 sg13g2_tiehi _34315__1301 (.L_HI(net1301));
 sg13g2_tiehi _35509__1302 (.L_HI(net1302));
 sg13g2_tiehi _34314__1303 (.L_HI(net1303));
 sg13g2_tiehi _35508__1304 (.L_HI(net1304));
 sg13g2_tiehi _34313__1305 (.L_HI(net1305));
 sg13g2_tiehi _34312__1306 (.L_HI(net1306));
 sg13g2_tiehi _34311__1307 (.L_HI(net1307));
 sg13g2_tiehi _33616__1308 (.L_HI(net1308));
 sg13g2_tiehi _34909__1309 (.L_HI(net1309));
 sg13g2_tiehi _34910__1310 (.L_HI(net1310));
 sg13g2_tiehi _34911__1311 (.L_HI(net1311));
 sg13g2_tiehi _34912__1312 (.L_HI(net1312));
 sg13g2_tiehi _34913__1313 (.L_HI(net1313));
 sg13g2_tiehi _34914__1314 (.L_HI(net1314));
 sg13g2_tiehi _34915__1315 (.L_HI(net1315));
 sg13g2_tiehi _34916__1316 (.L_HI(net1316));
 sg13g2_tiehi _34917__1317 (.L_HI(net1317));
 sg13g2_tiehi _34918__1318 (.L_HI(net1318));
 sg13g2_tiehi _34919__1319 (.L_HI(net1319));
 sg13g2_tiehi _34920__1320 (.L_HI(net1320));
 sg13g2_tiehi _34921__1321 (.L_HI(net1321));
 sg13g2_tiehi _34922__1322 (.L_HI(net1322));
 sg13g2_tiehi _34923__1323 (.L_HI(net1323));
 sg13g2_tiehi _34924__1324 (.L_HI(net1324));
 sg13g2_tiehi _34925__1325 (.L_HI(net1325));
 sg13g2_tiehi _34926__1326 (.L_HI(net1326));
 sg13g2_tiehi _34927__1327 (.L_HI(net1327));
 sg13g2_tiehi _34928__1328 (.L_HI(net1328));
 sg13g2_tiehi _34929__1329 (.L_HI(net1329));
 sg13g2_tiehi _34930__1330 (.L_HI(net1330));
 sg13g2_tiehi _34931__1331 (.L_HI(net1331));
 sg13g2_tiehi _34932__1332 (.L_HI(net1332));
 sg13g2_tiehi _34933__1333 (.L_HI(net1333));
 sg13g2_tiehi _34934__1334 (.L_HI(net1334));
 sg13g2_tiehi _34935__1335 (.L_HI(net1335));
 sg13g2_tiehi _34936__1336 (.L_HI(net1336));
 sg13g2_tiehi _34937__1337 (.L_HI(net1337));
 sg13g2_tiehi _34938__1338 (.L_HI(net1338));
 sg13g2_tiehi _34939__1339 (.L_HI(net1339));
 sg13g2_tiehi _34940__1340 (.L_HI(net1340));
 sg13g2_tiehi _34941__1341 (.L_HI(net1341));
 sg13g2_tiehi _34942__1342 (.L_HI(net1342));
 sg13g2_tiehi _34943__1343 (.L_HI(net1343));
 sg13g2_tiehi _34944__1344 (.L_HI(net1344));
 sg13g2_tiehi _34945__1345 (.L_HI(net1345));
 sg13g2_tiehi _34946__1346 (.L_HI(net1346));
 sg13g2_tiehi _34947__1347 (.L_HI(net1347));
 sg13g2_tiehi _34948__1348 (.L_HI(net1348));
 sg13g2_tiehi _34949__1349 (.L_HI(net1349));
 sg13g2_tiehi _34950__1350 (.L_HI(net1350));
 sg13g2_tiehi _34951__1351 (.L_HI(net1351));
 sg13g2_tiehi _34952__1352 (.L_HI(net1352));
 sg13g2_tiehi _34953__1353 (.L_HI(net1353));
 sg13g2_tiehi _34954__1354 (.L_HI(net1354));
 sg13g2_tiehi _34955__1355 (.L_HI(net1355));
 sg13g2_tiehi _34956__1356 (.L_HI(net1356));
 sg13g2_tiehi _34957__1357 (.L_HI(net1357));
 sg13g2_tiehi _34958__1358 (.L_HI(net1358));
 sg13g2_tiehi _34959__1359 (.L_HI(net1359));
 sg13g2_tiehi _34960__1360 (.L_HI(net1360));
 sg13g2_tiehi _34961__1361 (.L_HI(net1361));
 sg13g2_tiehi _34962__1362 (.L_HI(net1362));
 sg13g2_tiehi _34963__1363 (.L_HI(net1363));
 sg13g2_tiehi _34964__1364 (.L_HI(net1364));
 sg13g2_tiehi _34965__1365 (.L_HI(net1365));
 sg13g2_tiehi _34966__1366 (.L_HI(net1366));
 sg13g2_tiehi _34967__1367 (.L_HI(net1367));
 sg13g2_tiehi _34968__1368 (.L_HI(net1368));
 sg13g2_tiehi _34969__1369 (.L_HI(net1369));
 sg13g2_tiehi _34970__1370 (.L_HI(net1370));
 sg13g2_tiehi _34971__1371 (.L_HI(net1371));
 sg13g2_tiehi _34972__1372 (.L_HI(net1372));
 sg13g2_tiehi _34973__1373 (.L_HI(net1373));
 sg13g2_tiehi _34974__1374 (.L_HI(net1374));
 sg13g2_tiehi _34975__1375 (.L_HI(net1375));
 sg13g2_tiehi _34976__1376 (.L_HI(net1376));
 sg13g2_tiehi _34977__1377 (.L_HI(net1377));
 sg13g2_tiehi _34978__1378 (.L_HI(net1378));
 sg13g2_tiehi _34979__1379 (.L_HI(net1379));
 sg13g2_tiehi _34980__1380 (.L_HI(net1380));
 sg13g2_tiehi _34981__1381 (.L_HI(net1381));
 sg13g2_tiehi _34982__1382 (.L_HI(net1382));
 sg13g2_tiehi _34983__1383 (.L_HI(net1383));
 sg13g2_tiehi _34984__1384 (.L_HI(net1384));
 sg13g2_tiehi _34985__1385 (.L_HI(net1385));
 sg13g2_tiehi _34986__1386 (.L_HI(net1386));
 sg13g2_tiehi _34987__1387 (.L_HI(net1387));
 sg13g2_tiehi _34988__1388 (.L_HI(net1388));
 sg13g2_tiehi _34989__1389 (.L_HI(net1389));
 sg13g2_tiehi _34990__1390 (.L_HI(net1390));
 sg13g2_tiehi _34991__1391 (.L_HI(net1391));
 sg13g2_tiehi _34992__1392 (.L_HI(net1392));
 sg13g2_tiehi _34993__1393 (.L_HI(net1393));
 sg13g2_tiehi _34994__1394 (.L_HI(net1394));
 sg13g2_tiehi _34995__1395 (.L_HI(net1395));
 sg13g2_tiehi _34996__1396 (.L_HI(net1396));
 sg13g2_tiehi _34997__1397 (.L_HI(net1397));
 sg13g2_tiehi _34998__1398 (.L_HI(net1398));
 sg13g2_tiehi _34999__1399 (.L_HI(net1399));
 sg13g2_tiehi _35000__1400 (.L_HI(net1400));
 sg13g2_tiehi _35001__1401 (.L_HI(net1401));
 sg13g2_tiehi _35002__1402 (.L_HI(net1402));
 sg13g2_tiehi _35003__1403 (.L_HI(net1403));
 sg13g2_tiehi _34310__1404 (.L_HI(net1404));
 sg13g2_tiehi _35004__1405 (.L_HI(net1405));
 sg13g2_tiehi _35006__1406 (.L_HI(net1406));
 sg13g2_tiehi _35507__1407 (.L_HI(net1407));
 sg13g2_tiehi _34309__1408 (.L_HI(net1408));
 sg13g2_tiehi _35506__1409 (.L_HI(net1409));
 sg13g2_tiehi _34308__1410 (.L_HI(net1410));
 sg13g2_tiehi _36073__1411 (.L_HI(net1411));
 sg13g2_tiehi _34307__1412 (.L_HI(net1412));
 sg13g2_tiehi _35505__1413 (.L_HI(net1413));
 sg13g2_tiehi _34306__1414 (.L_HI(net1414));
 sg13g2_tiehi _36072__1415 (.L_HI(net1415));
 sg13g2_tiehi _34305__1416 (.L_HI(net1416));
 sg13g2_tiehi _35504__1417 (.L_HI(net1417));
 sg13g2_tiehi _34304__1418 (.L_HI(net1418));
 sg13g2_tiehi _36071__1419 (.L_HI(net1419));
 sg13g2_tiehi _34303__1420 (.L_HI(net1420));
 sg13g2_tiehi _35503__1421 (.L_HI(net1421));
 sg13g2_tiehi _34302__1422 (.L_HI(net1422));
 sg13g2_tiehi _36070__1423 (.L_HI(net1423));
 sg13g2_tiehi _34301__1424 (.L_HI(net1424));
 sg13g2_tiehi _35502__1425 (.L_HI(net1425));
 sg13g2_tiehi _34300__1426 (.L_HI(net1426));
 sg13g2_tiehi _36069__1427 (.L_HI(net1427));
 sg13g2_tiehi _34299__1428 (.L_HI(net1428));
 sg13g2_tiehi _35501__1429 (.L_HI(net1429));
 sg13g2_tiehi _34298__1430 (.L_HI(net1430));
 sg13g2_tiehi _36068__1431 (.L_HI(net1431));
 sg13g2_tiehi _34297__1432 (.L_HI(net1432));
 sg13g2_tiehi _35500__1433 (.L_HI(net1433));
 sg13g2_tiehi _34296__1434 (.L_HI(net1434));
 sg13g2_tiehi _36067__1435 (.L_HI(net1435));
 sg13g2_tiehi _34295__1436 (.L_HI(net1436));
 sg13g2_tiehi _35499__1437 (.L_HI(net1437));
 sg13g2_tiehi _34294__1438 (.L_HI(net1438));
 sg13g2_tiehi _36066__1439 (.L_HI(net1439));
 sg13g2_tiehi _34293__1440 (.L_HI(net1440));
 sg13g2_tiehi _35498__1441 (.L_HI(net1441));
 sg13g2_tiehi _34292__1442 (.L_HI(net1442));
 sg13g2_tiehi _36065__1443 (.L_HI(net1443));
 sg13g2_tiehi _34291__1444 (.L_HI(net1444));
 sg13g2_tiehi _35497__1445 (.L_HI(net1445));
 sg13g2_tiehi _34290__1446 (.L_HI(net1446));
 sg13g2_tiehi _36064__1447 (.L_HI(net1447));
 sg13g2_tiehi _34289__1448 (.L_HI(net1448));
 sg13g2_tiehi _35496__1449 (.L_HI(net1449));
 sg13g2_tiehi _34288__1450 (.L_HI(net1450));
 sg13g2_tiehi _36063__1451 (.L_HI(net1451));
 sg13g2_tiehi _34287__1452 (.L_HI(net1452));
 sg13g2_tiehi _35495__1453 (.L_HI(net1453));
 sg13g2_tiehi _34286__1454 (.L_HI(net1454));
 sg13g2_tiehi _36062__1455 (.L_HI(net1455));
 sg13g2_tiehi _34285__1456 (.L_HI(net1456));
 sg13g2_tiehi _35494__1457 (.L_HI(net1457));
 sg13g2_tiehi _34284__1458 (.L_HI(net1458));
 sg13g2_tiehi _36061__1459 (.L_HI(net1459));
 sg13g2_tiehi _34283__1460 (.L_HI(net1460));
 sg13g2_tiehi _35493__1461 (.L_HI(net1461));
 sg13g2_tiehi _34282__1462 (.L_HI(net1462));
 sg13g2_tiehi _36060__1463 (.L_HI(net1463));
 sg13g2_tiehi _34281__1464 (.L_HI(net1464));
 sg13g2_tiehi _35492__1465 (.L_HI(net1465));
 sg13g2_tiehi _34280__1466 (.L_HI(net1466));
 sg13g2_tiehi _36059__1467 (.L_HI(net1467));
 sg13g2_tiehi _34279__1468 (.L_HI(net1468));
 sg13g2_tiehi _35491__1469 (.L_HI(net1469));
 sg13g2_tiehi _34278__1470 (.L_HI(net1470));
 sg13g2_tiehi _36058__1471 (.L_HI(net1471));
 sg13g2_tiehi _34277__1472 (.L_HI(net1472));
 sg13g2_tiehi _35490__1473 (.L_HI(net1473));
 sg13g2_tiehi _34276__1474 (.L_HI(net1474));
 sg13g2_tiehi _36057__1475 (.L_HI(net1475));
 sg13g2_tiehi _34275__1476 (.L_HI(net1476));
 sg13g2_tiehi _35489__1477 (.L_HI(net1477));
 sg13g2_tiehi _34274__1478 (.L_HI(net1478));
 sg13g2_tiehi _36056__1479 (.L_HI(net1479));
 sg13g2_tiehi _34273__1480 (.L_HI(net1480));
 sg13g2_tiehi _35488__1481 (.L_HI(net1481));
 sg13g2_tiehi _34272__1482 (.L_HI(net1482));
 sg13g2_tiehi _36055__1483 (.L_HI(net1483));
 sg13g2_tiehi _34271__1484 (.L_HI(net1484));
 sg13g2_tiehi _35487__1485 (.L_HI(net1485));
 sg13g2_tiehi _34270__1486 (.L_HI(net1486));
 sg13g2_tiehi _36054__1487 (.L_HI(net1487));
 sg13g2_tiehi _34269__1488 (.L_HI(net1488));
 sg13g2_tiehi _35486__1489 (.L_HI(net1489));
 sg13g2_tiehi _34268__1490 (.L_HI(net1490));
 sg13g2_tiehi _36053__1491 (.L_HI(net1491));
 sg13g2_tiehi _34267__1492 (.L_HI(net1492));
 sg13g2_tiehi _35485__1493 (.L_HI(net1493));
 sg13g2_tiehi _34266__1494 (.L_HI(net1494));
 sg13g2_tiehi _36052__1495 (.L_HI(net1495));
 sg13g2_tiehi _34265__1496 (.L_HI(net1496));
 sg13g2_tiehi _35484__1497 (.L_HI(net1497));
 sg13g2_tiehi _34264__1498 (.L_HI(net1498));
 sg13g2_tiehi _36051__1499 (.L_HI(net1499));
 sg13g2_tiehi _34263__1500 (.L_HI(net1500));
 sg13g2_tiehi _35483__1501 (.L_HI(net1501));
 sg13g2_tiehi _34262__1502 (.L_HI(net1502));
 sg13g2_tiehi _36050__1503 (.L_HI(net1503));
 sg13g2_tiehi _34261__1504 (.L_HI(net1504));
 sg13g2_tiehi _35482__1505 (.L_HI(net1505));
 sg13g2_tiehi _34260__1506 (.L_HI(net1506));
 sg13g2_tiehi _36049__1507 (.L_HI(net1507));
 sg13g2_tiehi _34259__1508 (.L_HI(net1508));
 sg13g2_tiehi _35481__1509 (.L_HI(net1509));
 sg13g2_tiehi _34258__1510 (.L_HI(net1510));
 sg13g2_tiehi _36048__1511 (.L_HI(net1511));
 sg13g2_tiehi _34257__1512 (.L_HI(net1512));
 sg13g2_tiehi _35480__1513 (.L_HI(net1513));
 sg13g2_tiehi _34256__1514 (.L_HI(net1514));
 sg13g2_tiehi _36047__1515 (.L_HI(net1515));
 sg13g2_tiehi _34255__1516 (.L_HI(net1516));
 sg13g2_tiehi _35479__1517 (.L_HI(net1517));
 sg13g2_tiehi _34254__1518 (.L_HI(net1518));
 sg13g2_tiehi _36046__1519 (.L_HI(net1519));
 sg13g2_tiehi _34253__1520 (.L_HI(net1520));
 sg13g2_tiehi _35478__1521 (.L_HI(net1521));
 sg13g2_tiehi _34252__1522 (.L_HI(net1522));
 sg13g2_tiehi _36045__1523 (.L_HI(net1523));
 sg13g2_tiehi _34251__1524 (.L_HI(net1524));
 sg13g2_tiehi _35477__1525 (.L_HI(net1525));
 sg13g2_tiehi _34250__1526 (.L_HI(net1526));
 sg13g2_tiehi _36044__1527 (.L_HI(net1527));
 sg13g2_tiehi _34249__1528 (.L_HI(net1528));
 sg13g2_tiehi _35476__1529 (.L_HI(net1529));
 sg13g2_tiehi _34248__1530 (.L_HI(net1530));
 sg13g2_tiehi _36043__1531 (.L_HI(net1531));
 sg13g2_tiehi _34247__1532 (.L_HI(net1532));
 sg13g2_tiehi _35475__1533 (.L_HI(net1533));
 sg13g2_tiehi _34246__1534 (.L_HI(net1534));
 sg13g2_tiehi _36042__1535 (.L_HI(net1535));
 sg13g2_tiehi _34245__1536 (.L_HI(net1536));
 sg13g2_tiehi _35474__1537 (.L_HI(net1537));
 sg13g2_tiehi _34244__1538 (.L_HI(net1538));
 sg13g2_tiehi _35473__1539 (.L_HI(net1539));
 sg13g2_tiehi _34243__1540 (.L_HI(net1540));
 sg13g2_tiehi _36041__1541 (.L_HI(net1541));
 sg13g2_tiehi _34242__1542 (.L_HI(net1542));
 sg13g2_tiehi _35472__1543 (.L_HI(net1543));
 sg13g2_tiehi _34241__1544 (.L_HI(net1544));
 sg13g2_tiehi _36040__1545 (.L_HI(net1545));
 sg13g2_tiehi _34240__1546 (.L_HI(net1546));
 sg13g2_tiehi _35471__1547 (.L_HI(net1547));
 sg13g2_tiehi _34239__1548 (.L_HI(net1548));
 sg13g2_tiehi _36039__1549 (.L_HI(net1549));
 sg13g2_tiehi _34238__1550 (.L_HI(net1550));
 sg13g2_tiehi _35470__1551 (.L_HI(net1551));
 sg13g2_tiehi _34237__1552 (.L_HI(net1552));
 sg13g2_tiehi _36038__1553 (.L_HI(net1553));
 sg13g2_tiehi _34236__1554 (.L_HI(net1554));
 sg13g2_tiehi _35469__1555 (.L_HI(net1555));
 sg13g2_tiehi _34235__1556 (.L_HI(net1556));
 sg13g2_tiehi _36037__1557 (.L_HI(net1557));
 sg13g2_tiehi _34234__1558 (.L_HI(net1558));
 sg13g2_tiehi _35468__1559 (.L_HI(net1559));
 sg13g2_tiehi _34233__1560 (.L_HI(net1560));
 sg13g2_tiehi _36036__1561 (.L_HI(net1561));
 sg13g2_tiehi _34232__1562 (.L_HI(net1562));
 sg13g2_tiehi _35467__1563 (.L_HI(net1563));
 sg13g2_tiehi _34231__1564 (.L_HI(net1564));
 sg13g2_tiehi _36035__1565 (.L_HI(net1565));
 sg13g2_tiehi _34230__1566 (.L_HI(net1566));
 sg13g2_tiehi _35466__1567 (.L_HI(net1567));
 sg13g2_tiehi _34229__1568 (.L_HI(net1568));
 sg13g2_tiehi _36034__1569 (.L_HI(net1569));
 sg13g2_tiehi _34228__1570 (.L_HI(net1570));
 sg13g2_tiehi _35465__1571 (.L_HI(net1571));
 sg13g2_tiehi _34227__1572 (.L_HI(net1572));
 sg13g2_tiehi _36033__1573 (.L_HI(net1573));
 sg13g2_tiehi _34226__1574 (.L_HI(net1574));
 sg13g2_tiehi _35464__1575 (.L_HI(net1575));
 sg13g2_tiehi _34225__1576 (.L_HI(net1576));
 sg13g2_tiehi _36032__1577 (.L_HI(net1577));
 sg13g2_tiehi _34224__1578 (.L_HI(net1578));
 sg13g2_tiehi _35463__1579 (.L_HI(net1579));
 sg13g2_tiehi _34223__1580 (.L_HI(net1580));
 sg13g2_tiehi _36031__1581 (.L_HI(net1581));
 sg13g2_tiehi _34222__1582 (.L_HI(net1582));
 sg13g2_tiehi _35462__1583 (.L_HI(net1583));
 sg13g2_tiehi _34221__1584 (.L_HI(net1584));
 sg13g2_tiehi _36030__1585 (.L_HI(net1585));
 sg13g2_tiehi _34220__1586 (.L_HI(net1586));
 sg13g2_tiehi _35461__1587 (.L_HI(net1587));
 sg13g2_tiehi _34219__1588 (.L_HI(net1588));
 sg13g2_tiehi _36029__1589 (.L_HI(net1589));
 sg13g2_tiehi _34218__1590 (.L_HI(net1590));
 sg13g2_tiehi _35460__1591 (.L_HI(net1591));
 sg13g2_tiehi _34217__1592 (.L_HI(net1592));
 sg13g2_tiehi _36028__1593 (.L_HI(net1593));
 sg13g2_tiehi _34216__1594 (.L_HI(net1594));
 sg13g2_tiehi _35459__1595 (.L_HI(net1595));
 sg13g2_tiehi _34215__1596 (.L_HI(net1596));
 sg13g2_tiehi _36027__1597 (.L_HI(net1597));
 sg13g2_tiehi _34214__1598 (.L_HI(net1598));
 sg13g2_tiehi _35458__1599 (.L_HI(net1599));
 sg13g2_tiehi _34213__1600 (.L_HI(net1600));
 sg13g2_tiehi _36026__1601 (.L_HI(net1601));
 sg13g2_tiehi _34212__1602 (.L_HI(net1602));
 sg13g2_tiehi _35457__1603 (.L_HI(net1603));
 sg13g2_tiehi _34211__1604 (.L_HI(net1604));
 sg13g2_tiehi _36025__1605 (.L_HI(net1605));
 sg13g2_tiehi _34210__1606 (.L_HI(net1606));
 sg13g2_tiehi _35456__1607 (.L_HI(net1607));
 sg13g2_tiehi _34209__1608 (.L_HI(net1608));
 sg13g2_tiehi _36024__1609 (.L_HI(net1609));
 sg13g2_tiehi _34208__1610 (.L_HI(net1610));
 sg13g2_tiehi _35455__1611 (.L_HI(net1611));
 sg13g2_tiehi _34207__1612 (.L_HI(net1612));
 sg13g2_tiehi _36023__1613 (.L_HI(net1613));
 sg13g2_tiehi _34206__1614 (.L_HI(net1614));
 sg13g2_tiehi _35454__1615 (.L_HI(net1615));
 sg13g2_tiehi _34205__1616 (.L_HI(net1616));
 sg13g2_tiehi _36022__1617 (.L_HI(net1617));
 sg13g2_tiehi _34204__1618 (.L_HI(net1618));
 sg13g2_tiehi _35453__1619 (.L_HI(net1619));
 sg13g2_tiehi _34203__1620 (.L_HI(net1620));
 sg13g2_tiehi _36021__1621 (.L_HI(net1621));
 sg13g2_tiehi _34202__1622 (.L_HI(net1622));
 sg13g2_tiehi _35452__1623 (.L_HI(net1623));
 sg13g2_tiehi _34201__1624 (.L_HI(net1624));
 sg13g2_tiehi _36020__1625 (.L_HI(net1625));
 sg13g2_tiehi _34200__1626 (.L_HI(net1626));
 sg13g2_tiehi _35451__1627 (.L_HI(net1627));
 sg13g2_tiehi _34199__1628 (.L_HI(net1628));
 sg13g2_tiehi _36019__1629 (.L_HI(net1629));
 sg13g2_tiehi _34198__1630 (.L_HI(net1630));
 sg13g2_tiehi _35450__1631 (.L_HI(net1631));
 sg13g2_tiehi _34197__1632 (.L_HI(net1632));
 sg13g2_tiehi _36018__1633 (.L_HI(net1633));
 sg13g2_tiehi _34196__1634 (.L_HI(net1634));
 sg13g2_tiehi _35449__1635 (.L_HI(net1635));
 sg13g2_tiehi _34195__1636 (.L_HI(net1636));
 sg13g2_tiehi _36017__1637 (.L_HI(net1637));
 sg13g2_tiehi _34194__1638 (.L_HI(net1638));
 sg13g2_tiehi _35448__1639 (.L_HI(net1639));
 sg13g2_tiehi _34193__1640 (.L_HI(net1640));
 sg13g2_tiehi _36016__1641 (.L_HI(net1641));
 sg13g2_tiehi _34192__1642 (.L_HI(net1642));
 sg13g2_tiehi _35447__1643 (.L_HI(net1643));
 sg13g2_tiehi _34191__1644 (.L_HI(net1644));
 sg13g2_tiehi _36015__1645 (.L_HI(net1645));
 sg13g2_tiehi _34190__1646 (.L_HI(net1646));
 sg13g2_tiehi _35446__1647 (.L_HI(net1647));
 sg13g2_tiehi _34189__1648 (.L_HI(net1648));
 sg13g2_tiehi _36014__1649 (.L_HI(net1649));
 sg13g2_tiehi _34188__1650 (.L_HI(net1650));
 sg13g2_tiehi _35445__1651 (.L_HI(net1651));
 sg13g2_tiehi _34187__1652 (.L_HI(net1652));
 sg13g2_tiehi _36013__1653 (.L_HI(net1653));
 sg13g2_tiehi _34186__1654 (.L_HI(net1654));
 sg13g2_tiehi _35444__1655 (.L_HI(net1655));
 sg13g2_tiehi _34185__1656 (.L_HI(net1656));
 sg13g2_tiehi _36012__1657 (.L_HI(net1657));
 sg13g2_tiehi _34184__1658 (.L_HI(net1658));
 sg13g2_tiehi _35443__1659 (.L_HI(net1659));
 sg13g2_tiehi _34183__1660 (.L_HI(net1660));
 sg13g2_tiehi _36011__1661 (.L_HI(net1661));
 sg13g2_tiehi _34182__1662 (.L_HI(net1662));
 sg13g2_tiehi _35442__1663 (.L_HI(net1663));
 sg13g2_tiehi _34181__1664 (.L_HI(net1664));
 sg13g2_tiehi _36010__1665 (.L_HI(net1665));
 sg13g2_tiehi _34180__1666 (.L_HI(net1666));
 sg13g2_tiehi _35441__1667 (.L_HI(net1667));
 sg13g2_tiehi _34179__1668 (.L_HI(net1668));
 sg13g2_tiehi _35440__1669 (.L_HI(net1669));
 sg13g2_tiehi _34178__1670 (.L_HI(net1670));
 sg13g2_tiehi _35439__1671 (.L_HI(net1671));
 sg13g2_tiehi _34177__1672 (.L_HI(net1672));
 sg13g2_tiehi _36009__1673 (.L_HI(net1673));
 sg13g2_tiehi _34176__1674 (.L_HI(net1674));
 sg13g2_tiehi _35438__1675 (.L_HI(net1675));
 sg13g2_tiehi _34175__1676 (.L_HI(net1676));
 sg13g2_tiehi _36008__1677 (.L_HI(net1677));
 sg13g2_tiehi _34174__1678 (.L_HI(net1678));
 sg13g2_tiehi _35437__1679 (.L_HI(net1679));
 sg13g2_tiehi _34173__1680 (.L_HI(net1680));
 sg13g2_tiehi _36007__1681 (.L_HI(net1681));
 sg13g2_tiehi _34172__1682 (.L_HI(net1682));
 sg13g2_tiehi _35436__1683 (.L_HI(net1683));
 sg13g2_tiehi _34171__1684 (.L_HI(net1684));
 sg13g2_tiehi _36006__1685 (.L_HI(net1685));
 sg13g2_tiehi _34170__1686 (.L_HI(net1686));
 sg13g2_tiehi _35435__1687 (.L_HI(net1687));
 sg13g2_tiehi _34169__1688 (.L_HI(net1688));
 sg13g2_tiehi _36005__1689 (.L_HI(net1689));
 sg13g2_tiehi _34168__1690 (.L_HI(net1690));
 sg13g2_tiehi _35434__1691 (.L_HI(net1691));
 sg13g2_tiehi _34167__1692 (.L_HI(net1692));
 sg13g2_tiehi _36004__1693 (.L_HI(net1693));
 sg13g2_tiehi _34166__1694 (.L_HI(net1694));
 sg13g2_tiehi _35433__1695 (.L_HI(net1695));
 sg13g2_tiehi _34165__1696 (.L_HI(net1696));
 sg13g2_tiehi _36003__1697 (.L_HI(net1697));
 sg13g2_tiehi _34164__1698 (.L_HI(net1698));
 sg13g2_tiehi _35432__1699 (.L_HI(net1699));
 sg13g2_tiehi _34163__1700 (.L_HI(net1700));
 sg13g2_tiehi _36002__1701 (.L_HI(net1701));
 sg13g2_tiehi _34162__1702 (.L_HI(net1702));
 sg13g2_tiehi _35431__1703 (.L_HI(net1703));
 sg13g2_tiehi _34161__1704 (.L_HI(net1704));
 sg13g2_tiehi _36001__1705 (.L_HI(net1705));
 sg13g2_tiehi _34160__1706 (.L_HI(net1706));
 sg13g2_tiehi _35430__1707 (.L_HI(net1707));
 sg13g2_tiehi _34159__1708 (.L_HI(net1708));
 sg13g2_tiehi _36000__1709 (.L_HI(net1709));
 sg13g2_tiehi _34158__1710 (.L_HI(net1710));
 sg13g2_tiehi _35429__1711 (.L_HI(net1711));
 sg13g2_tiehi _34157__1712 (.L_HI(net1712));
 sg13g2_tiehi _35999__1713 (.L_HI(net1713));
 sg13g2_tiehi _34156__1714 (.L_HI(net1714));
 sg13g2_tiehi _35428__1715 (.L_HI(net1715));
 sg13g2_tiehi _34155__1716 (.L_HI(net1716));
 sg13g2_tiehi _35998__1717 (.L_HI(net1717));
 sg13g2_tiehi _34154__1718 (.L_HI(net1718));
 sg13g2_tiehi _35427__1719 (.L_HI(net1719));
 sg13g2_tiehi _34153__1720 (.L_HI(net1720));
 sg13g2_tiehi _35997__1721 (.L_HI(net1721));
 sg13g2_tiehi _34152__1722 (.L_HI(net1722));
 sg13g2_tiehi _35426__1723 (.L_HI(net1723));
 sg13g2_tiehi _34151__1724 (.L_HI(net1724));
 sg13g2_tiehi _35996__1725 (.L_HI(net1725));
 sg13g2_tiehi _34150__1726 (.L_HI(net1726));
 sg13g2_tiehi _34149__1727 (.L_HI(net1727));
 sg13g2_tiehi _34148__1728 (.L_HI(net1728));
 sg13g2_tiehi _34147__1729 (.L_HI(net1729));
 sg13g2_tiehi _34146__1730 (.L_HI(net1730));
 sg13g2_tiehi _34145__1731 (.L_HI(net1731));
 sg13g2_tiehi _34144__1732 (.L_HI(net1732));
 sg13g2_tiehi _34143__1733 (.L_HI(net1733));
 sg13g2_tiehi _34142__1734 (.L_HI(net1734));
 sg13g2_tiehi _34141__1735 (.L_HI(net1735));
 sg13g2_tiehi _34140__1736 (.L_HI(net1736));
 sg13g2_tiehi _34139__1737 (.L_HI(net1737));
 sg13g2_tiehi _34138__1738 (.L_HI(net1738));
 sg13g2_tiehi _34137__1739 (.L_HI(net1739));
 sg13g2_tiehi _34136__1740 (.L_HI(net1740));
 sg13g2_tiehi _34135__1741 (.L_HI(net1741));
 sg13g2_tiehi _34134__1742 (.L_HI(net1742));
 sg13g2_tiehi _34133__1743 (.L_HI(net1743));
 sg13g2_tiehi _34132__1744 (.L_HI(net1744));
 sg13g2_tiehi _34131__1745 (.L_HI(net1745));
 sg13g2_tiehi _34130__1746 (.L_HI(net1746));
 sg13g2_tiehi _34129__1747 (.L_HI(net1747));
 sg13g2_tiehi _34128__1748 (.L_HI(net1748));
 sg13g2_tiehi _34127__1749 (.L_HI(net1749));
 sg13g2_tiehi _34126__1750 (.L_HI(net1750));
 sg13g2_tiehi _34125__1751 (.L_HI(net1751));
 sg13g2_tiehi _34124__1752 (.L_HI(net1752));
 sg13g2_tiehi _34123__1753 (.L_HI(net1753));
 sg13g2_tiehi _34122__1754 (.L_HI(net1754));
 sg13g2_tiehi _34121__1755 (.L_HI(net1755));
 sg13g2_tiehi _34120__1756 (.L_HI(net1756));
 sg13g2_tiehi _34119__1757 (.L_HI(net1757));
 sg13g2_tiehi _34118__1758 (.L_HI(net1758));
 sg13g2_tiehi _34117__1759 (.L_HI(net1759));
 sg13g2_tiehi _34116__1760 (.L_HI(net1760));
 sg13g2_tiehi _34115__1761 (.L_HI(net1761));
 sg13g2_tiehi _34114__1762 (.L_HI(net1762));
 sg13g2_tiehi _34113__1763 (.L_HI(net1763));
 sg13g2_tiehi _34112__1764 (.L_HI(net1764));
 sg13g2_tiehi _34111__1765 (.L_HI(net1765));
 sg13g2_tiehi _34110__1766 (.L_HI(net1766));
 sg13g2_tiehi _34109__1767 (.L_HI(net1767));
 sg13g2_tiehi _34108__1768 (.L_HI(net1768));
 sg13g2_tiehi _34107__1769 (.L_HI(net1769));
 sg13g2_tiehi _34106__1770 (.L_HI(net1770));
 sg13g2_tiehi _34105__1771 (.L_HI(net1771));
 sg13g2_tiehi _34104__1772 (.L_HI(net1772));
 sg13g2_tiehi _34103__1773 (.L_HI(net1773));
 sg13g2_tiehi _34102__1774 (.L_HI(net1774));
 sg13g2_tiehi _34101__1775 (.L_HI(net1775));
 sg13g2_tiehi _34100__1776 (.L_HI(net1776));
 sg13g2_tiehi _34099__1777 (.L_HI(net1777));
 sg13g2_tiehi _34098__1778 (.L_HI(net1778));
 sg13g2_tiehi _34097__1779 (.L_HI(net1779));
 sg13g2_tiehi _34096__1780 (.L_HI(net1780));
 sg13g2_tiehi _34095__1781 (.L_HI(net1781));
 sg13g2_tiehi _34094__1782 (.L_HI(net1782));
 sg13g2_tiehi _34093__1783 (.L_HI(net1783));
 sg13g2_tiehi _34092__1784 (.L_HI(net1784));
 sg13g2_tiehi _34091__1785 (.L_HI(net1785));
 sg13g2_tiehi _34090__1786 (.L_HI(net1786));
 sg13g2_tiehi _34089__1787 (.L_HI(net1787));
 sg13g2_tiehi _34088__1788 (.L_HI(net1788));
 sg13g2_tiehi _34087__1789 (.L_HI(net1789));
 sg13g2_tiehi _34086__1790 (.L_HI(net1790));
 sg13g2_tiehi _35425__1791 (.L_HI(net1791));
 sg13g2_tiehi _34085__1792 (.L_HI(net1792));
 sg13g2_tiehi _35424__1793 (.L_HI(net1793));
 sg13g2_tiehi _34084__1794 (.L_HI(net1794));
 sg13g2_tiehi _34083__1795 (.L_HI(net1795));
 sg13g2_tiehi _34082__1796 (.L_HI(net1796));
 sg13g2_tiehi _34081__1797 (.L_HI(net1797));
 sg13g2_tiehi _34080__1798 (.L_HI(net1798));
 sg13g2_tiehi _34079__1799 (.L_HI(net1799));
 sg13g2_tiehi _34078__1800 (.L_HI(net1800));
 sg13g2_tiehi _34077__1801 (.L_HI(net1801));
 sg13g2_tiehi _34076__1802 (.L_HI(net1802));
 sg13g2_tiehi _34075__1803 (.L_HI(net1803));
 sg13g2_tiehi _34074__1804 (.L_HI(net1804));
 sg13g2_tiehi _34073__1805 (.L_HI(net1805));
 sg13g2_tiehi _34072__1806 (.L_HI(net1806));
 sg13g2_tiehi _34071__1807 (.L_HI(net1807));
 sg13g2_tiehi _34070__1808 (.L_HI(net1808));
 sg13g2_tiehi _34069__1809 (.L_HI(net1809));
 sg13g2_tiehi _34068__1810 (.L_HI(net1810));
 sg13g2_tiehi _34067__1811 (.L_HI(net1811));
 sg13g2_tiehi _34066__1812 (.L_HI(net1812));
 sg13g2_tiehi _34065__1813 (.L_HI(net1813));
 sg13g2_tiehi _34064__1814 (.L_HI(net1814));
 sg13g2_tiehi _34063__1815 (.L_HI(net1815));
 sg13g2_tiehi _34062__1816 (.L_HI(net1816));
 sg13g2_tiehi _34061__1817 (.L_HI(net1817));
 sg13g2_tiehi _34060__1818 (.L_HI(net1818));
 sg13g2_tiehi _34059__1819 (.L_HI(net1819));
 sg13g2_tiehi _34058__1820 (.L_HI(net1820));
 sg13g2_tiehi _34057__1821 (.L_HI(net1821));
 sg13g2_tiehi _34056__1822 (.L_HI(net1822));
 sg13g2_tiehi _34055__1823 (.L_HI(net1823));
 sg13g2_tiehi _34054__1824 (.L_HI(net1824));
 sg13g2_tiehi _34053__1825 (.L_HI(net1825));
 sg13g2_tiehi _34052__1826 (.L_HI(net1826));
 sg13g2_tiehi _34051__1827 (.L_HI(net1827));
 sg13g2_tiehi _34050__1828 (.L_HI(net1828));
 sg13g2_tiehi _34049__1829 (.L_HI(net1829));
 sg13g2_tiehi _34048__1830 (.L_HI(net1830));
 sg13g2_tiehi _34047__1831 (.L_HI(net1831));
 sg13g2_tiehi _34046__1832 (.L_HI(net1832));
 sg13g2_tiehi _34045__1833 (.L_HI(net1833));
 sg13g2_tiehi _34044__1834 (.L_HI(net1834));
 sg13g2_tiehi _34043__1835 (.L_HI(net1835));
 sg13g2_tiehi _34042__1836 (.L_HI(net1836));
 sg13g2_tiehi _34041__1837 (.L_HI(net1837));
 sg13g2_tiehi _34040__1838 (.L_HI(net1838));
 sg13g2_tiehi _34039__1839 (.L_HI(net1839));
 sg13g2_tiehi _34038__1840 (.L_HI(net1840));
 sg13g2_tiehi _34037__1841 (.L_HI(net1841));
 sg13g2_tiehi _34036__1842 (.L_HI(net1842));
 sg13g2_tiehi _34035__1843 (.L_HI(net1843));
 sg13g2_tiehi _34034__1844 (.L_HI(net1844));
 sg13g2_tiehi _34033__1845 (.L_HI(net1845));
 sg13g2_tiehi _34032__1846 (.L_HI(net1846));
 sg13g2_tiehi _34031__1847 (.L_HI(net1847));
 sg13g2_tiehi _34030__1848 (.L_HI(net1848));
 sg13g2_tiehi _34029__1849 (.L_HI(net1849));
 sg13g2_tiehi _34028__1850 (.L_HI(net1850));
 sg13g2_tiehi _34027__1851 (.L_HI(net1851));
 sg13g2_tiehi _34026__1852 (.L_HI(net1852));
 sg13g2_tiehi _34025__1853 (.L_HI(net1853));
 sg13g2_tiehi _34024__1854 (.L_HI(net1854));
 sg13g2_tiehi _34023__1855 (.L_HI(net1855));
 sg13g2_tiehi _34022__1856 (.L_HI(net1856));
 sg13g2_tiehi _34021__1857 (.L_HI(net1857));
 sg13g2_tiehi _34020__1858 (.L_HI(net1858));
 sg13g2_tiehi _34019__1859 (.L_HI(net1859));
 sg13g2_tiehi _34018__1860 (.L_HI(net1860));
 sg13g2_tiehi _34017__1861 (.L_HI(net1861));
 sg13g2_tiehi _34016__1862 (.L_HI(net1862));
 sg13g2_tiehi _34015__1863 (.L_HI(net1863));
 sg13g2_tiehi _34014__1864 (.L_HI(net1864));
 sg13g2_tiehi _34013__1865 (.L_HI(net1865));
 sg13g2_tiehi _34012__1866 (.L_HI(net1866));
 sg13g2_tiehi _34011__1867 (.L_HI(net1867));
 sg13g2_tiehi _34010__1868 (.L_HI(net1868));
 sg13g2_tiehi _34009__1869 (.L_HI(net1869));
 sg13g2_tiehi _34008__1870 (.L_HI(net1870));
 sg13g2_tiehi _34007__1871 (.L_HI(net1871));
 sg13g2_tiehi _34006__1872 (.L_HI(net1872));
 sg13g2_tiehi _34005__1873 (.L_HI(net1873));
 sg13g2_tiehi _34004__1874 (.L_HI(net1874));
 sg13g2_tiehi _34003__1875 (.L_HI(net1875));
 sg13g2_tiehi _34002__1876 (.L_HI(net1876));
 sg13g2_tiehi _34001__1877 (.L_HI(net1877));
 sg13g2_tiehi _34000__1878 (.L_HI(net1878));
 sg13g2_tiehi _33999__1879 (.L_HI(net1879));
 sg13g2_tiehi _33998__1880 (.L_HI(net1880));
 sg13g2_tiehi _33997__1881 (.L_HI(net1881));
 sg13g2_tiehi _33996__1882 (.L_HI(net1882));
 sg13g2_tiehi _33995__1883 (.L_HI(net1883));
 sg13g2_tiehi _33994__1884 (.L_HI(net1884));
 sg13g2_tiehi _33993__1885 (.L_HI(net1885));
 sg13g2_tiehi _33992__1886 (.L_HI(net1886));
 sg13g2_tiehi _33991__1887 (.L_HI(net1887));
 sg13g2_tiehi _33990__1888 (.L_HI(net1888));
 sg13g2_tiehi _33989__1889 (.L_HI(net1889));
 sg13g2_tiehi _33988__1890 (.L_HI(net1890));
 sg13g2_tiehi _33987__1891 (.L_HI(net1891));
 sg13g2_tiehi _33986__1892 (.L_HI(net1892));
 sg13g2_tiehi _33985__1893 (.L_HI(net1893));
 sg13g2_tiehi _33984__1894 (.L_HI(net1894));
 sg13g2_tiehi _33983__1895 (.L_HI(net1895));
 sg13g2_tiehi _33982__1896 (.L_HI(net1896));
 sg13g2_tiehi _33981__1897 (.L_HI(net1897));
 sg13g2_tiehi _33980__1898 (.L_HI(net1898));
 sg13g2_tiehi _33979__1899 (.L_HI(net1899));
 sg13g2_tiehi _33978__1900 (.L_HI(net1900));
 sg13g2_tiehi _33977__1901 (.L_HI(net1901));
 sg13g2_tiehi _33976__1902 (.L_HI(net1902));
 sg13g2_tiehi _33975__1903 (.L_HI(net1903));
 sg13g2_tiehi _33974__1904 (.L_HI(net1904));
 sg13g2_tiehi _33973__1905 (.L_HI(net1905));
 sg13g2_tiehi _33972__1906 (.L_HI(net1906));
 sg13g2_tiehi _33971__1907 (.L_HI(net1907));
 sg13g2_tiehi _33970__1908 (.L_HI(net1908));
 sg13g2_tiehi _33969__1909 (.L_HI(net1909));
 sg13g2_tiehi _33968__1910 (.L_HI(net1910));
 sg13g2_tiehi _33967__1911 (.L_HI(net1911));
 sg13g2_tiehi _33966__1912 (.L_HI(net1912));
 sg13g2_tiehi _33965__1913 (.L_HI(net1913));
 sg13g2_tiehi _33964__1914 (.L_HI(net1914));
 sg13g2_tiehi _33963__1915 (.L_HI(net1915));
 sg13g2_tiehi _33962__1916 (.L_HI(net1916));
 sg13g2_tiehi _33961__1917 (.L_HI(net1917));
 sg13g2_tiehi _33960__1918 (.L_HI(net1918));
 sg13g2_tiehi _33959__1919 (.L_HI(net1919));
 sg13g2_tiehi _33958__1920 (.L_HI(net1920));
 sg13g2_tiehi _33957__1921 (.L_HI(net1921));
 sg13g2_tiehi _33956__1922 (.L_HI(net1922));
 sg13g2_tiehi _33955__1923 (.L_HI(net1923));
 sg13g2_tiehi _33954__1924 (.L_HI(net1924));
 sg13g2_tiehi _33953__1925 (.L_HI(net1925));
 sg13g2_tiehi _33952__1926 (.L_HI(net1926));
 sg13g2_tiehi _33951__1927 (.L_HI(net1927));
 sg13g2_tiehi _33950__1928 (.L_HI(net1928));
 sg13g2_tiehi _33949__1929 (.L_HI(net1929));
 sg13g2_tiehi _33948__1930 (.L_HI(net1930));
 sg13g2_tiehi _33947__1931 (.L_HI(net1931));
 sg13g2_tiehi _33946__1932 (.L_HI(net1932));
 sg13g2_tiehi _33945__1933 (.L_HI(net1933));
 sg13g2_tiehi _33944__1934 (.L_HI(net1934));
 sg13g2_tiehi _33943__1935 (.L_HI(net1935));
 sg13g2_tiehi _33942__1936 (.L_HI(net1936));
 sg13g2_tiehi _33941__1937 (.L_HI(net1937));
 sg13g2_tiehi _33940__1938 (.L_HI(net1938));
 sg13g2_tiehi _35423__1939 (.L_HI(net1939));
 sg13g2_tiehi _33939__1940 (.L_HI(net1940));
 sg13g2_tiehi _35422__1941 (.L_HI(net1941));
 sg13g2_tiehi _33938__1942 (.L_HI(net1942));
 sg13g2_tiehi _35421__1943 (.L_HI(net1943));
 sg13g2_tiehi _33937__1944 (.L_HI(net1944));
 sg13g2_tiehi _35420__1945 (.L_HI(net1945));
 sg13g2_tiehi _33936__1946 (.L_HI(net1946));
 sg13g2_tiehi _35419__1947 (.L_HI(net1947));
 sg13g2_tiehi _33935__1948 (.L_HI(net1948));
 sg13g2_tiehi _35418__1949 (.L_HI(net1949));
 sg13g2_tiehi _33934__1950 (.L_HI(net1950));
 sg13g2_tiehi _35417__1951 (.L_HI(net1951));
 sg13g2_tiehi _33933__1952 (.L_HI(net1952));
 sg13g2_tiehi _35416__1953 (.L_HI(net1953));
 sg13g2_tiehi _33932__1954 (.L_HI(net1954));
 sg13g2_tiehi _35415__1955 (.L_HI(net1955));
 sg13g2_tiehi _33931__1956 (.L_HI(net1956));
 sg13g2_tiehi _35414__1957 (.L_HI(net1957));
 sg13g2_tiehi _33930__1958 (.L_HI(net1958));
 sg13g2_tiehi _35413__1959 (.L_HI(net1959));
 sg13g2_tiehi _33929__1960 (.L_HI(net1960));
 sg13g2_tiehi _35412__1961 (.L_HI(net1961));
 sg13g2_tiehi _33928__1962 (.L_HI(net1962));
 sg13g2_tiehi _35411__1963 (.L_HI(net1963));
 sg13g2_tiehi _33927__1964 (.L_HI(net1964));
 sg13g2_tiehi _35410__1965 (.L_HI(net1965));
 sg13g2_tiehi _33926__1966 (.L_HI(net1966));
 sg13g2_tiehi _35409__1967 (.L_HI(net1967));
 sg13g2_tiehi _33925__1968 (.L_HI(net1968));
 sg13g2_tiehi _35408__1969 (.L_HI(net1969));
 sg13g2_tiehi _33924__1970 (.L_HI(net1970));
 sg13g2_tiehi _35407__1971 (.L_HI(net1971));
 sg13g2_tiehi _33923__1972 (.L_HI(net1972));
 sg13g2_tiehi _35406__1973 (.L_HI(net1973));
 sg13g2_tiehi _33922__1974 (.L_HI(net1974));
 sg13g2_tiehi _35405__1975 (.L_HI(net1975));
 sg13g2_tiehi _33921__1976 (.L_HI(net1976));
 sg13g2_tiehi _35404__1977 (.L_HI(net1977));
 sg13g2_tiehi _33920__1978 (.L_HI(net1978));
 sg13g2_tiehi _35403__1979 (.L_HI(net1979));
 sg13g2_tiehi _33919__1980 (.L_HI(net1980));
 sg13g2_tiehi _35402__1981 (.L_HI(net1981));
 sg13g2_tiehi _33918__1982 (.L_HI(net1982));
 sg13g2_tiehi _35401__1983 (.L_HI(net1983));
 sg13g2_tiehi _33917__1984 (.L_HI(net1984));
 sg13g2_tiehi _35400__1985 (.L_HI(net1985));
 sg13g2_tiehi _33916__1986 (.L_HI(net1986));
 sg13g2_tiehi _35399__1987 (.L_HI(net1987));
 sg13g2_tiehi _33915__1988 (.L_HI(net1988));
 sg13g2_tiehi _35398__1989 (.L_HI(net1989));
 sg13g2_tiehi _33914__1990 (.L_HI(net1990));
 sg13g2_tiehi _35397__1991 (.L_HI(net1991));
 sg13g2_tiehi _33913__1992 (.L_HI(net1992));
 sg13g2_tiehi _35396__1993 (.L_HI(net1993));
 sg13g2_tiehi _33912__1994 (.L_HI(net1994));
 sg13g2_tiehi _35395__1995 (.L_HI(net1995));
 sg13g2_tiehi _33911__1996 (.L_HI(net1996));
 sg13g2_tiehi _35394__1997 (.L_HI(net1997));
 sg13g2_tiehi _33910__1998 (.L_HI(net1998));
 sg13g2_tiehi _35393__1999 (.L_HI(net1999));
 sg13g2_tiehi _33909__2000 (.L_HI(net2000));
 sg13g2_tiehi _35995__2001 (.L_HI(net2001));
 sg13g2_tiehi _33908__2002 (.L_HI(net2002));
 sg13g2_tiehi _33907__2003 (.L_HI(net2003));
 sg13g2_tiehi _33906__2004 (.L_HI(net2004));
 sg13g2_tiehi _33905__2005 (.L_HI(net2005));
 sg13g2_tiehi _33904__2006 (.L_HI(net2006));
 sg13g2_tiehi _33903__2007 (.L_HI(net2007));
 sg13g2_tiehi _33902__2008 (.L_HI(net2008));
 sg13g2_tiehi _33901__2009 (.L_HI(net2009));
 sg13g2_tiehi _33900__2010 (.L_HI(net2010));
 sg13g2_tiehi _33899__2011 (.L_HI(net2011));
 sg13g2_tiehi _33898__2012 (.L_HI(net2012));
 sg13g2_tiehi _33897__2013 (.L_HI(net2013));
 sg13g2_tiehi _33896__2014 (.L_HI(net2014));
 sg13g2_tiehi _33895__2015 (.L_HI(net2015));
 sg13g2_tiehi _33894__2016 (.L_HI(net2016));
 sg13g2_tiehi _33893__2017 (.L_HI(net2017));
 sg13g2_tiehi _33892__2018 (.L_HI(net2018));
 sg13g2_tiehi _33891__2019 (.L_HI(net2019));
 sg13g2_tiehi _33890__2020 (.L_HI(net2020));
 sg13g2_tiehi _33889__2021 (.L_HI(net2021));
 sg13g2_tiehi _33888__2022 (.L_HI(net2022));
 sg13g2_tiehi _33887__2023 (.L_HI(net2023));
 sg13g2_tiehi _33886__2024 (.L_HI(net2024));
 sg13g2_tiehi _33885__2025 (.L_HI(net2025));
 sg13g2_tiehi _33884__2026 (.L_HI(net2026));
 sg13g2_tiehi _33883__2027 (.L_HI(net2027));
 sg13g2_tiehi _33882__2028 (.L_HI(net2028));
 sg13g2_tiehi _33881__2029 (.L_HI(net2029));
 sg13g2_tiehi _33880__2030 (.L_HI(net2030));
 sg13g2_tiehi _33879__2031 (.L_HI(net2031));
 sg13g2_tiehi _33878__2032 (.L_HI(net2032));
 sg13g2_tiehi _33877__2033 (.L_HI(net2033));
 sg13g2_tiehi _33876__2034 (.L_HI(net2034));
 sg13g2_tiehi _33875__2035 (.L_HI(net2035));
 sg13g2_tiehi _33874__2036 (.L_HI(net2036));
 sg13g2_tiehi _33873__2037 (.L_HI(net2037));
 sg13g2_tiehi _33872__2038 (.L_HI(net2038));
 sg13g2_tiehi _33871__2039 (.L_HI(net2039));
 sg13g2_tiehi _33870__2040 (.L_HI(net2040));
 sg13g2_tiehi _33869__2041 (.L_HI(net2041));
 sg13g2_tiehi _33868__2042 (.L_HI(net2042));
 sg13g2_tiehi _33867__2043 (.L_HI(net2043));
 sg13g2_tiehi _33866__2044 (.L_HI(net2044));
 sg13g2_tiehi _33865__2045 (.L_HI(net2045));
 sg13g2_tiehi _33864__2046 (.L_HI(net2046));
 sg13g2_tiehi _33863__2047 (.L_HI(net2047));
 sg13g2_tiehi _33862__2048 (.L_HI(net2048));
 sg13g2_tiehi _33861__2049 (.L_HI(net2049));
 sg13g2_tiehi _33860__2050 (.L_HI(net2050));
 sg13g2_tiehi _33859__2051 (.L_HI(net2051));
 sg13g2_tiehi _33858__2052 (.L_HI(net2052));
 sg13g2_tiehi _33857__2053 (.L_HI(net2053));
 sg13g2_tiehi _33856__2054 (.L_HI(net2054));
 sg13g2_tiehi _33855__2055 (.L_HI(net2055));
 sg13g2_tiehi _33854__2056 (.L_HI(net2056));
 sg13g2_tiehi _33853__2057 (.L_HI(net2057));
 sg13g2_tiehi _33852__2058 (.L_HI(net2058));
 sg13g2_tiehi _33851__2059 (.L_HI(net2059));
 sg13g2_tiehi _33850__2060 (.L_HI(net2060));
 sg13g2_tiehi _33849__2061 (.L_HI(net2061));
 sg13g2_tiehi _33848__2062 (.L_HI(net2062));
 sg13g2_tiehi _33847__2063 (.L_HI(net2063));
 sg13g2_tiehi _33846__2064 (.L_HI(net2064));
 sg13g2_tiehi _33845__2065 (.L_HI(net2065));
 sg13g2_tiehi _33844__2066 (.L_HI(net2066));
 sg13g2_tiehi _33843__2067 (.L_HI(net2067));
 sg13g2_tiehi _33842__2068 (.L_HI(net2068));
 sg13g2_tiehi _33841__2069 (.L_HI(net2069));
 sg13g2_tiehi _33840__2070 (.L_HI(net2070));
 sg13g2_tiehi _33839__2071 (.L_HI(net2071));
 sg13g2_tiehi _33838__2072 (.L_HI(net2072));
 sg13g2_tiehi _33837__2073 (.L_HI(net2073));
 sg13g2_tiehi _33836__2074 (.L_HI(net2074));
 sg13g2_tiehi _33835__2075 (.L_HI(net2075));
 sg13g2_tiehi _33834__2076 (.L_HI(net2076));
 sg13g2_tiehi _33833__2077 (.L_HI(net2077));
 sg13g2_tiehi _33832__2078 (.L_HI(net2078));
 sg13g2_tiehi _33831__2079 (.L_HI(net2079));
 sg13g2_tiehi _33830__2080 (.L_HI(net2080));
 sg13g2_tiehi _33829__2081 (.L_HI(net2081));
 sg13g2_tiehi _33828__2082 (.L_HI(net2082));
 sg13g2_tiehi _33827__2083 (.L_HI(net2083));
 sg13g2_tiehi _33826__2084 (.L_HI(net2084));
 sg13g2_tiehi _33825__2085 (.L_HI(net2085));
 sg13g2_tiehi _33824__2086 (.L_HI(net2086));
 sg13g2_tiehi _33823__2087 (.L_HI(net2087));
 sg13g2_tiehi _33822__2088 (.L_HI(net2088));
 sg13g2_tiehi _33821__2089 (.L_HI(net2089));
 sg13g2_tiehi _33820__2090 (.L_HI(net2090));
 sg13g2_tiehi _33819__2091 (.L_HI(net2091));
 sg13g2_tiehi _33818__2092 (.L_HI(net2092));
 sg13g2_tiehi _33817__2093 (.L_HI(net2093));
 sg13g2_tiehi _33816__2094 (.L_HI(net2094));
 sg13g2_tiehi _33815__2095 (.L_HI(net2095));
 sg13g2_tiehi _33814__2096 (.L_HI(net2096));
 sg13g2_tiehi _33813__2097 (.L_HI(net2097));
 sg13g2_tiehi _33812__2098 (.L_HI(net2098));
 sg13g2_tiehi _33811__2099 (.L_HI(net2099));
 sg13g2_tiehi _33810__2100 (.L_HI(net2100));
 sg13g2_tiehi _33809__2101 (.L_HI(net2101));
 sg13g2_tiehi _33808__2102 (.L_HI(net2102));
 sg13g2_tiehi _33807__2103 (.L_HI(net2103));
 sg13g2_tiehi _33806__2104 (.L_HI(net2104));
 sg13g2_tiehi _33805__2105 (.L_HI(net2105));
 sg13g2_tiehi _33804__2106 (.L_HI(net2106));
 sg13g2_tiehi _33803__2107 (.L_HI(net2107));
 sg13g2_tiehi _33802__2108 (.L_HI(net2108));
 sg13g2_tiehi _33801__2109 (.L_HI(net2109));
 sg13g2_tiehi _33800__2110 (.L_HI(net2110));
 sg13g2_tiehi _33799__2111 (.L_HI(net2111));
 sg13g2_tiehi _33798__2112 (.L_HI(net2112));
 sg13g2_tiehi _33797__2113 (.L_HI(net2113));
 sg13g2_tiehi _33796__2114 (.L_HI(net2114));
 sg13g2_tiehi _33795__2115 (.L_HI(net2115));
 sg13g2_tiehi _33794__2116 (.L_HI(net2116));
 sg13g2_tiehi _33793__2117 (.L_HI(net2117));
 sg13g2_tiehi _33792__2118 (.L_HI(net2118));
 sg13g2_tiehi _33791__2119 (.L_HI(net2119));
 sg13g2_tiehi _33790__2120 (.L_HI(net2120));
 sg13g2_tiehi _33789__2121 (.L_HI(net2121));
 sg13g2_tiehi _33788__2122 (.L_HI(net2122));
 sg13g2_tiehi _33787__2123 (.L_HI(net2123));
 sg13g2_tiehi _33786__2124 (.L_HI(net2124));
 sg13g2_tiehi _33785__2125 (.L_HI(net2125));
 sg13g2_tiehi _33784__2126 (.L_HI(net2126));
 sg13g2_tiehi _33783__2127 (.L_HI(net2127));
 sg13g2_tiehi _33782__2128 (.L_HI(net2128));
 sg13g2_tiehi _33781__2129 (.L_HI(net2129));
 sg13g2_tiehi _33780__2130 (.L_HI(net2130));
 sg13g2_tiehi _35392__2131 (.L_HI(net2131));
 sg13g2_tiehi _33779__2132 (.L_HI(net2132));
 sg13g2_tiehi _35994__2133 (.L_HI(net2133));
 sg13g2_tiehi _33778__2134 (.L_HI(net2134));
 sg13g2_tiehi _35391__2135 (.L_HI(net2135));
 sg13g2_tiehi _33777__2136 (.L_HI(net2136));
 sg13g2_tiehi _35993__2137 (.L_HI(net2137));
 sg13g2_tiehi _33776__2138 (.L_HI(net2138));
 sg13g2_tiehi _33775__2139 (.L_HI(net2139));
 sg13g2_tiehi _33774__2140 (.L_HI(net2140));
 sg13g2_tiehi _33773__2141 (.L_HI(net2141));
 sg13g2_tiehi _33772__2142 (.L_HI(net2142));
 sg13g2_tiehi _33771__2143 (.L_HI(net2143));
 sg13g2_tiehi _33770__2144 (.L_HI(net2144));
 sg13g2_tiehi _33769__2145 (.L_HI(net2145));
 sg13g2_tiehi _33768__2146 (.L_HI(net2146));
 sg13g2_tiehi _33767__2147 (.L_HI(net2147));
 sg13g2_tiehi _33766__2148 (.L_HI(net2148));
 sg13g2_tiehi _33765__2149 (.L_HI(net2149));
 sg13g2_tiehi _33764__2150 (.L_HI(net2150));
 sg13g2_tiehi _33763__2151 (.L_HI(net2151));
 sg13g2_tiehi _33762__2152 (.L_HI(net2152));
 sg13g2_tiehi _33761__2153 (.L_HI(net2153));
 sg13g2_tiehi _33760__2154 (.L_HI(net2154));
 sg13g2_tiehi _33759__2155 (.L_HI(net2155));
 sg13g2_tiehi _33758__2156 (.L_HI(net2156));
 sg13g2_tiehi _33757__2157 (.L_HI(net2157));
 sg13g2_tiehi _33756__2158 (.L_HI(net2158));
 sg13g2_tiehi _33755__2159 (.L_HI(net2159));
 sg13g2_tiehi _33754__2160 (.L_HI(net2160));
 sg13g2_tiehi _33753__2161 (.L_HI(net2161));
 sg13g2_tiehi _33752__2162 (.L_HI(net2162));
 sg13g2_tiehi _33751__2163 (.L_HI(net2163));
 sg13g2_tiehi _33750__2164 (.L_HI(net2164));
 sg13g2_tiehi _33749__2165 (.L_HI(net2165));
 sg13g2_tiehi _33748__2166 (.L_HI(net2166));
 sg13g2_tiehi _33747__2167 (.L_HI(net2167));
 sg13g2_tiehi _33746__2168 (.L_HI(net2168));
 sg13g2_tiehi _33745__2169 (.L_HI(net2169));
 sg13g2_tiehi _33744__2170 (.L_HI(net2170));
 sg13g2_tiehi _33743__2171 (.L_HI(net2171));
 sg13g2_tiehi _33742__2172 (.L_HI(net2172));
 sg13g2_tiehi _33741__2173 (.L_HI(net2173));
 sg13g2_tiehi _33740__2174 (.L_HI(net2174));
 sg13g2_tiehi _33739__2175 (.L_HI(net2175));
 sg13g2_tiehi _33738__2176 (.L_HI(net2176));
 sg13g2_tiehi _33737__2177 (.L_HI(net2177));
 sg13g2_tiehi _33736__2178 (.L_HI(net2178));
 sg13g2_tiehi _33735__2179 (.L_HI(net2179));
 sg13g2_tiehi _33734__2180 (.L_HI(net2180));
 sg13g2_tiehi _33733__2181 (.L_HI(net2181));
 sg13g2_tiehi _33732__2182 (.L_HI(net2182));
 sg13g2_tiehi _33731__2183 (.L_HI(net2183));
 sg13g2_tiehi _33730__2184 (.L_HI(net2184));
 sg13g2_tiehi _33729__2185 (.L_HI(net2185));
 sg13g2_tiehi _33728__2186 (.L_HI(net2186));
 sg13g2_tiehi _33727__2187 (.L_HI(net2187));
 sg13g2_tiehi _33726__2188 (.L_HI(net2188));
 sg13g2_tiehi _33725__2189 (.L_HI(net2189));
 sg13g2_tiehi _33724__2190 (.L_HI(net2190));
 sg13g2_tiehi _33723__2191 (.L_HI(net2191));
 sg13g2_tiehi _33722__2192 (.L_HI(net2192));
 sg13g2_tiehi _33721__2193 (.L_HI(net2193));
 sg13g2_tiehi _33720__2194 (.L_HI(net2194));
 sg13g2_tiehi _33719__2195 (.L_HI(net2195));
 sg13g2_tiehi _33718__2196 (.L_HI(net2196));
 sg13g2_tiehi _33717__2197 (.L_HI(net2197));
 sg13g2_tiehi _33716__2198 (.L_HI(net2198));
 sg13g2_tiehi _33715__2199 (.L_HI(net2199));
 sg13g2_tiehi _33714__2200 (.L_HI(net2200));
 sg13g2_tiehi _33713__2201 (.L_HI(net2201));
 sg13g2_tiehi _33712__2202 (.L_HI(net2202));
 sg13g2_tiehi _33711__2203 (.L_HI(net2203));
 sg13g2_tiehi _33710__2204 (.L_HI(net2204));
 sg13g2_tiehi _33709__2205 (.L_HI(net2205));
 sg13g2_tiehi _33708__2206 (.L_HI(net2206));
 sg13g2_tiehi _33707__2207 (.L_HI(net2207));
 sg13g2_tiehi _33706__2208 (.L_HI(net2208));
 sg13g2_tiehi _33705__2209 (.L_HI(net2209));
 sg13g2_tiehi _33704__2210 (.L_HI(net2210));
 sg13g2_tiehi _33703__2211 (.L_HI(net2211));
 sg13g2_tiehi _33702__2212 (.L_HI(net2212));
 sg13g2_tiehi _33701__2213 (.L_HI(net2213));
 sg13g2_tiehi _33700__2214 (.L_HI(net2214));
 sg13g2_tiehi _33699__2215 (.L_HI(net2215));
 sg13g2_tiehi _33698__2216 (.L_HI(net2216));
 sg13g2_tiehi _33697__2217 (.L_HI(net2217));
 sg13g2_tiehi _33696__2218 (.L_HI(net2218));
 sg13g2_tiehi _33695__2219 (.L_HI(net2219));
 sg13g2_tiehi _33694__2220 (.L_HI(net2220));
 sg13g2_tiehi _33693__2221 (.L_HI(net2221));
 sg13g2_tiehi _33692__2222 (.L_HI(net2222));
 sg13g2_tiehi _33691__2223 (.L_HI(net2223));
 sg13g2_tiehi _33690__2224 (.L_HI(net2224));
 sg13g2_tiehi _33689__2225 (.L_HI(net2225));
 sg13g2_tiehi _33688__2226 (.L_HI(net2226));
 sg13g2_tiehi _33687__2227 (.L_HI(net2227));
 sg13g2_tiehi _33686__2228 (.L_HI(net2228));
 sg13g2_tiehi _33685__2229 (.L_HI(net2229));
 sg13g2_tiehi _33684__2230 (.L_HI(net2230));
 sg13g2_tiehi _33683__2231 (.L_HI(net2231));
 sg13g2_tiehi _33682__2232 (.L_HI(net2232));
 sg13g2_tiehi _33681__2233 (.L_HI(net2233));
 sg13g2_tiehi _33680__2234 (.L_HI(net2234));
 sg13g2_tiehi _33679__2235 (.L_HI(net2235));
 sg13g2_tiehi _33678__2236 (.L_HI(net2236));
 sg13g2_tiehi _33677__2237 (.L_HI(net2237));
 sg13g2_tiehi _33676__2238 (.L_HI(net2238));
 sg13g2_tiehi _33675__2239 (.L_HI(net2239));
 sg13g2_tiehi _33674__2240 (.L_HI(net2240));
 sg13g2_tiehi _33673__2241 (.L_HI(net2241));
 sg13g2_tiehi _33672__2242 (.L_HI(net2242));
 sg13g2_tiehi _33671__2243 (.L_HI(net2243));
 sg13g2_tiehi _33670__2244 (.L_HI(net2244));
 sg13g2_tiehi _33669__2245 (.L_HI(net2245));
 sg13g2_tiehi _33668__2246 (.L_HI(net2246));
 sg13g2_tiehi _33667__2247 (.L_HI(net2247));
 sg13g2_tiehi _33666__2248 (.L_HI(net2248));
 sg13g2_tiehi _33665__2249 (.L_HI(net2249));
 sg13g2_tiehi _33664__2250 (.L_HI(net2250));
 sg13g2_tiehi _33663__2251 (.L_HI(net2251));
 sg13g2_tiehi _33662__2252 (.L_HI(net2252));
 sg13g2_tiehi _33661__2253 (.L_HI(net2253));
 sg13g2_tiehi _33660__2254 (.L_HI(net2254));
 sg13g2_tiehi _33659__2255 (.L_HI(net2255));
 sg13g2_tiehi _33658__2256 (.L_HI(net2256));
 sg13g2_tiehi _33657__2257 (.L_HI(net2257));
 sg13g2_tiehi _33656__2258 (.L_HI(net2258));
 sg13g2_tiehi _33655__2259 (.L_HI(net2259));
 sg13g2_tiehi _33654__2260 (.L_HI(net2260));
 sg13g2_tiehi _33653__2261 (.L_HI(net2261));
 sg13g2_tiehi _33652__2262 (.L_HI(net2262));
 sg13g2_tiehi _33651__2263 (.L_HI(net2263));
 sg13g2_tiehi _33650__2264 (.L_HI(net2264));
 sg13g2_tiehi _33649__2265 (.L_HI(net2265));
 sg13g2_tiehi _33648__2266 (.L_HI(net2266));
 sg13g2_tiehi _33647__2267 (.L_HI(net2267));
 sg13g2_tiehi _33646__2268 (.L_HI(net2268));
 sg13g2_tiehi _33645__2269 (.L_HI(net2269));
 sg13g2_tiehi _33644__2270 (.L_HI(net2270));
 sg13g2_tiehi _33643__2271 (.L_HI(net2271));
 sg13g2_tiehi _33642__2272 (.L_HI(net2272));
 sg13g2_tiehi _33641__2273 (.L_HI(net2273));
 sg13g2_tiehi _33640__2274 (.L_HI(net2274));
 sg13g2_tiehi _35390__2275 (.L_HI(net2275));
 sg13g2_tiehi _33639__2276 (.L_HI(net2276));
 sg13g2_tiehi _35992__2277 (.L_HI(net2277));
 sg13g2_tiehi _33638__2278 (.L_HI(net2278));
 sg13g2_tiehi _35389__2279 (.L_HI(net2279));
 sg13g2_tiehi _33637__2280 (.L_HI(net2280));
 sg13g2_tiehi _35991__2281 (.L_HI(net2281));
 sg13g2_tiehi _33636__2282 (.L_HI(net2282));
 sg13g2_tiehi _35388__2283 (.L_HI(net2283));
 sg13g2_tiehi _33635__2284 (.L_HI(net2284));
 sg13g2_tiehi _35990__2285 (.L_HI(net2285));
 sg13g2_tiehi _33634__2286 (.L_HI(net2286));
 sg13g2_tiehi _35387__2287 (.L_HI(net2287));
 sg13g2_tiehi _33633__2288 (.L_HI(net2288));
 sg13g2_tiehi _35989__2289 (.L_HI(net2289));
 sg13g2_tiehi _33632__2290 (.L_HI(net2290));
 sg13g2_tiehi _35386__2291 (.L_HI(net2291));
 sg13g2_tiehi _33631__2292 (.L_HI(net2292));
 sg13g2_tiehi _35988__2293 (.L_HI(net2293));
 sg13g2_tiehi _33630__2294 (.L_HI(net2294));
 sg13g2_tiehi _35385__2295 (.L_HI(net2295));
 sg13g2_tiehi _33629__2296 (.L_HI(net2296));
 sg13g2_tiehi _35987__2297 (.L_HI(net2297));
 sg13g2_tiehi _33628__2298 (.L_HI(net2298));
 sg13g2_tiehi _35384__2299 (.L_HI(net2299));
 sg13g2_tiehi _33627__2300 (.L_HI(net2300));
 sg13g2_tiehi _35986__2301 (.L_HI(net2301));
 sg13g2_tiehi _33626__2302 (.L_HI(net2302));
 sg13g2_tiehi _35383__2303 (.L_HI(net2303));
 sg13g2_tiehi _33625__2304 (.L_HI(net2304));
 sg13g2_tiehi _35985__2305 (.L_HI(net2305));
 sg13g2_tiehi _33624__2306 (.L_HI(net2306));
 sg13g2_tiehi _35382__2307 (.L_HI(net2307));
 sg13g2_tiehi _33623__2308 (.L_HI(net2308));
 sg13g2_tiehi _35984__2309 (.L_HI(net2309));
 sg13g2_tiehi _33622__2310 (.L_HI(net2310));
 sg13g2_tiehi _35381__2311 (.L_HI(net2311));
 sg13g2_tiehi _33621__2312 (.L_HI(net2312));
 sg13g2_tiehi _35983__2313 (.L_HI(net2313));
 sg13g2_tiehi _33620__2314 (.L_HI(net2314));
 sg13g2_tiehi _35380__2315 (.L_HI(net2315));
 sg13g2_tiehi _33619__2316 (.L_HI(net2316));
 sg13g2_tiehi _35982__2317 (.L_HI(net2317));
 sg13g2_tiehi _33618__2318 (.L_HI(net2318));
 sg13g2_tiehi _35379__2319 (.L_HI(net2319));
 sg13g2_tiehi _33617__2320 (.L_HI(net2320));
 sg13g2_tiehi _35378__2321 (.L_HI(net2321));
 sg13g2_tiehi _35377__2322 (.L_HI(net2322));
 sg13g2_tiehi _35376__2323 (.L_HI(net2323));
 sg13g2_tiehi _35375__2324 (.L_HI(net2324));
 sg13g2_tiehi _35374__2325 (.L_HI(net2325));
 sg13g2_tiehi _35373__2326 (.L_HI(net2326));
 sg13g2_tiehi _35372__2327 (.L_HI(net2327));
 sg13g2_tiehi _35371__2328 (.L_HI(net2328));
 sg13g2_tiehi _35370__2329 (.L_HI(net2329));
 sg13g2_tiehi _35369__2330 (.L_HI(net2330));
 sg13g2_tiehi _35368__2331 (.L_HI(net2331));
 sg13g2_tiehi _35367__2332 (.L_HI(net2332));
 sg13g2_tiehi _35007__2333 (.L_HI(net2333));
 sg13g2_tiehi _35934__2334 (.L_HI(net2334));
 sg13g2_tiehi _35935__2335 (.L_HI(net2335));
 sg13g2_tiehi _35936__2336 (.L_HI(net2336));
 sg13g2_tiehi _35937__2337 (.L_HI(net2337));
 sg13g2_tiehi _35938__2338 (.L_HI(net2338));
 sg13g2_tiehi _35939__2339 (.L_HI(net2339));
 sg13g2_tiehi _35366__2340 (.L_HI(net2340));
 sg13g2_tiehi _35365__2341 (.L_HI(net2341));
 sg13g2_tiehi _35364__2342 (.L_HI(net2342));
 sg13g2_tiehi _35363__2343 (.L_HI(net2343));
 sg13g2_tiehi _35362__2344 (.L_HI(net2344));
 sg13g2_tiehi _35361__2345 (.L_HI(net2345));
 sg13g2_tiehi _35360__2346 (.L_HI(net2346));
 sg13g2_tiehi _35359__2347 (.L_HI(net2347));
 sg13g2_tiehi _35358__2348 (.L_HI(net2348));
 sg13g2_tiehi _35357__2349 (.L_HI(net2349));
 sg13g2_tiehi _35356__2350 (.L_HI(net2350));
 sg13g2_tiehi _35355__2351 (.L_HI(net2351));
 sg13g2_tiehi _35354__2352 (.L_HI(net2352));
 sg13g2_tiehi _35353__2353 (.L_HI(net2353));
 sg13g2_tiehi _35352__2354 (.L_HI(net2354));
 sg13g2_tiehi _35351__2355 (.L_HI(net2355));
 sg13g2_tiehi _35350__2356 (.L_HI(net2356));
 sg13g2_tiehi _35349__2357 (.L_HI(net2357));
 sg13g2_tiehi _35348__2358 (.L_HI(net2358));
 sg13g2_tiehi _35347__2359 (.L_HI(net2359));
 sg13g2_tiehi _35346__2360 (.L_HI(net2360));
 sg13g2_tiehi _35345__2361 (.L_HI(net2361));
 sg13g2_tiehi _35344__2362 (.L_HI(net2362));
 sg13g2_tiehi _35343__2363 (.L_HI(net2363));
 sg13g2_tiehi _35342__2364 (.L_HI(net2364));
 sg13g2_tiehi _35341__2365 (.L_HI(net2365));
 sg13g2_tiehi _35340__2366 (.L_HI(net2366));
 sg13g2_tiehi _35339__2367 (.L_HI(net2367));
 sg13g2_tiehi _35338__2368 (.L_HI(net2368));
 sg13g2_tiehi _35337__2369 (.L_HI(net2369));
 sg13g2_tiehi _35336__2370 (.L_HI(net2370));
 sg13g2_tiehi _35335__2371 (.L_HI(net2371));
 sg13g2_tiehi _35334__2372 (.L_HI(net2372));
 sg13g2_tiehi _35333__2373 (.L_HI(net2373));
 sg13g2_tiehi _35332__2374 (.L_HI(net2374));
 sg13g2_tiehi _35331__2375 (.L_HI(net2375));
 sg13g2_tiehi _35330__2376 (.L_HI(net2376));
 sg13g2_tiehi _35329__2377 (.L_HI(net2377));
 sg13g2_tiehi _35328__2378 (.L_HI(net2378));
 sg13g2_tiehi _35327__2379 (.L_HI(net2379));
 sg13g2_tiehi _35326__2380 (.L_HI(net2380));
 sg13g2_tiehi _35325__2381 (.L_HI(net2381));
 sg13g2_tiehi _35324__2382 (.L_HI(net2382));
 sg13g2_tiehi _35323__2383 (.L_HI(net2383));
 sg13g2_tiehi _35322__2384 (.L_HI(net2384));
 sg13g2_tiehi _35321__2385 (.L_HI(net2385));
 sg13g2_tiehi _35320__2386 (.L_HI(net2386));
 sg13g2_tiehi _35319__2387 (.L_HI(net2387));
 sg13g2_tiehi _35318__2388 (.L_HI(net2388));
 sg13g2_tiehi _35317__2389 (.L_HI(net2389));
 sg13g2_tiehi _35316__2390 (.L_HI(net2390));
 sg13g2_tiehi _35315__2391 (.L_HI(net2391));
 sg13g2_tiehi _35314__2392 (.L_HI(net2392));
 sg13g2_tiehi _35313__2393 (.L_HI(net2393));
 sg13g2_tiehi _35312__2394 (.L_HI(net2394));
 sg13g2_tiehi _35311__2395 (.L_HI(net2395));
 sg13g2_tiehi _35310__2396 (.L_HI(net2396));
 sg13g2_tiehi _35309__2397 (.L_HI(net2397));
 sg13g2_tiehi _35308__2398 (.L_HI(net2398));
 sg13g2_tiehi _35307__2399 (.L_HI(net2399));
 sg13g2_tiehi _35306__2400 (.L_HI(net2400));
 sg13g2_tiehi _35305__2401 (.L_HI(net2401));
 sg13g2_tiehi _35304__2402 (.L_HI(net2402));
 sg13g2_tiehi _35303__2403 (.L_HI(net2403));
 sg13g2_tiehi _35302__2404 (.L_HI(net2404));
 sg13g2_tiehi _35301__2405 (.L_HI(net2405));
 sg13g2_tiehi _35300__2406 (.L_HI(net2406));
 sg13g2_tiehi _35299__2407 (.L_HI(net2407));
 sg13g2_tiehi _35298__2408 (.L_HI(net2408));
 sg13g2_tiehi _35297__2409 (.L_HI(net2409));
 sg13g2_tiehi _35296__2410 (.L_HI(net2410));
 sg13g2_tiehi _35295__2411 (.L_HI(net2411));
 sg13g2_tiehi _35294__2412 (.L_HI(net2412));
 sg13g2_tiehi _35293__2413 (.L_HI(net2413));
 sg13g2_tiehi _35292__2414 (.L_HI(net2414));
 sg13g2_tiehi _35981__2415 (.L_HI(net2415));
 sg13g2_tiehi _35291__2416 (.L_HI(net2416));
 sg13g2_tiehi _35980__2417 (.L_HI(net2417));
 sg13g2_tiehi _35290__2418 (.L_HI(net2418));
 sg13g2_tiehi _35979__2419 (.L_HI(net2419));
 sg13g2_tiehi _35289__2420 (.L_HI(net2420));
 sg13g2_tiehi _35978__2421 (.L_HI(net2421));
 sg13g2_tiehi _35288__2422 (.L_HI(net2422));
 sg13g2_tiehi _35977__2423 (.L_HI(net2423));
 sg13g2_tiehi _35287__2424 (.L_HI(net2424));
 sg13g2_tiehi _35976__2425 (.L_HI(net2425));
 sg13g2_tiehi _35286__2426 (.L_HI(net2426));
 sg13g2_tiehi _35975__2427 (.L_HI(net2427));
 sg13g2_tiehi _35285__2428 (.L_HI(net2428));
 sg13g2_tiehi _35974__2429 (.L_HI(net2429));
 sg13g2_tiehi _35284__2430 (.L_HI(net2430));
 sg13g2_tiehi _35973__2431 (.L_HI(net2431));
 sg13g2_tiehi _35283__2432 (.L_HI(net2432));
 sg13g2_tiehi _35972__2433 (.L_HI(net2433));
 sg13g2_tiehi _35282__2434 (.L_HI(net2434));
 sg13g2_tiehi _35971__2435 (.L_HI(net2435));
 sg13g2_tiehi _35281__2436 (.L_HI(net2436));
 sg13g2_tiehi _35280__2437 (.L_HI(net2437));
 sg13g2_tiehi _35970__2438 (.L_HI(net2438));
 sg13g2_tiehi _35279__2439 (.L_HI(net2439));
 sg13g2_tiehi _35969__2440 (.L_HI(net2440));
 sg13g2_tiehi _35278__2441 (.L_HI(net2441));
 sg13g2_tiehi _35277__2442 (.L_HI(net2442));
 sg13g2_tiehi _35276__2443 (.L_HI(net2443));
 sg13g2_tiehi _35275__2444 (.L_HI(net2444));
 sg13g2_tiehi _35968__2445 (.L_HI(net2445));
 sg13g2_tiehi _35274__2446 (.L_HI(net2446));
 sg13g2_tiehi _35940__2447 (.L_HI(net2447));
 sg13g2_tiehi _35273__2448 (.L_HI(net2448));
 sg13g2_tiehi _35967__2449 (.L_HI(net2449));
 sg13g2_tiehi _35272__2450 (.L_HI(net2450));
 sg13g2_tiehi _36195__2451 (.L_HI(net2451));
 sg13g2_tiehi _35271__2452 (.L_HI(net2452));
 sg13g2_tiehi _35966__2453 (.L_HI(net2453));
 sg13g2_tiehi _35270__2454 (.L_HI(net2454));
 sg13g2_tiehi _36194__2455 (.L_HI(net2455));
 sg13g2_tiehi _35269__2456 (.L_HI(net2456));
 sg13g2_tiehi _35965__2457 (.L_HI(net2457));
 sg13g2_tiehi _35268__2458 (.L_HI(net2458));
 sg13g2_tiehi _36193__2459 (.L_HI(net2459));
 sg13g2_tiehi _35267__2460 (.L_HI(net2460));
 sg13g2_tiehi _35964__2461 (.L_HI(net2461));
 sg13g2_tiehi _35266__2462 (.L_HI(net2462));
 sg13g2_tiehi _36192__2463 (.L_HI(net2463));
 sg13g2_tiehi _35265__2464 (.L_HI(net2464));
 sg13g2_tiehi _35963__2465 (.L_HI(net2465));
 sg13g2_tiehi _35264__2466 (.L_HI(net2466));
 sg13g2_tiehi _36191__2467 (.L_HI(net2467));
 sg13g2_tiehi _35263__2468 (.L_HI(net2468));
 sg13g2_tiehi _35962__2469 (.L_HI(net2469));
 sg13g2_tiehi _35262__2470 (.L_HI(net2470));
 sg13g2_tiehi _36190__2471 (.L_HI(net2471));
 sg13g2_tiehi _35261__2472 (.L_HI(net2472));
 sg13g2_tiehi _35961__2473 (.L_HI(net2473));
 sg13g2_tiehi _35260__2474 (.L_HI(net2474));
 sg13g2_tiehi _36189__2475 (.L_HI(net2475));
 sg13g2_tiehi _35259__2476 (.L_HI(net2476));
 sg13g2_tiehi _35960__2477 (.L_HI(net2477));
 sg13g2_tiehi _35258__2478 (.L_HI(net2478));
 sg13g2_tiehi _36188__2479 (.L_HI(net2479));
 sg13g2_tiehi _35257__2480 (.L_HI(net2480));
 sg13g2_tiehi _35959__2481 (.L_HI(net2481));
 sg13g2_tiehi _35256__2482 (.L_HI(net2482));
 sg13g2_tiehi _36187__2483 (.L_HI(net2483));
 sg13g2_tiehi _35255__2484 (.L_HI(net2484));
 sg13g2_tiehi _35958__2485 (.L_HI(net2485));
 sg13g2_tiehi _35254__2486 (.L_HI(net2486));
 sg13g2_tiehi _36186__2487 (.L_HI(net2487));
 sg13g2_tiehi _35253__2488 (.L_HI(net2488));
 sg13g2_tiehi _35957__2489 (.L_HI(net2489));
 sg13g2_tiehi _35252__2490 (.L_HI(net2490));
 sg13g2_tiehi _36185__2491 (.L_HI(net2491));
 sg13g2_tiehi _35251__2492 (.L_HI(net2492));
 sg13g2_tiehi _35956__2493 (.L_HI(net2493));
 sg13g2_tiehi _35250__2494 (.L_HI(net2494));
 sg13g2_tiehi _36184__2495 (.L_HI(net2495));
 sg13g2_tiehi _35249__2496 (.L_HI(net2496));
 sg13g2_tiehi _35955__2497 (.L_HI(net2497));
 sg13g2_tiehi _35248__2498 (.L_HI(net2498));
 sg13g2_tiehi _36183__2499 (.L_HI(net2499));
 sg13g2_tiehi _35247__2500 (.L_HI(net2500));
 sg13g2_tiehi _35954__2501 (.L_HI(net2501));
 sg13g2_tiehi _35246__2502 (.L_HI(net2502));
 sg13g2_tiehi _36182__2503 (.L_HI(net2503));
 sg13g2_tiehi _35245__2504 (.L_HI(net2504));
 sg13g2_tiehi _35953__2505 (.L_HI(net2505));
 sg13g2_tiehi _35244__2506 (.L_HI(net2506));
 sg13g2_tiehi _36181__2507 (.L_HI(net2507));
 sg13g2_tiehi _35243__2508 (.L_HI(net2508));
 sg13g2_tiehi _35952__2509 (.L_HI(net2509));
 sg13g2_tiehi _35242__2510 (.L_HI(net2510));
 sg13g2_tiehi _36180__2511 (.L_HI(net2511));
 sg13g2_tiehi _35241__2512 (.L_HI(net2512));
 sg13g2_tiehi _35951__2513 (.L_HI(net2513));
 sg13g2_tiehi _35240__2514 (.L_HI(net2514));
 sg13g2_tiehi _36179__2515 (.L_HI(net2515));
 sg13g2_tiehi _35239__2516 (.L_HI(net2516));
 sg13g2_tiehi _35950__2517 (.L_HI(net2517));
 sg13g2_tiehi _35238__2518 (.L_HI(net2518));
 sg13g2_tiehi _36178__2519 (.L_HI(net2519));
 sg13g2_tiehi _35237__2520 (.L_HI(net2520));
 sg13g2_tiehi _35949__2521 (.L_HI(net2521));
 sg13g2_tiehi _35236__2522 (.L_HI(net2522));
 sg13g2_tiehi _35235__2523 (.L_HI(net2523));
 sg13g2_tiehi _35234__2524 (.L_HI(net2524));
 sg13g2_tiehi _35233__2525 (.L_HI(net2525));
 sg13g2_tiehi _35232__2526 (.L_HI(net2526));
 sg13g2_tiehi _35231__2527 (.L_HI(net2527));
 sg13g2_tiehi _35230__2528 (.L_HI(net2528));
 sg13g2_tiehi _35229__2529 (.L_HI(net2529));
 sg13g2_tiehi _35228__2530 (.L_HI(net2530));
 sg13g2_tiehi _35227__2531 (.L_HI(net2531));
 sg13g2_tiehi _35226__2532 (.L_HI(net2532));
 sg13g2_tiehi _35225__2533 (.L_HI(net2533));
 sg13g2_tiehi _35224__2534 (.L_HI(net2534));
 sg13g2_tiehi _35223__2535 (.L_HI(net2535));
 sg13g2_tiehi _35222__2536 (.L_HI(net2536));
 sg13g2_tiehi _35221__2537 (.L_HI(net2537));
 sg13g2_tiehi _35220__2538 (.L_HI(net2538));
 sg13g2_tiehi _35219__2539 (.L_HI(net2539));
 sg13g2_tiehi _35218__2540 (.L_HI(net2540));
 sg13g2_tiehi _35217__2541 (.L_HI(net2541));
 sg13g2_tiehi _35216__2542 (.L_HI(net2542));
 sg13g2_tiehi _35215__2543 (.L_HI(net2543));
 sg13g2_tiehi _35214__2544 (.L_HI(net2544));
 sg13g2_tiehi _35213__2545 (.L_HI(net2545));
 sg13g2_tiehi _35212__2546 (.L_HI(net2546));
 sg13g2_tiehi _35211__2547 (.L_HI(net2547));
 sg13g2_tiehi _35210__2548 (.L_HI(net2548));
 sg13g2_tiehi _35209__2549 (.L_HI(net2549));
 sg13g2_tiehi _35208__2550 (.L_HI(net2550));
 sg13g2_tiehi _35207__2551 (.L_HI(net2551));
 sg13g2_tiehi _35206__2552 (.L_HI(net2552));
 sg13g2_tiehi _35205__2553 (.L_HI(net2553));
 sg13g2_tiehi _35204__2554 (.L_HI(net2554));
 sg13g2_tiehi _36177__2555 (.L_HI(net2555));
 sg13g2_tiehi _35203__2556 (.L_HI(net2556));
 sg13g2_tiehi _35948__2557 (.L_HI(net2557));
 sg13g2_tiehi _35202__2558 (.L_HI(net2558));
 sg13g2_tiehi _36176__2559 (.L_HI(net2559));
 sg13g2_tiehi _35201__2560 (.L_HI(net2560));
 sg13g2_tiehi _35947__2561 (.L_HI(net2561));
 sg13g2_tiehi _35200__2562 (.L_HI(net2562));
 sg13g2_tiehi _36175__2563 (.L_HI(net2563));
 sg13g2_tiehi _35199__2564 (.L_HI(net2564));
 sg13g2_tiehi _35946__2565 (.L_HI(net2565));
 sg13g2_tiehi _35198__2566 (.L_HI(net2566));
 sg13g2_tiehi _36174__2567 (.L_HI(net2567));
 sg13g2_tiehi _35197__2568 (.L_HI(net2568));
 sg13g2_tiehi _35945__2569 (.L_HI(net2569));
 sg13g2_tiehi _35196__2570 (.L_HI(net2570));
 sg13g2_tiehi _36173__2571 (.L_HI(net2571));
 sg13g2_tiehi _35195__2572 (.L_HI(net2572));
 sg13g2_tiehi _35194__2573 (.L_HI(net2573));
 sg13g2_tiehi _35193__2574 (.L_HI(net2574));
 sg13g2_tiehi _35192__2575 (.L_HI(net2575));
 sg13g2_tiehi _35191__2576 (.L_HI(net2576));
 sg13g2_tiehi _35190__2577 (.L_HI(net2577));
 sg13g2_tiehi _35944__2578 (.L_HI(net2578));
 sg13g2_tiehi _35189__2579 (.L_HI(net2579));
 sg13g2_tiehi _36172__2580 (.L_HI(net2580));
 sg13g2_tiehi _35188__2581 (.L_HI(net2581));
 sg13g2_tiehi _35943__2582 (.L_HI(net2582));
 sg13g2_tiehi _35187__2583 (.L_HI(net2583));
 sg13g2_tiehi _36171__2584 (.L_HI(net2584));
 sg13g2_tiehi _35186__2585 (.L_HI(net2585));
 sg13g2_tiehi _35942__2586 (.L_HI(net2586));
 sg13g2_tiehi _35185__2587 (.L_HI(net2587));
 sg13g2_tiehi _35941__2588 (.L_HI(net2588));
 sg13g2_tiehi _35184__2589 (.L_HI(net2589));
 sg13g2_tiehi _35933__2590 (.L_HI(net2590));
 sg13g2_tiehi _35183__2591 (.L_HI(net2591));
 sg13g2_tiehi _35932__2592 (.L_HI(net2592));
 sg13g2_tiehi _35182__2593 (.L_HI(net2593));
 sg13g2_tiehi tt_um_kianV_rv32ima_uLinux_SoC_2594 (.L_HI(net2594));
 sg13g2_tiehi tt_um_kianV_rv32ima_uLinux_SoC_2595 (.L_HI(net2595));
 sg13g2_tiehi tt_um_kianV_rv32ima_uLinux_SoC_2596 (.L_HI(net2596));
 sg13g2_tiehi tt_um_kianV_rv32ima_uLinux_SoC_2597 (.L_HI(net2597));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_4 _38780_ (.X(uio_oe[2]),
    .A(uio_oe[5]));
 sg13g2_buf_4 _38781_ (.X(uio_oe[4]),
    .A(uio_oe[5]));
 sg13g2_buf_4 _38782_ (.X(uio_out[1]),
    .A(sio0_si_mosi_o));
 sg13g2_buf_4 _38783_ (.X(uio_out[2]),
    .A(sio1_so_miso_o));
 sg13g2_buf_4 _38784_ (.X(uio_out[3]),
    .A(sclk));
 sg13g2_buf_4 _38785_ (.X(uio_out[4]),
    .A(sio2_o));
 sg13g2_buf_4 _38786_ (.X(uio_out[5]),
    .A(sio3_o));
 sg13g2_buf_4 fanout7326 (.X(net7326),
    .A(_05313_));
 sg13g2_buf_4 fanout7327 (.X(net7327),
    .A(net7328));
 sg13g2_buf_4 fanout7328 (.X(net7328),
    .A(net7329));
 sg13g2_buf_4 fanout7329 (.X(net7329),
    .A(_05312_));
 sg13g2_buf_4 fanout7330 (.X(net7330),
    .A(_05022_));
 sg13g2_buf_4 fanout7331 (.X(net7331),
    .A(net7332));
 sg13g2_buf_4 fanout7332 (.X(net7332),
    .A(net7333));
 sg13g2_buf_4 fanout7333 (.X(net7333),
    .A(_05021_));
 sg13g2_buf_4 fanout7334 (.X(net7334),
    .A(net7335));
 sg13g2_buf_2 fanout7335 (.A(_13829_),
    .X(net7335));
 sg13g2_buf_2 fanout7336 (.A(_13809_),
    .X(net7336));
 sg13g2_buf_2 fanout7337 (.A(net7338),
    .X(net7337));
 sg13g2_buf_2 fanout7338 (.A(net7341),
    .X(net7338));
 sg13g2_buf_2 fanout7339 (.A(net7340),
    .X(net7339));
 sg13g2_buf_2 fanout7340 (.A(net7341),
    .X(net7340));
 sg13g2_buf_4 fanout7341 (.X(net7341),
    .A(_05965_));
 sg13g2_buf_4 fanout7342 (.X(net7342),
    .A(net7347));
 sg13g2_buf_1 fanout7343 (.A(net7347),
    .X(net7343));
 sg13g2_buf_4 fanout7344 (.X(net7344),
    .A(net7347));
 sg13g2_buf_1 fanout7345 (.A(net7347),
    .X(net7345));
 sg13g2_buf_2 fanout7346 (.A(net7347),
    .X(net7346));
 sg13g2_buf_4 fanout7347 (.X(net7347),
    .A(_05965_));
 sg13g2_buf_4 fanout7348 (.X(net7348),
    .A(net7350));
 sg13g2_buf_2 fanout7349 (.A(net7350),
    .X(net7349));
 sg13g2_buf_4 fanout7350 (.X(net7350),
    .A(_05853_));
 sg13g2_buf_2 fanout7351 (.A(net7353),
    .X(net7351));
 sg13g2_buf_1 fanout7352 (.A(net7353),
    .X(net7352));
 sg13g2_buf_1 fanout7353 (.A(net7354),
    .X(net7353));
 sg13g2_buf_4 fanout7354 (.X(net7354),
    .A(net7360));
 sg13g2_buf_4 fanout7355 (.X(net7355),
    .A(net7357));
 sg13g2_buf_2 fanout7356 (.A(net7357),
    .X(net7356));
 sg13g2_buf_1 fanout7357 (.A(net7359),
    .X(net7357));
 sg13g2_buf_4 fanout7358 (.X(net7358),
    .A(net7359));
 sg13g2_buf_2 fanout7359 (.A(net7360),
    .X(net7359));
 sg13g2_buf_4 fanout7360 (.X(net7360),
    .A(_05853_));
 sg13g2_buf_4 fanout7361 (.X(net7361),
    .A(_13328_));
 sg13g2_buf_2 fanout7362 (.A(_13328_),
    .X(net7362));
 sg13g2_buf_2 fanout7363 (.A(_06665_),
    .X(net7363));
 sg13g2_buf_1 fanout7364 (.A(_06665_),
    .X(net7364));
 sg13g2_buf_4 fanout7365 (.X(net7365),
    .A(net7366));
 sg13g2_buf_4 fanout7366 (.X(net7366),
    .A(net7375));
 sg13g2_buf_4 fanout7367 (.X(net7367),
    .A(net7369));
 sg13g2_buf_4 fanout7368 (.X(net7368),
    .A(net7369));
 sg13g2_buf_2 fanout7369 (.A(net7370),
    .X(net7369));
 sg13g2_buf_4 fanout7370 (.X(net7370),
    .A(net7375));
 sg13g2_buf_2 fanout7371 (.A(net7374),
    .X(net7371));
 sg13g2_buf_2 fanout7372 (.A(net7373),
    .X(net7372));
 sg13g2_buf_2 fanout7373 (.A(net7374),
    .X(net7373));
 sg13g2_buf_4 fanout7374 (.X(net7374),
    .A(net7375));
 sg13g2_buf_2 fanout7375 (.A(_05854_),
    .X(net7375));
 sg13g2_buf_2 fanout7376 (.A(net7378),
    .X(net7376));
 sg13g2_buf_2 fanout7377 (.A(net7378),
    .X(net7377));
 sg13g2_buf_1 fanout7378 (.A(net7379),
    .X(net7378));
 sg13g2_buf_1 fanout7379 (.A(net7380),
    .X(net7379));
 sg13g2_buf_2 fanout7380 (.A(net7388),
    .X(net7380));
 sg13g2_buf_2 fanout7381 (.A(net7383),
    .X(net7381));
 sg13g2_buf_1 fanout7382 (.A(net7383),
    .X(net7382));
 sg13g2_buf_2 fanout7383 (.A(net7387),
    .X(net7383));
 sg13g2_buf_2 fanout7384 (.A(net7385),
    .X(net7384));
 sg13g2_buf_2 fanout7385 (.A(net7386),
    .X(net7385));
 sg13g2_buf_2 fanout7386 (.A(net7387),
    .X(net7386));
 sg13g2_buf_2 fanout7387 (.A(net7388),
    .X(net7387));
 sg13g2_buf_4 fanout7388 (.X(net7388),
    .A(_05031_));
 sg13g2_buf_2 fanout7389 (.A(_14277_),
    .X(net7389));
 sg13g2_buf_2 fanout7390 (.A(net7392),
    .X(net7390));
 sg13g2_buf_2 fanout7391 (.A(net7392),
    .X(net7391));
 sg13g2_buf_2 fanout7392 (.A(_07037_),
    .X(net7392));
 sg13g2_buf_2 fanout7393 (.A(_07037_),
    .X(net7393));
 sg13g2_buf_1 fanout7394 (.A(_07037_),
    .X(net7394));
 sg13g2_buf_4 fanout7395 (.X(net7395),
    .A(_07358_));
 sg13g2_buf_2 fanout7396 (.A(_06984_),
    .X(net7396));
 sg13g2_buf_4 fanout7397 (.X(net7397),
    .A(_14461_));
 sg13g2_buf_2 fanout7398 (.A(_14461_),
    .X(net7398));
 sg13g2_buf_2 fanout7399 (.A(net7404),
    .X(net7399));
 sg13g2_buf_2 fanout7400 (.A(net7401),
    .X(net7400));
 sg13g2_buf_2 fanout7401 (.A(net7404),
    .X(net7401));
 sg13g2_buf_2 fanout7402 (.A(net7404),
    .X(net7402));
 sg13g2_buf_1 fanout7403 (.A(net7404),
    .X(net7403));
 sg13g2_buf_2 fanout7404 (.A(_14034_),
    .X(net7404));
 sg13g2_buf_2 fanout7405 (.A(_13981_),
    .X(net7405));
 sg13g2_buf_2 fanout7406 (.A(_13981_),
    .X(net7406));
 sg13g2_buf_2 fanout7407 (.A(net7411),
    .X(net7407));
 sg13g2_buf_2 fanout7408 (.A(net7409),
    .X(net7408));
 sg13g2_buf_2 fanout7409 (.A(net7410),
    .X(net7409));
 sg13g2_buf_2 fanout7410 (.A(net7411),
    .X(net7410));
 sg13g2_buf_1 fanout7411 (.A(net7417),
    .X(net7411));
 sg13g2_buf_2 fanout7412 (.A(net7413),
    .X(net7412));
 sg13g2_buf_2 fanout7413 (.A(net7414),
    .X(net7413));
 sg13g2_buf_2 fanout7414 (.A(net7417),
    .X(net7414));
 sg13g2_buf_2 fanout7415 (.A(net7416),
    .X(net7415));
 sg13g2_buf_2 fanout7416 (.A(net7417),
    .X(net7416));
 sg13g2_buf_2 fanout7417 (.A(_07396_),
    .X(net7417));
 sg13g2_buf_4 fanout7418 (.X(net7418),
    .A(_07360_));
 sg13g2_buf_2 fanout7419 (.A(_06454_),
    .X(net7419));
 sg13g2_buf_2 fanout7420 (.A(_06444_),
    .X(net7420));
 sg13g2_buf_2 fanout7421 (.A(net7423),
    .X(net7421));
 sg13g2_buf_2 fanout7422 (.A(net7423),
    .X(net7422));
 sg13g2_buf_2 fanout7423 (.A(_14460_),
    .X(net7423));
 sg13g2_buf_4 fanout7424 (.X(net7424),
    .A(_13188_));
 sg13g2_buf_2 fanout7425 (.A(_13188_),
    .X(net7425));
 sg13g2_buf_2 fanout7426 (.A(net7427),
    .X(net7426));
 sg13g2_buf_2 fanout7427 (.A(net7428),
    .X(net7427));
 sg13g2_buf_1 fanout7428 (.A(net7429),
    .X(net7428));
 sg13g2_buf_2 fanout7429 (.A(net7430),
    .X(net7429));
 sg13g2_buf_2 fanout7430 (.A(_07359_),
    .X(net7430));
 sg13g2_buf_2 fanout7431 (.A(net7433),
    .X(net7431));
 sg13g2_buf_2 fanout7432 (.A(net7433),
    .X(net7432));
 sg13g2_buf_2 fanout7433 (.A(_07359_),
    .X(net7433));
 sg13g2_buf_2 fanout7434 (.A(_06257_),
    .X(net7434));
 sg13g2_buf_2 fanout7435 (.A(_14440_),
    .X(net7435));
 sg13g2_buf_1 fanout7436 (.A(_14440_),
    .X(net7436));
 sg13g2_buf_4 fanout7437 (.X(net7437),
    .A(net7439));
 sg13g2_buf_4 fanout7438 (.X(net7438),
    .A(net7439));
 sg13g2_buf_4 fanout7439 (.X(net7439),
    .A(_13230_));
 sg13g2_buf_2 fanout7440 (.A(net7441),
    .X(net7440));
 sg13g2_buf_4 fanout7441 (.X(net7441),
    .A(_13228_));
 sg13g2_buf_2 fanout7442 (.A(net7444),
    .X(net7442));
 sg13g2_buf_2 fanout7443 (.A(net7444),
    .X(net7443));
 sg13g2_buf_2 fanout7444 (.A(_13228_),
    .X(net7444));
 sg13g2_buf_2 fanout7445 (.A(net7446),
    .X(net7445));
 sg13g2_buf_4 fanout7446 (.X(net7446),
    .A(net7449));
 sg13g2_buf_4 fanout7447 (.X(net7447),
    .A(net7448));
 sg13g2_buf_4 fanout7448 (.X(net7448),
    .A(net7449));
 sg13g2_buf_2 fanout7449 (.A(_13215_),
    .X(net7449));
 sg13g2_buf_4 fanout7450 (.X(net7450),
    .A(net7451));
 sg13g2_buf_4 fanout7451 (.X(net7451),
    .A(_13214_));
 sg13g2_buf_4 fanout7452 (.X(net7452),
    .A(_13214_));
 sg13g2_buf_2 fanout7453 (.A(_13214_),
    .X(net7453));
 sg13g2_buf_2 fanout7454 (.A(_12555_),
    .X(net7454));
 sg13g2_buf_2 fanout7455 (.A(_12555_),
    .X(net7455));
 sg13g2_buf_2 fanout7456 (.A(net7457),
    .X(net7456));
 sg13g2_buf_2 fanout7457 (.A(net7458),
    .X(net7457));
 sg13g2_buf_2 fanout7458 (.A(_12555_),
    .X(net7458));
 sg13g2_buf_2 fanout7459 (.A(net7460),
    .X(net7459));
 sg13g2_buf_1 fanout7460 (.A(net7461),
    .X(net7460));
 sg13g2_buf_2 fanout7461 (.A(_12554_),
    .X(net7461));
 sg13g2_buf_2 fanout7462 (.A(net7463),
    .X(net7462));
 sg13g2_buf_2 fanout7463 (.A(net7464),
    .X(net7463));
 sg13g2_buf_2 fanout7464 (.A(_12554_),
    .X(net7464));
 sg13g2_buf_4 fanout7465 (.X(net7465),
    .A(net7466));
 sg13g2_buf_4 fanout7466 (.X(net7466),
    .A(_13213_));
 sg13g2_buf_4 fanout7467 (.X(net7467),
    .A(_13050_));
 sg13g2_buf_2 fanout7468 (.A(_13047_),
    .X(net7468));
 sg13g2_buf_2 fanout7469 (.A(_09005_),
    .X(net7469));
 sg13g2_buf_2 fanout7470 (.A(_12883_),
    .X(net7470));
 sg13g2_buf_2 fanout7471 (.A(net7472),
    .X(net7471));
 sg13g2_buf_4 fanout7472 (.X(net7472),
    .A(net7478));
 sg13g2_buf_2 fanout7473 (.A(net7474),
    .X(net7473));
 sg13g2_buf_2 fanout7474 (.A(net7477),
    .X(net7474));
 sg13g2_buf_2 fanout7475 (.A(net7477),
    .X(net7475));
 sg13g2_buf_1 fanout7476 (.A(net7477),
    .X(net7476));
 sg13g2_buf_4 fanout7477 (.X(net7477),
    .A(net7478));
 sg13g2_buf_4 fanout7478 (.X(net7478),
    .A(net7479));
 sg13g2_buf_4 fanout7479 (.X(net7479),
    .A(_12468_));
 sg13g2_buf_4 fanout7480 (.X(net7480),
    .A(_12467_));
 sg13g2_buf_4 fanout7481 (.X(net7481),
    .A(net7483));
 sg13g2_buf_2 fanout7482 (.A(net7483),
    .X(net7482));
 sg13g2_buf_4 fanout7483 (.X(net7483),
    .A(net7484));
 sg13g2_buf_2 fanout7484 (.A(_12467_),
    .X(net7484));
 sg13g2_buf_4 fanout7485 (.X(net7485),
    .A(net7487));
 sg13g2_buf_4 fanout7486 (.X(net7486),
    .A(net7487));
 sg13g2_buf_2 fanout7487 (.A(net7490),
    .X(net7487));
 sg13g2_buf_2 fanout7488 (.A(net7490),
    .X(net7488));
 sg13g2_buf_1 fanout7489 (.A(net7490),
    .X(net7489));
 sg13g2_buf_8 fanout7490 (.A(_11756_),
    .X(net7490));
 sg13g2_buf_4 fanout7491 (.X(net7491),
    .A(net7493));
 sg13g2_buf_2 fanout7492 (.A(net7493),
    .X(net7492));
 sg13g2_buf_4 fanout7493 (.X(net7493),
    .A(_12894_));
 sg13g2_buf_2 fanout7494 (.A(net7498),
    .X(net7494));
 sg13g2_buf_2 fanout7495 (.A(net7497),
    .X(net7495));
 sg13g2_buf_2 fanout7496 (.A(net7498),
    .X(net7496));
 sg13g2_buf_4 fanout7497 (.X(net7497),
    .A(net7498));
 sg13g2_buf_8 fanout7498 (.A(_13145_),
    .X(net7498));
 sg13g2_buf_4 fanout7499 (.X(net7499),
    .A(net7500));
 sg13g2_buf_4 fanout7500 (.X(net7500),
    .A(net7501));
 sg13g2_buf_4 fanout7501 (.X(net7501),
    .A(net7503));
 sg13g2_buf_2 fanout7502 (.A(net7503),
    .X(net7502));
 sg13g2_buf_8 fanout7503 (.A(_13132_),
    .X(net7503));
 sg13g2_buf_2 fanout7504 (.A(net7509),
    .X(net7504));
 sg13g2_buf_1 fanout7505 (.A(net7509),
    .X(net7505));
 sg13g2_buf_4 fanout7506 (.X(net7506),
    .A(net7508));
 sg13g2_buf_2 fanout7507 (.A(net7508),
    .X(net7507));
 sg13g2_buf_2 fanout7508 (.A(net7509),
    .X(net7508));
 sg13g2_buf_4 fanout7509 (.X(net7509),
    .A(net7510));
 sg13g2_buf_8 fanout7510 (.A(_13119_),
    .X(net7510));
 sg13g2_buf_2 fanout7511 (.A(net7512),
    .X(net7511));
 sg13g2_buf_4 fanout7512 (.X(net7512),
    .A(net7515));
 sg13g2_buf_2 fanout7513 (.A(net7514),
    .X(net7513));
 sg13g2_buf_4 fanout7514 (.X(net7514),
    .A(net7515));
 sg13g2_buf_8 fanout7515 (.A(_13108_),
    .X(net7515));
 sg13g2_buf_4 fanout7516 (.X(net7516),
    .A(net7517));
 sg13g2_buf_1 fanout7517 (.A(net7521),
    .X(net7517));
 sg13g2_buf_4 fanout7518 (.X(net7518),
    .A(net7519));
 sg13g2_buf_2 fanout7519 (.A(net7520),
    .X(net7519));
 sg13g2_buf_2 fanout7520 (.A(net7521),
    .X(net7520));
 sg13g2_buf_4 fanout7521 (.X(net7521),
    .A(_13095_));
 sg13g2_buf_2 fanout7522 (.A(net7523),
    .X(net7522));
 sg13g2_buf_2 fanout7523 (.A(net7525),
    .X(net7523));
 sg13g2_buf_4 fanout7524 (.X(net7524),
    .A(net7525));
 sg13g2_buf_4 fanout7525 (.X(net7525),
    .A(net7527));
 sg13g2_buf_4 fanout7526 (.X(net7526),
    .A(net7527));
 sg13g2_buf_4 fanout7527 (.X(net7527),
    .A(_13084_));
 sg13g2_buf_2 fanout7528 (.A(net7529),
    .X(net7528));
 sg13g2_buf_2 fanout7529 (.A(net7533),
    .X(net7529));
 sg13g2_buf_4 fanout7530 (.X(net7530),
    .A(net7532));
 sg13g2_buf_2 fanout7531 (.A(net7532),
    .X(net7531));
 sg13g2_buf_2 fanout7532 (.A(net7533),
    .X(net7532));
 sg13g2_buf_8 fanout7533 (.A(_13073_),
    .X(net7533));
 sg13g2_buf_4 fanout7534 (.X(net7534),
    .A(net7535));
 sg13g2_buf_1 fanout7535 (.A(net7536),
    .X(net7535));
 sg13g2_buf_4 fanout7536 (.X(net7536),
    .A(net7539));
 sg13g2_buf_4 fanout7537 (.X(net7537),
    .A(net7538));
 sg13g2_buf_2 fanout7538 (.A(net7539),
    .X(net7538));
 sg13g2_buf_8 fanout7539 (.A(_13062_),
    .X(net7539));
 sg13g2_buf_2 fanout7540 (.A(net7542),
    .X(net7540));
 sg13g2_buf_2 fanout7541 (.A(net7542),
    .X(net7541));
 sg13g2_buf_2 fanout7542 (.A(net7545),
    .X(net7542));
 sg13g2_buf_2 fanout7543 (.A(net7544),
    .X(net7543));
 sg13g2_buf_4 fanout7544 (.X(net7544),
    .A(net7545));
 sg13g2_buf_8 fanout7545 (.A(_13039_),
    .X(net7545));
 sg13g2_buf_2 fanout7546 (.A(net7547),
    .X(net7546));
 sg13g2_buf_2 fanout7547 (.A(net7550),
    .X(net7547));
 sg13g2_buf_2 fanout7548 (.A(net7549),
    .X(net7548));
 sg13g2_buf_2 fanout7549 (.A(net7550),
    .X(net7549));
 sg13g2_buf_8 fanout7550 (.A(_13029_),
    .X(net7550));
 sg13g2_buf_2 fanout7551 (.A(net7556),
    .X(net7551));
 sg13g2_buf_2 fanout7552 (.A(net7555),
    .X(net7552));
 sg13g2_buf_1 fanout7553 (.A(net7554),
    .X(net7553));
 sg13g2_buf_2 fanout7554 (.A(net7555),
    .X(net7554));
 sg13g2_buf_2 fanout7555 (.A(net7556),
    .X(net7555));
 sg13g2_buf_8 fanout7556 (.A(_13018_),
    .X(net7556));
 sg13g2_buf_4 fanout7557 (.X(net7557),
    .A(net7559));
 sg13g2_buf_2 fanout7558 (.A(net7559),
    .X(net7558));
 sg13g2_buf_1 fanout7559 (.A(net7562),
    .X(net7559));
 sg13g2_buf_2 fanout7560 (.A(net7561),
    .X(net7560));
 sg13g2_buf_2 fanout7561 (.A(net7562),
    .X(net7561));
 sg13g2_buf_4 fanout7562 (.X(net7562),
    .A(_13007_));
 sg13g2_buf_2 fanout7563 (.A(net7564),
    .X(net7563));
 sg13g2_buf_4 fanout7564 (.X(net7564),
    .A(net7565));
 sg13g2_buf_4 fanout7565 (.X(net7565),
    .A(net7567));
 sg13g2_buf_4 fanout7566 (.X(net7566),
    .A(net7567));
 sg13g2_buf_4 fanout7567 (.X(net7567),
    .A(_12997_));
 sg13g2_buf_4 fanout7568 (.X(net7568),
    .A(net7572));
 sg13g2_buf_2 fanout7569 (.A(net7572),
    .X(net7569));
 sg13g2_buf_4 fanout7570 (.X(net7570),
    .A(net7572));
 sg13g2_buf_2 fanout7571 (.A(net7572),
    .X(net7571));
 sg13g2_buf_2 fanout7572 (.A(net7573),
    .X(net7572));
 sg13g2_buf_8 fanout7573 (.A(_12986_),
    .X(net7573));
 sg13g2_buf_2 fanout7574 (.A(net7577),
    .X(net7574));
 sg13g2_buf_2 fanout7575 (.A(net7577),
    .X(net7575));
 sg13g2_buf_4 fanout7576 (.X(net7576),
    .A(net7577));
 sg13g2_buf_2 fanout7577 (.A(net7579),
    .X(net7577));
 sg13g2_buf_2 fanout7578 (.A(net7579),
    .X(net7578));
 sg13g2_buf_8 fanout7579 (.A(_12975_),
    .X(net7579));
 sg13g2_buf_2 fanout7580 (.A(net7581),
    .X(net7580));
 sg13g2_buf_2 fanout7581 (.A(net7582),
    .X(net7581));
 sg13g2_buf_4 fanout7582 (.X(net7582),
    .A(_12964_));
 sg13g2_buf_2 fanout7583 (.A(net7584),
    .X(net7583));
 sg13g2_buf_1 fanout7584 (.A(net7585),
    .X(net7584));
 sg13g2_buf_4 fanout7585 (.X(net7585),
    .A(_12964_));
 sg13g2_buf_4 fanout7586 (.X(net7586),
    .A(net7591));
 sg13g2_buf_1 fanout7587 (.A(net7591),
    .X(net7587));
 sg13g2_buf_2 fanout7588 (.A(net7590),
    .X(net7588));
 sg13g2_buf_2 fanout7589 (.A(net7590),
    .X(net7589));
 sg13g2_buf_2 fanout7590 (.A(net7591),
    .X(net7590));
 sg13g2_buf_8 fanout7591 (.A(_12951_),
    .X(net7591));
 sg13g2_buf_2 fanout7592 (.A(net7596),
    .X(net7592));
 sg13g2_buf_2 fanout7593 (.A(net7596),
    .X(net7593));
 sg13g2_buf_2 fanout7594 (.A(net7595),
    .X(net7594));
 sg13g2_buf_2 fanout7595 (.A(net7596),
    .X(net7595));
 sg13g2_buf_8 fanout7596 (.A(_12939_),
    .X(net7596));
 sg13g2_buf_2 fanout7597 (.A(net7598),
    .X(net7597));
 sg13g2_buf_4 fanout7598 (.X(net7598),
    .A(net7601));
 sg13g2_buf_2 fanout7599 (.A(net7600),
    .X(net7599));
 sg13g2_buf_2 fanout7600 (.A(net7601),
    .X(net7600));
 sg13g2_buf_2 fanout7601 (.A(_12928_),
    .X(net7601));
 sg13g2_buf_4 fanout7602 (.X(net7602),
    .A(net7603));
 sg13g2_buf_4 fanout7603 (.X(net7603),
    .A(_12918_));
 sg13g2_buf_2 fanout7604 (.A(net7605),
    .X(net7604));
 sg13g2_buf_2 fanout7605 (.A(net7606),
    .X(net7605));
 sg13g2_buf_8 fanout7606 (.A(_12918_),
    .X(net7606));
 sg13g2_buf_2 fanout7607 (.A(net7608),
    .X(net7607));
 sg13g2_buf_4 fanout7608 (.X(net7608),
    .A(net7611));
 sg13g2_buf_4 fanout7609 (.X(net7609),
    .A(net7610));
 sg13g2_buf_2 fanout7610 (.A(net7611),
    .X(net7610));
 sg13g2_buf_4 fanout7611 (.X(net7611),
    .A(_12905_));
 sg13g2_buf_4 fanout7612 (.X(net7612),
    .A(net7616));
 sg13g2_buf_2 fanout7613 (.A(net7616),
    .X(net7613));
 sg13g2_buf_4 fanout7614 (.X(net7614),
    .A(net7615));
 sg13g2_buf_4 fanout7615 (.X(net7615),
    .A(net7616));
 sg13g2_buf_2 fanout7616 (.A(net7617),
    .X(net7616));
 sg13g2_buf_2 fanout7617 (.A(net7618),
    .X(net7617));
 sg13g2_buf_8 fanout7618 (.A(_12892_),
    .X(net7618));
 sg13g2_buf_4 fanout7619 (.X(net7619),
    .A(net7620));
 sg13g2_buf_2 fanout7620 (.A(net7624),
    .X(net7620));
 sg13g2_buf_4 fanout7621 (.X(net7621),
    .A(net7623));
 sg13g2_buf_4 fanout7622 (.X(net7622),
    .A(net7623));
 sg13g2_buf_2 fanout7623 (.A(net7624),
    .X(net7623));
 sg13g2_buf_4 fanout7624 (.X(net7624),
    .A(_12548_));
 sg13g2_buf_2 fanout7625 (.A(net7629),
    .X(net7625));
 sg13g2_buf_4 fanout7626 (.X(net7626),
    .A(net7629));
 sg13g2_buf_2 fanout7627 (.A(net7629),
    .X(net7627));
 sg13g2_buf_4 fanout7628 (.X(net7628),
    .A(net7629));
 sg13g2_buf_4 fanout7629 (.X(net7629),
    .A(_12539_));
 sg13g2_buf_4 fanout7630 (.X(net7630),
    .A(net7631));
 sg13g2_buf_2 fanout7631 (.A(net7632),
    .X(net7631));
 sg13g2_buf_2 fanout7632 (.A(net7635),
    .X(net7632));
 sg13g2_buf_4 fanout7633 (.X(net7633),
    .A(net7635));
 sg13g2_buf_2 fanout7634 (.A(net7635),
    .X(net7634));
 sg13g2_buf_2 fanout7635 (.A(_12530_),
    .X(net7635));
 sg13g2_buf_2 fanout7636 (.A(net7639),
    .X(net7636));
 sg13g2_buf_2 fanout7637 (.A(net7639),
    .X(net7637));
 sg13g2_buf_4 fanout7638 (.X(net7638),
    .A(net7639));
 sg13g2_buf_2 fanout7639 (.A(net7640),
    .X(net7639));
 sg13g2_buf_4 fanout7640 (.X(net7640),
    .A(net7641));
 sg13g2_buf_8 fanout7641 (.A(_12519_),
    .X(net7641));
 sg13g2_buf_2 fanout7642 (.A(net7645),
    .X(net7642));
 sg13g2_buf_2 fanout7643 (.A(net7644),
    .X(net7643));
 sg13g2_buf_2 fanout7644 (.A(net7645),
    .X(net7644));
 sg13g2_buf_2 fanout7645 (.A(net7646),
    .X(net7645));
 sg13g2_buf_4 fanout7646 (.X(net7646),
    .A(net7647));
 sg13g2_buf_8 fanout7647 (.A(_12509_),
    .X(net7647));
 sg13g2_buf_4 fanout7648 (.X(net7648),
    .A(net7652));
 sg13g2_buf_2 fanout7649 (.A(net7652),
    .X(net7649));
 sg13g2_buf_2 fanout7650 (.A(net7651),
    .X(net7650));
 sg13g2_buf_2 fanout7651 (.A(net7652),
    .X(net7651));
 sg13g2_buf_4 fanout7652 (.X(net7652),
    .A(_12497_));
 sg13g2_buf_2 fanout7653 (.A(net7656),
    .X(net7653));
 sg13g2_buf_2 fanout7654 (.A(net7655),
    .X(net7654));
 sg13g2_buf_4 fanout7655 (.X(net7655),
    .A(net7656));
 sg13g2_buf_2 fanout7656 (.A(net7657),
    .X(net7656));
 sg13g2_buf_4 fanout7657 (.X(net7657),
    .A(_12486_));
 sg13g2_buf_2 fanout7658 (.A(net7661),
    .X(net7658));
 sg13g2_buf_2 fanout7659 (.A(net7660),
    .X(net7659));
 sg13g2_buf_2 fanout7660 (.A(net7661),
    .X(net7660));
 sg13g2_buf_2 fanout7661 (.A(net7662),
    .X(net7661));
 sg13g2_buf_4 fanout7662 (.X(net7662),
    .A(_12477_));
 sg13g2_buf_4 fanout7663 (.X(net7663),
    .A(net7667));
 sg13g2_buf_4 fanout7664 (.X(net7664),
    .A(net7666));
 sg13g2_buf_2 fanout7665 (.A(net7666),
    .X(net7665));
 sg13g2_buf_2 fanout7666 (.A(net7667),
    .X(net7666));
 sg13g2_buf_2 fanout7667 (.A(net7668),
    .X(net7667));
 sg13g2_buf_8 fanout7668 (.A(_11846_),
    .X(net7668));
 sg13g2_buf_2 fanout7669 (.A(net7671),
    .X(net7669));
 sg13g2_buf_2 fanout7670 (.A(net7671),
    .X(net7670));
 sg13g2_buf_2 fanout7671 (.A(_11631_),
    .X(net7671));
 sg13g2_buf_2 fanout7672 (.A(net7674),
    .X(net7672));
 sg13g2_buf_2 fanout7673 (.A(net7674),
    .X(net7673));
 sg13g2_buf_2 fanout7674 (.A(_11624_),
    .X(net7674));
 sg13g2_buf_4 fanout7675 (.X(net7675),
    .A(_11630_));
 sg13g2_buf_4 fanout7676 (.X(net7676),
    .A(_11629_));
 sg13g2_buf_4 fanout7677 (.X(net7677),
    .A(_11623_));
 sg13g2_buf_2 fanout7678 (.A(_11623_),
    .X(net7678));
 sg13g2_buf_4 fanout7679 (.X(net7679),
    .A(_11618_));
 sg13g2_buf_2 fanout7680 (.A(_11618_),
    .X(net7680));
 sg13g2_buf_2 fanout7681 (.A(net7682),
    .X(net7681));
 sg13g2_buf_2 fanout7682 (.A(_06611_),
    .X(net7682));
 sg13g2_buf_2 fanout7683 (.A(net7684),
    .X(net7683));
 sg13g2_buf_2 fanout7684 (.A(_06222_),
    .X(net7684));
 sg13g2_buf_4 fanout7685 (.X(net7685),
    .A(net7687));
 sg13g2_buf_8 fanout7686 (.A(net7687),
    .X(net7686));
 sg13g2_buf_4 fanout7687 (.X(net7687),
    .A(_12612_));
 sg13g2_buf_4 fanout7688 (.X(net7688),
    .A(net7689));
 sg13g2_buf_8 fanout7689 (.A(_12612_),
    .X(net7689));
 sg13g2_buf_4 fanout7690 (.X(net7690),
    .A(net7695));
 sg13g2_buf_2 fanout7691 (.A(net7695),
    .X(net7691));
 sg13g2_buf_4 fanout7692 (.X(net7692),
    .A(net7693));
 sg13g2_buf_2 fanout7693 (.A(net7694),
    .X(net7693));
 sg13g2_buf_4 fanout7694 (.X(net7694),
    .A(net7695));
 sg13g2_buf_2 fanout7695 (.A(_08182_),
    .X(net7695));
 sg13g2_buf_4 fanout7696 (.X(net7696),
    .A(net7697));
 sg13g2_buf_8 fanout7697 (.A(net7700),
    .X(net7697));
 sg13g2_buf_8 fanout7698 (.A(net7700),
    .X(net7698));
 sg13g2_buf_4 fanout7699 (.X(net7699),
    .A(net7700));
 sg13g2_buf_4 fanout7700 (.X(net7700),
    .A(_04075_));
 sg13g2_buf_4 fanout7701 (.X(net7701),
    .A(net7702));
 sg13g2_buf_4 fanout7702 (.X(net7702),
    .A(_03854_));
 sg13g2_buf_4 fanout7703 (.X(net7703),
    .A(net7704));
 sg13g2_buf_4 fanout7704 (.X(net7704),
    .A(_03854_));
 sg13g2_buf_4 fanout7705 (.X(net7705),
    .A(net7706));
 sg13g2_buf_4 fanout7706 (.X(net7706),
    .A(_03853_));
 sg13g2_buf_4 fanout7707 (.X(net7707),
    .A(net7708));
 sg13g2_buf_4 fanout7708 (.X(net7708),
    .A(net7709));
 sg13g2_buf_4 fanout7709 (.X(net7709),
    .A(_08181_));
 sg13g2_buf_4 fanout7710 (.X(net7710),
    .A(_07483_));
 sg13g2_buf_2 fanout7711 (.A(_07483_),
    .X(net7711));
 sg13g2_buf_4 fanout7712 (.X(net7712),
    .A(_07483_));
 sg13g2_buf_2 fanout7713 (.A(net7714),
    .X(net7713));
 sg13g2_buf_4 fanout7714 (.X(net7714),
    .A(net7718));
 sg13g2_buf_2 fanout7715 (.A(net7717),
    .X(net7715));
 sg13g2_buf_2 fanout7716 (.A(net7717),
    .X(net7716));
 sg13g2_buf_4 fanout7717 (.X(net7717),
    .A(net7718));
 sg13g2_buf_4 fanout7718 (.X(net7718),
    .A(net7722));
 sg13g2_buf_4 fanout7719 (.X(net7719),
    .A(net7722));
 sg13g2_buf_2 fanout7720 (.A(net7722),
    .X(net7720));
 sg13g2_buf_2 fanout7721 (.A(net7722),
    .X(net7721));
 sg13g2_buf_4 fanout7722 (.X(net7722),
    .A(_04560_));
 sg13g2_buf_2 fanout7723 (.A(net7725),
    .X(net7723));
 sg13g2_buf_1 fanout7724 (.A(net7725),
    .X(net7724));
 sg13g2_buf_2 fanout7725 (.A(net7729),
    .X(net7725));
 sg13g2_buf_2 fanout7726 (.A(net7728),
    .X(net7726));
 sg13g2_buf_2 fanout7727 (.A(net7728),
    .X(net7727));
 sg13g2_buf_2 fanout7728 (.A(net7729),
    .X(net7728));
 sg13g2_buf_2 fanout7729 (.A(_04185_),
    .X(net7729));
 sg13g2_buf_2 fanout7730 (.A(net7733),
    .X(net7730));
 sg13g2_buf_2 fanout7731 (.A(net7733),
    .X(net7731));
 sg13g2_buf_4 fanout7732 (.X(net7732),
    .A(net7733));
 sg13g2_buf_4 fanout7733 (.X(net7733),
    .A(_04185_));
 sg13g2_buf_4 fanout7734 (.X(net7734),
    .A(net7737));
 sg13g2_buf_2 fanout7735 (.A(net7737),
    .X(net7735));
 sg13g2_buf_4 fanout7736 (.X(net7736),
    .A(net7737));
 sg13g2_buf_8 fanout7737 (.A(_04121_),
    .X(net7737));
 sg13g2_buf_4 fanout7738 (.X(net7738),
    .A(net7741));
 sg13g2_buf_2 fanout7739 (.A(net7741),
    .X(net7739));
 sg13g2_buf_4 fanout7740 (.X(net7740),
    .A(net7741));
 sg13g2_buf_4 fanout7741 (.X(net7741),
    .A(_04120_));
 sg13g2_buf_4 fanout7742 (.X(net7742),
    .A(net7743));
 sg13g2_buf_4 fanout7743 (.X(net7743),
    .A(net7746));
 sg13g2_buf_2 fanout7744 (.A(net7745),
    .X(net7744));
 sg13g2_buf_4 fanout7745 (.X(net7745),
    .A(net7746));
 sg13g2_buf_2 fanout7746 (.A(_04074_),
    .X(net7746));
 sg13g2_buf_4 fanout7747 (.X(net7747),
    .A(net7748));
 sg13g2_buf_4 fanout7748 (.X(net7748),
    .A(_03852_));
 sg13g2_buf_2 fanout7749 (.A(net7756),
    .X(net7749));
 sg13g2_buf_2 fanout7750 (.A(net7756),
    .X(net7750));
 sg13g2_buf_2 fanout7751 (.A(net7756),
    .X(net7751));
 sg13g2_buf_2 fanout7752 (.A(net7753),
    .X(net7752));
 sg13g2_buf_2 fanout7753 (.A(net7756),
    .X(net7753));
 sg13g2_buf_4 fanout7754 (.X(net7754),
    .A(net7756));
 sg13g2_buf_2 fanout7755 (.A(net7756),
    .X(net7755));
 sg13g2_buf_4 fanout7756 (.X(net7756),
    .A(_07482_));
 sg13g2_buf_4 fanout7757 (.X(net7757),
    .A(net7761));
 sg13g2_buf_4 fanout7758 (.X(net7758),
    .A(net7759));
 sg13g2_buf_4 fanout7759 (.X(net7759),
    .A(net7760));
 sg13g2_buf_4 fanout7760 (.X(net7760),
    .A(net7761));
 sg13g2_buf_2 fanout7761 (.A(_05303_),
    .X(net7761));
 sg13g2_buf_4 fanout7762 (.X(net7762),
    .A(net7771));
 sg13g2_buf_2 fanout7763 (.A(net7766),
    .X(net7763));
 sg13g2_buf_1 fanout7764 (.A(net7766),
    .X(net7764));
 sg13g2_buf_2 fanout7765 (.A(net7766),
    .X(net7765));
 sg13g2_buf_2 fanout7766 (.A(net7771),
    .X(net7766));
 sg13g2_buf_2 fanout7767 (.A(net7770),
    .X(net7767));
 sg13g2_buf_2 fanout7768 (.A(net7770),
    .X(net7768));
 sg13g2_buf_2 fanout7769 (.A(net7770),
    .X(net7769));
 sg13g2_buf_4 fanout7770 (.X(net7770),
    .A(net7771));
 sg13g2_buf_4 fanout7771 (.X(net7771),
    .A(_04593_));
 sg13g2_buf_2 fanout7772 (.A(net7777),
    .X(net7772));
 sg13g2_buf_4 fanout7773 (.X(net7773),
    .A(net7777));
 sg13g2_buf_2 fanout7774 (.A(net7776),
    .X(net7774));
 sg13g2_buf_2 fanout7775 (.A(net7776),
    .X(net7775));
 sg13g2_buf_4 fanout7776 (.X(net7776),
    .A(net7777));
 sg13g2_buf_4 fanout7777 (.X(net7777),
    .A(net7781));
 sg13g2_buf_2 fanout7778 (.A(net7781),
    .X(net7778));
 sg13g2_buf_2 fanout7779 (.A(net7781),
    .X(net7779));
 sg13g2_buf_2 fanout7780 (.A(net7781),
    .X(net7780));
 sg13g2_buf_4 fanout7781 (.X(net7781),
    .A(_04218_));
 sg13g2_buf_4 fanout7782 (.X(net7782),
    .A(net7787));
 sg13g2_buf_2 fanout7783 (.A(net7784),
    .X(net7783));
 sg13g2_buf_8 fanout7784 (.A(net7787),
    .X(net7784));
 sg13g2_buf_8 fanout7785 (.A(net7787),
    .X(net7785));
 sg13g2_buf_2 fanout7786 (.A(net7787),
    .X(net7786));
 sg13g2_buf_4 fanout7787 (.X(net7787),
    .A(_12623_));
 sg13g2_buf_4 fanout7788 (.X(net7788),
    .A(net7789));
 sg13g2_buf_4 fanout7789 (.X(net7789),
    .A(net7792));
 sg13g2_buf_4 fanout7790 (.X(net7790),
    .A(net7791));
 sg13g2_buf_8 fanout7791 (.A(net7792),
    .X(net7791));
 sg13g2_buf_8 fanout7792 (.A(_12621_),
    .X(net7792));
 sg13g2_buf_4 fanout7793 (.X(net7793),
    .A(net7794));
 sg13g2_buf_4 fanout7794 (.X(net7794),
    .A(net7797));
 sg13g2_buf_2 fanout7795 (.A(net7797),
    .X(net7795));
 sg13g2_buf_4 fanout7796 (.X(net7796),
    .A(net7797));
 sg13g2_buf_8 fanout7797 (.A(_12620_),
    .X(net7797));
 sg13g2_buf_4 fanout7798 (.X(net7798),
    .A(net7801));
 sg13g2_buf_4 fanout7799 (.X(net7799),
    .A(net7801));
 sg13g2_buf_2 fanout7800 (.A(net7801),
    .X(net7800));
 sg13g2_buf_4 fanout7801 (.X(net7801),
    .A(_12619_));
 sg13g2_buf_4 fanout7802 (.X(net7802),
    .A(net7806));
 sg13g2_buf_2 fanout7803 (.A(net7804),
    .X(net7803));
 sg13g2_buf_2 fanout7804 (.A(net7805),
    .X(net7804));
 sg13g2_buf_4 fanout7805 (.X(net7805),
    .A(net7806));
 sg13g2_buf_2 fanout7806 (.A(_12619_),
    .X(net7806));
 sg13g2_buf_4 fanout7807 (.X(net7807),
    .A(net7810));
 sg13g2_buf_4 fanout7808 (.X(net7808),
    .A(net7810));
 sg13g2_buf_2 fanout7809 (.A(net7810),
    .X(net7809));
 sg13g2_buf_2 fanout7810 (.A(_12616_),
    .X(net7810));
 sg13g2_buf_4 fanout7811 (.X(net7811),
    .A(_12616_));
 sg13g2_buf_2 fanout7812 (.A(_12616_),
    .X(net7812));
 sg13g2_buf_4 fanout7813 (.X(net7813),
    .A(net7815));
 sg13g2_buf_2 fanout7814 (.A(net7815),
    .X(net7814));
 sg13g2_buf_4 fanout7815 (.X(net7815),
    .A(net7816));
 sg13g2_buf_4 fanout7816 (.X(net7816),
    .A(net7823));
 sg13g2_buf_4 fanout7817 (.X(net7817),
    .A(net7821));
 sg13g2_buf_4 fanout7818 (.X(net7818),
    .A(net7821));
 sg13g2_buf_2 fanout7819 (.A(net7820),
    .X(net7819));
 sg13g2_buf_4 fanout7820 (.X(net7820),
    .A(net7821));
 sg13g2_buf_2 fanout7821 (.A(net7823),
    .X(net7821));
 sg13g2_buf_4 fanout7822 (.X(net7822),
    .A(net7823));
 sg13g2_buf_8 fanout7823 (.A(_09124_),
    .X(net7823));
 sg13g2_buf_4 fanout7824 (.X(net7824),
    .A(net7825));
 sg13g2_buf_4 fanout7825 (.X(net7825),
    .A(net7826));
 sg13g2_buf_4 fanout7826 (.X(net7826),
    .A(net7827));
 sg13g2_buf_4 fanout7827 (.X(net7827),
    .A(net7834));
 sg13g2_buf_4 fanout7828 (.X(net7828),
    .A(net7834));
 sg13g2_buf_1 fanout7829 (.A(net7834),
    .X(net7829));
 sg13g2_buf_4 fanout7830 (.X(net7830),
    .A(net7832));
 sg13g2_buf_4 fanout7831 (.X(net7831),
    .A(net7832));
 sg13g2_buf_4 fanout7832 (.X(net7832),
    .A(net7833));
 sg13g2_buf_4 fanout7833 (.X(net7833),
    .A(net7834));
 sg13g2_buf_4 fanout7834 (.X(net7834),
    .A(_08792_));
 sg13g2_buf_4 fanout7835 (.X(net7835),
    .A(net7837));
 sg13g2_buf_2 fanout7836 (.A(net7837),
    .X(net7836));
 sg13g2_buf_2 fanout7837 (.A(net7838),
    .X(net7837));
 sg13g2_buf_2 fanout7838 (.A(net7839),
    .X(net7838));
 sg13g2_buf_4 fanout7839 (.X(net7839),
    .A(_08759_));
 sg13g2_buf_4 fanout7840 (.X(net7840),
    .A(net7845));
 sg13g2_buf_1 fanout7841 (.A(net7845),
    .X(net7841));
 sg13g2_buf_4 fanout7842 (.X(net7842),
    .A(net7843));
 sg13g2_buf_8 fanout7843 (.A(net7844),
    .X(net7843));
 sg13g2_buf_8 fanout7844 (.A(net7845),
    .X(net7844));
 sg13g2_buf_8 fanout7845 (.A(_08759_),
    .X(net7845));
 sg13g2_buf_4 fanout7846 (.X(net7846),
    .A(net7848));
 sg13g2_buf_1 fanout7847 (.A(net7848),
    .X(net7847));
 sg13g2_buf_4 fanout7848 (.X(net7848),
    .A(net7850));
 sg13g2_buf_4 fanout7849 (.X(net7849),
    .A(net7850));
 sg13g2_buf_4 fanout7850 (.X(net7850),
    .A(net7856));
 sg13g2_buf_4 fanout7851 (.X(net7851),
    .A(net7853));
 sg13g2_buf_4 fanout7852 (.X(net7852),
    .A(net7853));
 sg13g2_buf_4 fanout7853 (.X(net7853),
    .A(net7856));
 sg13g2_buf_4 fanout7854 (.X(net7854),
    .A(net7856));
 sg13g2_buf_4 fanout7855 (.X(net7855),
    .A(net7856));
 sg13g2_buf_8 fanout7856 (.A(_08688_),
    .X(net7856));
 sg13g2_buf_4 fanout7857 (.X(net7857),
    .A(net7858));
 sg13g2_buf_4 fanout7858 (.X(net7858),
    .A(net7859));
 sg13g2_buf_4 fanout7859 (.X(net7859),
    .A(net7860));
 sg13g2_buf_8 fanout7860 (.A(net7867),
    .X(net7860));
 sg13g2_buf_4 fanout7861 (.X(net7861),
    .A(net7866));
 sg13g2_buf_2 fanout7862 (.A(net7866),
    .X(net7862));
 sg13g2_buf_4 fanout7863 (.X(net7863),
    .A(net7866));
 sg13g2_buf_4 fanout7864 (.X(net7864),
    .A(net7866));
 sg13g2_buf_4 fanout7865 (.X(net7865),
    .A(net7867));
 sg13g2_buf_2 fanout7866 (.A(net7867),
    .X(net7866));
 sg13g2_buf_8 fanout7867 (.A(_08655_),
    .X(net7867));
 sg13g2_buf_4 fanout7868 (.X(net7868),
    .A(net7869));
 sg13g2_buf_4 fanout7869 (.X(net7869),
    .A(net7870));
 sg13g2_buf_4 fanout7870 (.X(net7870),
    .A(net7871));
 sg13g2_buf_4 fanout7871 (.X(net7871),
    .A(_06086_));
 sg13g2_buf_4 fanout7872 (.X(net7872),
    .A(net7877));
 sg13g2_buf_1 fanout7873 (.A(net7877),
    .X(net7873));
 sg13g2_buf_4 fanout7874 (.X(net7874),
    .A(net7875));
 sg13g2_buf_8 fanout7875 (.A(net7876),
    .X(net7875));
 sg13g2_buf_8 fanout7876 (.A(net7877),
    .X(net7876));
 sg13g2_buf_8 fanout7877 (.A(_06086_),
    .X(net7877));
 sg13g2_buf_2 fanout7878 (.A(net7879),
    .X(net7878));
 sg13g2_buf_2 fanout7879 (.A(_05302_),
    .X(net7879));
 sg13g2_buf_2 fanout7880 (.A(net7881),
    .X(net7880));
 sg13g2_buf_2 fanout7881 (.A(net7882),
    .X(net7881));
 sg13g2_buf_4 fanout7882 (.X(net7882),
    .A(_05302_));
 sg13g2_buf_4 fanout7883 (.X(net7883),
    .A(net7884));
 sg13g2_buf_2 fanout7884 (.A(net7885),
    .X(net7884));
 sg13g2_buf_4 fanout7885 (.X(net7885),
    .A(net7886));
 sg13g2_buf_4 fanout7886 (.X(net7886),
    .A(_03743_));
 sg13g2_buf_4 fanout7887 (.X(net7887),
    .A(net7892));
 sg13g2_buf_2 fanout7888 (.A(net7892),
    .X(net7888));
 sg13g2_buf_4 fanout7889 (.X(net7889),
    .A(net7890));
 sg13g2_buf_4 fanout7890 (.X(net7890),
    .A(net7891));
 sg13g2_buf_4 fanout7891 (.X(net7891),
    .A(net7892));
 sg13g2_buf_8 fanout7892 (.A(_03743_),
    .X(net7892));
 sg13g2_buf_4 fanout7893 (.X(net7893),
    .A(net7895));
 sg13g2_buf_2 fanout7894 (.A(net7895),
    .X(net7894));
 sg13g2_buf_4 fanout7895 (.X(net7895),
    .A(net7896));
 sg13g2_buf_2 fanout7896 (.A(net7897),
    .X(net7896));
 sg13g2_buf_8 fanout7897 (.A(net7903),
    .X(net7897));
 sg13g2_buf_4 fanout7898 (.X(net7898),
    .A(net7900));
 sg13g2_buf_4 fanout7899 (.X(net7899),
    .A(net7900));
 sg13g2_buf_4 fanout7900 (.X(net7900),
    .A(net7903));
 sg13g2_buf_4 fanout7901 (.X(net7901),
    .A(net7903));
 sg13g2_buf_4 fanout7902 (.X(net7902),
    .A(net7903));
 sg13g2_buf_8 fanout7903 (.A(_14371_),
    .X(net7903));
 sg13g2_buf_4 fanout7904 (.X(net7904),
    .A(net7907));
 sg13g2_buf_4 fanout7905 (.X(net7905),
    .A(net7907));
 sg13g2_buf_2 fanout7906 (.A(net7907),
    .X(net7906));
 sg13g2_buf_2 fanout7907 (.A(_12617_),
    .X(net7907));
 sg13g2_buf_8 fanout7908 (.A(_12617_),
    .X(net7908));
 sg13g2_buf_2 fanout7909 (.A(_12617_),
    .X(net7909));
 sg13g2_buf_4 fanout7910 (.X(net7910),
    .A(net7913));
 sg13g2_buf_4 fanout7911 (.X(net7911),
    .A(net7912));
 sg13g2_buf_4 fanout7912 (.X(net7912),
    .A(net7913));
 sg13g2_buf_4 fanout7913 (.X(net7913),
    .A(net7914));
 sg13g2_buf_8 fanout7914 (.A(_12598_),
    .X(net7914));
 sg13g2_buf_4 fanout7915 (.X(net7915),
    .A(net7916));
 sg13g2_buf_4 fanout7916 (.X(net7916),
    .A(net7917));
 sg13g2_buf_8 fanout7917 (.A(_12597_),
    .X(net7917));
 sg13g2_buf_8 fanout7918 (.A(_12597_),
    .X(net7918));
 sg13g2_buf_2 fanout7919 (.A(_12597_),
    .X(net7919));
 sg13g2_buf_4 fanout7920 (.X(net7920),
    .A(net7921));
 sg13g2_buf_4 fanout7921 (.X(net7921),
    .A(net7922));
 sg13g2_buf_8 fanout7922 (.A(net7924),
    .X(net7922));
 sg13g2_buf_8 fanout7923 (.A(net7924),
    .X(net7923));
 sg13g2_buf_8 fanout7924 (.A(_12593_),
    .X(net7924));
 sg13g2_buf_4 fanout7925 (.X(net7925),
    .A(net7930));
 sg13g2_buf_2 fanout7926 (.A(net7927),
    .X(net7926));
 sg13g2_buf_4 fanout7927 (.X(net7927),
    .A(net7930));
 sg13g2_buf_8 fanout7928 (.A(net7930),
    .X(net7928));
 sg13g2_buf_4 fanout7929 (.X(net7929),
    .A(net7930));
 sg13g2_buf_8 fanout7930 (.A(_12589_),
    .X(net7930));
 sg13g2_buf_4 fanout7931 (.X(net7931),
    .A(net7932));
 sg13g2_buf_4 fanout7932 (.X(net7932),
    .A(net7933));
 sg13g2_buf_4 fanout7933 (.X(net7933),
    .A(net7935));
 sg13g2_buf_8 fanout7934 (.A(net7935),
    .X(net7934));
 sg13g2_buf_8 fanout7935 (.A(_12583_),
    .X(net7935));
 sg13g2_buf_2 fanout7936 (.A(net7937),
    .X(net7936));
 sg13g2_buf_2 fanout7937 (.A(_11939_),
    .X(net7937));
 sg13g2_buf_2 fanout7938 (.A(_11895_),
    .X(net7938));
 sg13g2_buf_4 fanout7939 (.X(net7939),
    .A(net7941));
 sg13g2_buf_4 fanout7940 (.X(net7940),
    .A(net7941));
 sg13g2_buf_4 fanout7941 (.X(net7941),
    .A(net7942));
 sg13g2_buf_4 fanout7942 (.X(net7942),
    .A(_10342_));
 sg13g2_buf_4 fanout7943 (.X(net7943),
    .A(net7948));
 sg13g2_buf_4 fanout7944 (.X(net7944),
    .A(net7946));
 sg13g2_buf_2 fanout7945 (.A(net7946),
    .X(net7945));
 sg13g2_buf_4 fanout7946 (.X(net7946),
    .A(net7948));
 sg13g2_buf_4 fanout7947 (.X(net7947),
    .A(net7948));
 sg13g2_buf_8 fanout7948 (.A(_10342_),
    .X(net7948));
 sg13g2_buf_4 fanout7949 (.X(net7949),
    .A(net7950));
 sg13g2_buf_4 fanout7950 (.X(net7950),
    .A(net7951));
 sg13g2_buf_4 fanout7951 (.X(net7951),
    .A(net7952));
 sg13g2_buf_8 fanout7952 (.A(net7958),
    .X(net7952));
 sg13g2_buf_4 fanout7953 (.X(net7953),
    .A(net7958));
 sg13g2_buf_4 fanout7954 (.X(net7954),
    .A(net7956));
 sg13g2_buf_4 fanout7955 (.X(net7955),
    .A(net7956));
 sg13g2_buf_4 fanout7956 (.X(net7956),
    .A(net7958));
 sg13g2_buf_4 fanout7957 (.X(net7957),
    .A(net7958));
 sg13g2_buf_8 fanout7958 (.A(_10309_),
    .X(net7958));
 sg13g2_buf_4 fanout7959 (.X(net7959),
    .A(net7960));
 sg13g2_buf_4 fanout7960 (.X(net7960),
    .A(net7961));
 sg13g2_buf_8 fanout7961 (.A(net7969),
    .X(net7961));
 sg13g2_buf_2 fanout7962 (.A(net7969),
    .X(net7962));
 sg13g2_buf_4 fanout7963 (.X(net7963),
    .A(net7969));
 sg13g2_buf_2 fanout7964 (.A(net7969),
    .X(net7964));
 sg13g2_buf_4 fanout7965 (.X(net7965),
    .A(net7967));
 sg13g2_buf_4 fanout7966 (.X(net7966),
    .A(net7967));
 sg13g2_buf_4 fanout7967 (.X(net7967),
    .A(net7968));
 sg13g2_buf_8 fanout7968 (.A(net7969),
    .X(net7968));
 sg13g2_buf_8 fanout7969 (.A(_08925_),
    .X(net7969));
 sg13g2_buf_2 fanout7970 (.A(net7971),
    .X(net7970));
 sg13g2_buf_2 fanout7971 (.A(net7972),
    .X(net7971));
 sg13g2_buf_4 fanout7972 (.X(net7972),
    .A(_05653_));
 sg13g2_buf_2 fanout7973 (.A(net7975),
    .X(net7973));
 sg13g2_buf_2 fanout7974 (.A(net7975),
    .X(net7974));
 sg13g2_buf_2 fanout7975 (.A(net7976),
    .X(net7975));
 sg13g2_buf_2 fanout7976 (.A(_05652_),
    .X(net7976));
 sg13g2_buf_2 fanout7977 (.A(net7978),
    .X(net7977));
 sg13g2_buf_2 fanout7978 (.A(net7979),
    .X(net7978));
 sg13g2_buf_2 fanout7979 (.A(_05652_),
    .X(net7979));
 sg13g2_buf_2 fanout7980 (.A(net7981),
    .X(net7980));
 sg13g2_buf_4 fanout7981 (.X(net7981),
    .A(net7982));
 sg13g2_buf_4 fanout7982 (.X(net7982),
    .A(_05038_));
 sg13g2_buf_2 fanout7983 (.A(net7985),
    .X(net7983));
 sg13g2_buf_1 fanout7984 (.A(net7985),
    .X(net7984));
 sg13g2_buf_2 fanout7985 (.A(net7986),
    .X(net7985));
 sg13g2_buf_2 fanout7986 (.A(_05037_),
    .X(net7986));
 sg13g2_buf_2 fanout7987 (.A(net7988),
    .X(net7987));
 sg13g2_buf_2 fanout7988 (.A(net7989),
    .X(net7988));
 sg13g2_buf_2 fanout7989 (.A(_05037_),
    .X(net7989));
 sg13g2_buf_4 fanout7990 (.X(net7990),
    .A(_03850_));
 sg13g2_buf_2 fanout7991 (.A(_03850_),
    .X(net7991));
 sg13g2_buf_2 fanout7992 (.A(net7993),
    .X(net7992));
 sg13g2_buf_4 fanout7993 (.X(net7993),
    .A(_03850_));
 sg13g2_buf_4 fanout7994 (.X(net7994),
    .A(_11661_));
 sg13g2_buf_4 fanout7995 (.X(net7995),
    .A(_11660_));
 sg13g2_buf_2 fanout7996 (.A(net7997),
    .X(net7996));
 sg13g2_buf_2 fanout7997 (.A(net7999),
    .X(net7997));
 sg13g2_buf_4 fanout7998 (.X(net7998),
    .A(net7999));
 sg13g2_buf_4 fanout7999 (.X(net7999),
    .A(_11643_));
 sg13g2_buf_2 fanout8000 (.A(net8001),
    .X(net8000));
 sg13g2_buf_1 fanout8001 (.A(net8003),
    .X(net8001));
 sg13g2_buf_4 fanout8002 (.X(net8002),
    .A(net8003));
 sg13g2_buf_2 fanout8003 (.A(_11639_),
    .X(net8003));
 sg13g2_buf_4 fanout8004 (.X(net8004),
    .A(_11635_));
 sg13g2_buf_2 fanout8005 (.A(_11635_),
    .X(net8005));
 sg13g2_buf_4 fanout8006 (.X(net8006),
    .A(_11442_));
 sg13g2_buf_4 fanout8007 (.X(net8007),
    .A(_11080_));
 sg13g2_buf_4 fanout8008 (.X(net8008),
    .A(_11070_));
 sg13g2_buf_2 fanout8009 (.A(net8010),
    .X(net8009));
 sg13g2_buf_4 fanout8010 (.X(net8010),
    .A(net8012));
 sg13g2_buf_4 fanout8011 (.X(net8011),
    .A(net8012));
 sg13g2_buf_8 fanout8012 (.A(_09157_),
    .X(net8012));
 sg13g2_buf_4 fanout8013 (.X(net8013),
    .A(net8019));
 sg13g2_buf_4 fanout8014 (.X(net8014),
    .A(net8019));
 sg13g2_buf_4 fanout8015 (.X(net8015),
    .A(net8017));
 sg13g2_buf_2 fanout8016 (.A(net8017),
    .X(net8016));
 sg13g2_buf_8 fanout8017 (.A(net8019),
    .X(net8017));
 sg13g2_buf_4 fanout8018 (.X(net8018),
    .A(net8019));
 sg13g2_buf_4 fanout8019 (.X(net8019),
    .A(_09157_));
 sg13g2_buf_4 fanout8020 (.X(net8020),
    .A(net8021));
 sg13g2_buf_4 fanout8021 (.X(net8021),
    .A(net8022));
 sg13g2_buf_8 fanout8022 (.A(_09091_),
    .X(net8022));
 sg13g2_buf_2 fanout8023 (.A(_09091_),
    .X(net8023));
 sg13g2_buf_4 fanout8024 (.X(net8024),
    .A(net8029));
 sg13g2_buf_4 fanout8025 (.X(net8025),
    .A(net8026));
 sg13g2_buf_2 fanout8026 (.A(net8029),
    .X(net8026));
 sg13g2_buf_4 fanout8027 (.X(net8027),
    .A(net8029));
 sg13g2_buf_4 fanout8028 (.X(net8028),
    .A(net8029));
 sg13g2_buf_8 fanout8029 (.A(_09091_),
    .X(net8029));
 sg13g2_buf_4 fanout8030 (.X(net8030),
    .A(net8032));
 sg13g2_buf_2 fanout8031 (.A(net8032),
    .X(net8031));
 sg13g2_buf_4 fanout8032 (.X(net8032),
    .A(net8034));
 sg13g2_buf_4 fanout8033 (.X(net8033),
    .A(net8034));
 sg13g2_buf_4 fanout8034 (.X(net8034),
    .A(_08891_));
 sg13g2_buf_4 fanout8035 (.X(net8035),
    .A(net8041));
 sg13g2_buf_2 fanout8036 (.A(net8041),
    .X(net8036));
 sg13g2_buf_4 fanout8037 (.X(net8037),
    .A(net8039));
 sg13g2_buf_2 fanout8038 (.A(net8039),
    .X(net8038));
 sg13g2_buf_4 fanout8039 (.X(net8039),
    .A(net8041));
 sg13g2_buf_4 fanout8040 (.X(net8040),
    .A(net8041));
 sg13g2_buf_8 fanout8041 (.A(_08891_),
    .X(net8041));
 sg13g2_buf_4 fanout8042 (.X(net8042),
    .A(net8043));
 sg13g2_buf_4 fanout8043 (.X(net8043),
    .A(net8045));
 sg13g2_buf_4 fanout8044 (.X(net8044),
    .A(net8045));
 sg13g2_buf_8 fanout8045 (.A(_08858_),
    .X(net8045));
 sg13g2_buf_4 fanout8046 (.X(net8046),
    .A(net8052));
 sg13g2_buf_2 fanout8047 (.A(net8052),
    .X(net8047));
 sg13g2_buf_2 fanout8048 (.A(net8050),
    .X(net8048));
 sg13g2_buf_2 fanout8049 (.A(net8050),
    .X(net8049));
 sg13g2_buf_4 fanout8050 (.X(net8050),
    .A(net8052));
 sg13g2_buf_4 fanout8051 (.X(net8051),
    .A(net8052));
 sg13g2_buf_4 fanout8052 (.X(net8052),
    .A(_08858_));
 sg13g2_buf_2 fanout8053 (.A(net8054),
    .X(net8053));
 sg13g2_buf_4 fanout8054 (.X(net8054),
    .A(net8056));
 sg13g2_buf_4 fanout8055 (.X(net8055),
    .A(net8056));
 sg13g2_buf_8 fanout8056 (.A(_08825_),
    .X(net8056));
 sg13g2_buf_8 fanout8057 (.A(net8063),
    .X(net8057));
 sg13g2_buf_2 fanout8058 (.A(net8063),
    .X(net8058));
 sg13g2_buf_2 fanout8059 (.A(net8061),
    .X(net8059));
 sg13g2_buf_2 fanout8060 (.A(net8061),
    .X(net8060));
 sg13g2_buf_4 fanout8061 (.X(net8061),
    .A(net8063));
 sg13g2_buf_2 fanout8062 (.A(net8063),
    .X(net8062));
 sg13g2_buf_4 fanout8063 (.X(net8063),
    .A(_08825_));
 sg13g2_buf_4 fanout8064 (.X(net8064),
    .A(net8065));
 sg13g2_buf_4 fanout8065 (.X(net8065),
    .A(net8067));
 sg13g2_buf_4 fanout8066 (.X(net8066),
    .A(net8067));
 sg13g2_buf_8 fanout8067 (.A(net8075),
    .X(net8067));
 sg13g2_buf_4 fanout8068 (.X(net8068),
    .A(net8075));
 sg13g2_buf_2 fanout8069 (.A(net8075),
    .X(net8069));
 sg13g2_buf_4 fanout8070 (.X(net8070),
    .A(net8074));
 sg13g2_buf_4 fanout8071 (.X(net8071),
    .A(net8073));
 sg13g2_buf_2 fanout8072 (.A(net8073),
    .X(net8072));
 sg13g2_buf_4 fanout8073 (.X(net8073),
    .A(net8074));
 sg13g2_buf_4 fanout8074 (.X(net8074),
    .A(net8075));
 sg13g2_buf_8 fanout8075 (.A(_08726_),
    .X(net8075));
 sg13g2_buf_4 fanout8076 (.X(net8076),
    .A(net8078));
 sg13g2_buf_4 fanout8077 (.X(net8077),
    .A(net8078));
 sg13g2_buf_2 fanout8078 (.A(net8079),
    .X(net8078));
 sg13g2_buf_4 fanout8079 (.X(net8079),
    .A(_07143_));
 sg13g2_buf_4 fanout8080 (.X(net8080),
    .A(net8085));
 sg13g2_buf_4 fanout8081 (.X(net8081),
    .A(net8082));
 sg13g2_buf_4 fanout8082 (.X(net8082),
    .A(net8083));
 sg13g2_buf_4 fanout8083 (.X(net8083),
    .A(net8085));
 sg13g2_buf_4 fanout8084 (.X(net8084),
    .A(net8085));
 sg13g2_buf_8 fanout8085 (.A(_07143_),
    .X(net8085));
 sg13g2_buf_4 fanout8086 (.X(net8086),
    .A(net8087));
 sg13g2_buf_2 fanout8087 (.A(net8088),
    .X(net8087));
 sg13g2_buf_4 fanout8088 (.X(net8088),
    .A(net8096));
 sg13g2_buf_4 fanout8089 (.X(net8089),
    .A(net8096));
 sg13g2_buf_4 fanout8090 (.X(net8090),
    .A(net8095));
 sg13g2_buf_4 fanout8091 (.X(net8091),
    .A(net8092));
 sg13g2_buf_2 fanout8092 (.A(net8094),
    .X(net8092));
 sg13g2_buf_4 fanout8093 (.X(net8093),
    .A(net8094));
 sg13g2_buf_4 fanout8094 (.X(net8094),
    .A(net8095));
 sg13g2_buf_4 fanout8095 (.X(net8095),
    .A(net8096));
 sg13g2_buf_4 fanout8096 (.X(net8096),
    .A(_07003_));
 sg13g2_buf_4 fanout8097 (.X(net8097),
    .A(net8099));
 sg13g2_buf_2 fanout8098 (.A(net8099),
    .X(net8098));
 sg13g2_buf_4 fanout8099 (.X(net8099),
    .A(net8100));
 sg13g2_buf_4 fanout8100 (.X(net8100),
    .A(net8107));
 sg13g2_buf_4 fanout8101 (.X(net8101),
    .A(net8107));
 sg13g2_buf_1 fanout8102 (.A(net8107),
    .X(net8102));
 sg13g2_buf_4 fanout8103 (.X(net8103),
    .A(net8105));
 sg13g2_buf_4 fanout8104 (.X(net8104),
    .A(net8105));
 sg13g2_buf_4 fanout8105 (.X(net8105),
    .A(net8106));
 sg13g2_buf_4 fanout8106 (.X(net8106),
    .A(net8107));
 sg13g2_buf_8 fanout8107 (.A(_06464_),
    .X(net8107));
 sg13g2_buf_4 fanout8108 (.X(net8108),
    .A(net8109));
 sg13g2_buf_2 fanout8109 (.A(net8110),
    .X(net8109));
 sg13g2_buf_4 fanout8110 (.X(net8110),
    .A(net8111));
 sg13g2_buf_4 fanout8111 (.X(net8111),
    .A(_04617_));
 sg13g2_buf_4 fanout8112 (.X(net8112),
    .A(net8118));
 sg13g2_buf_4 fanout8113 (.X(net8113),
    .A(net8118));
 sg13g2_buf_4 fanout8114 (.X(net8114),
    .A(net8116));
 sg13g2_buf_2 fanout8115 (.A(net8116),
    .X(net8115));
 sg13g2_buf_4 fanout8116 (.X(net8116),
    .A(net8118));
 sg13g2_buf_4 fanout8117 (.X(net8117),
    .A(net8118));
 sg13g2_buf_4 fanout8118 (.X(net8118),
    .A(_04617_));
 sg13g2_buf_4 fanout8119 (.X(net8119),
    .A(net8121));
 sg13g2_buf_4 fanout8120 (.X(net8120),
    .A(net8124));
 sg13g2_buf_2 fanout8121 (.A(net8124),
    .X(net8121));
 sg13g2_buf_8 fanout8122 (.A(net8124),
    .X(net8122));
 sg13g2_buf_4 fanout8123 (.X(net8123),
    .A(net8124));
 sg13g2_buf_4 fanout8124 (.X(net8124),
    .A(_04253_));
 sg13g2_buf_4 fanout8125 (.X(net8125),
    .A(net8127));
 sg13g2_buf_2 fanout8126 (.A(net8127),
    .X(net8126));
 sg13g2_buf_4 fanout8127 (.X(net8127),
    .A(net8129));
 sg13g2_buf_4 fanout8128 (.X(net8128),
    .A(net8129));
 sg13g2_buf_4 fanout8129 (.X(net8129),
    .A(_03776_));
 sg13g2_buf_4 fanout8130 (.X(net8130),
    .A(net8136));
 sg13g2_buf_4 fanout8131 (.X(net8131),
    .A(net8136));
 sg13g2_buf_4 fanout8132 (.X(net8132),
    .A(net8134));
 sg13g2_buf_2 fanout8133 (.A(net8134),
    .X(net8133));
 sg13g2_buf_4 fanout8134 (.X(net8134),
    .A(net8136));
 sg13g2_buf_4 fanout8135 (.X(net8135),
    .A(net8136));
 sg13g2_buf_8 fanout8136 (.A(_03776_),
    .X(net8136));
 sg13g2_buf_2 fanout8137 (.A(net8139),
    .X(net8137));
 sg13g2_buf_2 fanout8138 (.A(net8139),
    .X(net8138));
 sg13g2_buf_4 fanout8139 (.X(net8139),
    .A(net8140));
 sg13g2_buf_2 fanout8140 (.A(net8141),
    .X(net8140));
 sg13g2_buf_4 fanout8141 (.X(net8141),
    .A(_02849_));
 sg13g2_buf_4 fanout8142 (.X(net8142),
    .A(net8147));
 sg13g2_buf_4 fanout8143 (.X(net8143),
    .A(net8146));
 sg13g2_buf_4 fanout8144 (.X(net8144),
    .A(net8146));
 sg13g2_buf_4 fanout8145 (.X(net8145),
    .A(net8147));
 sg13g2_buf_2 fanout8146 (.A(net8147),
    .X(net8146));
 sg13g2_buf_4 fanout8147 (.X(net8147),
    .A(_02849_));
 sg13g2_buf_4 fanout8148 (.X(net8148),
    .A(net8150));
 sg13g2_buf_2 fanout8149 (.A(net8150),
    .X(net8149));
 sg13g2_buf_4 fanout8150 (.X(net8150),
    .A(net8151));
 sg13g2_buf_4 fanout8151 (.X(net8151),
    .A(net8159));
 sg13g2_buf_4 fanout8152 (.X(net8152),
    .A(net8159));
 sg13g2_buf_2 fanout8153 (.A(net8159),
    .X(net8153));
 sg13g2_buf_4 fanout8154 (.X(net8154),
    .A(net8158));
 sg13g2_buf_4 fanout8155 (.X(net8155),
    .A(net8157));
 sg13g2_buf_2 fanout8156 (.A(net8157),
    .X(net8156));
 sg13g2_buf_4 fanout8157 (.X(net8157),
    .A(net8158));
 sg13g2_buf_2 fanout8158 (.A(net8159),
    .X(net8158));
 sg13g2_buf_8 fanout8159 (.A(_02815_),
    .X(net8159));
 sg13g2_buf_4 fanout8160 (.X(net8160),
    .A(net8161));
 sg13g2_buf_4 fanout8161 (.X(net8161),
    .A(net8163));
 sg13g2_buf_4 fanout8162 (.X(net8162),
    .A(net8163));
 sg13g2_buf_8 fanout8163 (.A(_14404_),
    .X(net8163));
 sg13g2_buf_4 fanout8164 (.X(net8164),
    .A(net8170));
 sg13g2_buf_2 fanout8165 (.A(net8170),
    .X(net8165));
 sg13g2_buf_2 fanout8166 (.A(net8168),
    .X(net8166));
 sg13g2_buf_1 fanout8167 (.A(net8168),
    .X(net8167));
 sg13g2_buf_4 fanout8168 (.X(net8168),
    .A(net8170));
 sg13g2_buf_4 fanout8169 (.X(net8169),
    .A(net8170));
 sg13g2_buf_4 fanout8170 (.X(net8170),
    .A(_14404_));
 sg13g2_buf_4 fanout8171 (.X(net8171),
    .A(net8173));
 sg13g2_buf_2 fanout8172 (.A(net8173),
    .X(net8172));
 sg13g2_buf_4 fanout8173 (.X(net8173),
    .A(net8175));
 sg13g2_buf_4 fanout8174 (.X(net8174),
    .A(net8175));
 sg13g2_buf_2 fanout8175 (.A(net8183),
    .X(net8175));
 sg13g2_buf_4 fanout8176 (.X(net8176),
    .A(net8183));
 sg13g2_buf_2 fanout8177 (.A(net8183),
    .X(net8177));
 sg13g2_buf_4 fanout8178 (.X(net8178),
    .A(net8182));
 sg13g2_buf_4 fanout8179 (.X(net8179),
    .A(net8181));
 sg13g2_buf_1 fanout8180 (.A(net8181),
    .X(net8180));
 sg13g2_buf_2 fanout8181 (.A(net8182),
    .X(net8181));
 sg13g2_buf_4 fanout8182 (.X(net8182),
    .A(net8183));
 sg13g2_buf_4 fanout8183 (.X(net8183),
    .A(_14336_));
 sg13g2_buf_2 fanout8184 (.A(net8186),
    .X(net8184));
 sg13g2_buf_2 fanout8185 (.A(net8186),
    .X(net8185));
 sg13g2_buf_4 fanout8186 (.X(net8186),
    .A(net8188));
 sg13g2_buf_4 fanout8187 (.X(net8187),
    .A(net8188));
 sg13g2_buf_4 fanout8188 (.X(net8188),
    .A(net8196));
 sg13g2_buf_4 fanout8189 (.X(net8189),
    .A(net8196));
 sg13g2_buf_2 fanout8190 (.A(net8196),
    .X(net8190));
 sg13g2_buf_4 fanout8191 (.X(net8191),
    .A(net8195));
 sg13g2_buf_4 fanout8192 (.X(net8192),
    .A(net8194));
 sg13g2_buf_2 fanout8193 (.A(net8194),
    .X(net8193));
 sg13g2_buf_4 fanout8194 (.X(net8194),
    .A(net8195));
 sg13g2_buf_4 fanout8195 (.X(net8195),
    .A(net8196));
 sg13g2_buf_4 fanout8196 (.X(net8196),
    .A(_14303_));
 sg13g2_buf_4 fanout8197 (.X(net8197),
    .A(net8198));
 sg13g2_buf_4 fanout8198 (.X(net8198),
    .A(net8200));
 sg13g2_buf_4 fanout8199 (.X(net8199),
    .A(net8200));
 sg13g2_buf_8 fanout8200 (.A(net8208),
    .X(net8200));
 sg13g2_buf_4 fanout8201 (.X(net8201),
    .A(net8208));
 sg13g2_buf_2 fanout8202 (.A(net8208),
    .X(net8202));
 sg13g2_buf_4 fanout8203 (.X(net8203),
    .A(net8207));
 sg13g2_buf_4 fanout8204 (.X(net8204),
    .A(net8206));
 sg13g2_buf_2 fanout8205 (.A(net8206),
    .X(net8205));
 sg13g2_buf_2 fanout8206 (.A(net8207),
    .X(net8206));
 sg13g2_buf_4 fanout8207 (.X(net8207),
    .A(net8208));
 sg13g2_buf_4 fanout8208 (.X(net8208),
    .A(_14233_));
 sg13g2_buf_2 fanout8209 (.A(net8210),
    .X(net8209));
 sg13g2_buf_2 fanout8210 (.A(net8211),
    .X(net8210));
 sg13g2_buf_4 fanout8211 (.X(net8211),
    .A(net8213));
 sg13g2_buf_4 fanout8212 (.X(net8212),
    .A(net8213));
 sg13g2_buf_2 fanout8213 (.A(_14200_),
    .X(net8213));
 sg13g2_buf_4 fanout8214 (.X(net8214),
    .A(net8220));
 sg13g2_buf_4 fanout8215 (.X(net8215),
    .A(net8220));
 sg13g2_buf_4 fanout8216 (.X(net8216),
    .A(net8218));
 sg13g2_buf_2 fanout8217 (.A(net8218),
    .X(net8217));
 sg13g2_buf_4 fanout8218 (.X(net8218),
    .A(net8220));
 sg13g2_buf_4 fanout8219 (.X(net8219),
    .A(net8220));
 sg13g2_buf_4 fanout8220 (.X(net8220),
    .A(_14200_));
 sg13g2_buf_4 fanout8221 (.X(net8221),
    .A(net8223));
 sg13g2_buf_1 fanout8222 (.A(net8223),
    .X(net8222));
 sg13g2_buf_2 fanout8223 (.A(net8225),
    .X(net8223));
 sg13g2_buf_4 fanout8224 (.X(net8224),
    .A(net8225));
 sg13g2_buf_8 fanout8225 (.A(_14166_),
    .X(net8225));
 sg13g2_buf_4 fanout8226 (.X(net8226),
    .A(net8232));
 sg13g2_buf_4 fanout8227 (.X(net8227),
    .A(net8232));
 sg13g2_buf_4 fanout8228 (.X(net8228),
    .A(net8230));
 sg13g2_buf_2 fanout8229 (.A(net8230),
    .X(net8229));
 sg13g2_buf_4 fanout8230 (.X(net8230),
    .A(net8232));
 sg13g2_buf_4 fanout8231 (.X(net8231),
    .A(net8232));
 sg13g2_buf_4 fanout8232 (.X(net8232),
    .A(_14166_));
 sg13g2_buf_4 fanout8233 (.X(net8233),
    .A(net8234));
 sg13g2_buf_2 fanout8234 (.A(net8235),
    .X(net8234));
 sg13g2_buf_2 fanout8235 (.A(net8237),
    .X(net8235));
 sg13g2_buf_4 fanout8236 (.X(net8236),
    .A(net8237));
 sg13g2_buf_4 fanout8237 (.X(net8237),
    .A(_14131_));
 sg13g2_buf_8 fanout8238 (.A(net8244),
    .X(net8238));
 sg13g2_buf_2 fanout8239 (.A(net8244),
    .X(net8239));
 sg13g2_buf_4 fanout8240 (.X(net8240),
    .A(net8242));
 sg13g2_buf_2 fanout8241 (.A(net8242),
    .X(net8241));
 sg13g2_buf_4 fanout8242 (.X(net8242),
    .A(net8244));
 sg13g2_buf_4 fanout8243 (.X(net8243),
    .A(net8244));
 sg13g2_buf_4 fanout8244 (.X(net8244),
    .A(_14131_));
 sg13g2_buf_2 fanout8245 (.A(net8247),
    .X(net8245));
 sg13g2_buf_1 fanout8246 (.A(net8247),
    .X(net8246));
 sg13g2_buf_2 fanout8247 (.A(net8248),
    .X(net8247));
 sg13g2_buf_2 fanout8248 (.A(_11707_),
    .X(net8248));
 sg13g2_buf_4 fanout8249 (.X(net8249),
    .A(_11706_));
 sg13g2_buf_2 fanout8250 (.A(_11706_),
    .X(net8250));
 sg13g2_buf_4 fanout8251 (.X(net8251),
    .A(_11701_));
 sg13g2_buf_4 fanout8252 (.X(net8252),
    .A(net8254));
 sg13g2_buf_4 fanout8253 (.X(net8253),
    .A(net8254));
 sg13g2_buf_2 fanout8254 (.A(_11700_),
    .X(net8254));
 sg13g2_buf_2 fanout8255 (.A(net8256),
    .X(net8255));
 sg13g2_buf_2 fanout8256 (.A(net8257),
    .X(net8256));
 sg13g2_buf_4 fanout8257 (.X(net8257),
    .A(_11646_));
 sg13g2_buf_4 fanout8258 (.X(net8258),
    .A(_11645_));
 sg13g2_buf_4 fanout8259 (.X(net8259),
    .A(net8261));
 sg13g2_buf_2 fanout8260 (.A(net8261),
    .X(net8260));
 sg13g2_buf_4 fanout8261 (.X(net8261),
    .A(_11637_));
 sg13g2_buf_2 fanout8262 (.A(net8264),
    .X(net8262));
 sg13g2_buf_4 fanout8263 (.X(net8263),
    .A(net8264));
 sg13g2_buf_4 fanout8264 (.X(net8264),
    .A(_11636_));
 sg13g2_buf_4 fanout8265 (.X(net8265),
    .A(net8267));
 sg13g2_buf_2 fanout8266 (.A(net8267),
    .X(net8266));
 sg13g2_buf_4 fanout8267 (.X(net8267),
    .A(_11634_));
 sg13g2_buf_4 fanout8268 (.X(net8268),
    .A(net8269));
 sg13g2_buf_2 fanout8269 (.A(_11491_),
    .X(net8269));
 sg13g2_buf_4 fanout8270 (.X(net8270),
    .A(_11472_));
 sg13g2_buf_4 fanout8271 (.X(net8271),
    .A(net8272));
 sg13g2_buf_4 fanout8272 (.X(net8272),
    .A(_11462_));
 sg13g2_buf_4 fanout8273 (.X(net8273),
    .A(net8274));
 sg13g2_buf_4 fanout8274 (.X(net8274),
    .A(_11450_));
 sg13g2_buf_4 fanout8275 (.X(net8275),
    .A(_11439_));
 sg13g2_buf_4 fanout8276 (.X(net8276),
    .A(net8278));
 sg13g2_buf_2 fanout8277 (.A(net8278),
    .X(net8277));
 sg13g2_buf_4 fanout8278 (.X(net8278),
    .A(_11413_));
 sg13g2_buf_4 fanout8279 (.X(net8279),
    .A(net8280));
 sg13g2_buf_4 fanout8280 (.X(net8280),
    .A(_11401_));
 sg13g2_buf_4 fanout8281 (.X(net8281),
    .A(net8282));
 sg13g2_buf_8 fanout8282 (.A(_11391_),
    .X(net8282));
 sg13g2_buf_8 fanout8283 (.A(_11378_),
    .X(net8283));
 sg13g2_buf_4 fanout8284 (.X(net8284),
    .A(net8285));
 sg13g2_buf_4 fanout8285 (.X(net8285),
    .A(_11362_));
 sg13g2_buf_4 fanout8286 (.X(net8286),
    .A(_11349_));
 sg13g2_buf_4 fanout8287 (.X(net8287),
    .A(_11335_));
 sg13g2_buf_4 fanout8288 (.X(net8288),
    .A(net8289));
 sg13g2_buf_4 fanout8289 (.X(net8289),
    .A(_11322_));
 sg13g2_buf_4 fanout8290 (.X(net8290),
    .A(_11307_));
 sg13g2_buf_8 fanout8291 (.A(_11303_),
    .X(net8291));
 sg13g2_buf_4 fanout8292 (.X(net8292),
    .A(_11291_));
 sg13g2_buf_4 fanout8293 (.X(net8293),
    .A(_11280_));
 sg13g2_buf_2 fanout8294 (.A(_11280_),
    .X(net8294));
 sg13g2_buf_8 fanout8295 (.A(_11267_),
    .X(net8295));
 sg13g2_buf_4 fanout8296 (.X(net8296),
    .A(_11234_));
 sg13g2_buf_2 fanout8297 (.A(_11234_),
    .X(net8297));
 sg13g2_buf_4 fanout8298 (.X(net8298),
    .A(_11185_));
 sg13g2_buf_4 fanout8299 (.X(net8299),
    .A(net8300));
 sg13g2_buf_4 fanout8300 (.X(net8300),
    .A(_11159_));
 sg13g2_buf_4 fanout8301 (.X(net8301),
    .A(net8302));
 sg13g2_buf_4 fanout8302 (.X(net8302),
    .A(_11132_));
 sg13g2_buf_4 fanout8303 (.X(net8303),
    .A(_11117_));
 sg13g2_buf_4 fanout8304 (.X(net8304),
    .A(net8306));
 sg13g2_buf_2 fanout8305 (.A(net8306),
    .X(net8305));
 sg13g2_buf_4 fanout8306 (.X(net8306),
    .A(_11106_));
 sg13g2_buf_4 fanout8307 (.X(net8307),
    .A(net8308));
 sg13g2_buf_4 fanout8308 (.X(net8308),
    .A(_11078_));
 sg13g2_buf_4 fanout8309 (.X(net8309),
    .A(_11068_));
 sg13g2_buf_4 fanout8310 (.X(net8310),
    .A(net8312));
 sg13g2_buf_4 fanout8311 (.X(net8311),
    .A(net8312));
 sg13g2_buf_8 fanout8312 (.A(_11043_),
    .X(net8312));
 sg13g2_buf_4 fanout8313 (.X(net8313),
    .A(_11042_));
 sg13g2_buf_4 fanout8314 (.X(net8314),
    .A(_10992_));
 sg13g2_buf_4 fanout8315 (.X(net8315),
    .A(_10992_));
 sg13g2_buf_2 fanout8316 (.A(_09056_),
    .X(net8316));
 sg13g2_buf_2 fanout8317 (.A(_09056_),
    .X(net8317));
 sg13g2_buf_2 fanout8318 (.A(net8319),
    .X(net8318));
 sg13g2_buf_2 fanout8319 (.A(net8322),
    .X(net8319));
 sg13g2_buf_2 fanout8320 (.A(net8321),
    .X(net8320));
 sg13g2_buf_2 fanout8321 (.A(net8322),
    .X(net8321));
 sg13g2_buf_2 fanout8322 (.A(_08962_),
    .X(net8322));
 sg13g2_buf_2 fanout8323 (.A(net8327),
    .X(net8323));
 sg13g2_buf_2 fanout8324 (.A(net8327),
    .X(net8324));
 sg13g2_buf_2 fanout8325 (.A(net8327),
    .X(net8325));
 sg13g2_buf_1 fanout8326 (.A(net8327),
    .X(net8326));
 sg13g2_buf_1 fanout8327 (.A(_07212_),
    .X(net8327));
 sg13g2_buf_2 fanout8328 (.A(_07211_),
    .X(net8328));
 sg13g2_buf_2 fanout8329 (.A(_07211_),
    .X(net8329));
 sg13g2_buf_2 fanout8330 (.A(net8332),
    .X(net8330));
 sg13g2_buf_1 fanout8331 (.A(net8332),
    .X(net8331));
 sg13g2_buf_1 fanout8332 (.A(net8333),
    .X(net8332));
 sg13g2_buf_2 fanout8333 (.A(_07211_),
    .X(net8333));
 sg13g2_buf_4 fanout8334 (.X(net8334),
    .A(net8336));
 sg13g2_buf_4 fanout8335 (.X(net8335),
    .A(net8336));
 sg13g2_buf_4 fanout8336 (.X(net8336),
    .A(_03839_));
 sg13g2_buf_4 fanout8337 (.X(net8337),
    .A(_03839_));
 sg13g2_buf_1 fanout8338 (.A(_03839_),
    .X(net8338));
 sg13g2_buf_4 fanout8339 (.X(net8339),
    .A(net8340));
 sg13g2_buf_4 fanout8340 (.X(net8340),
    .A(_03835_));
 sg13g2_buf_4 fanout8341 (.X(net8341),
    .A(net8342));
 sg13g2_buf_8 fanout8342 (.A(_03835_),
    .X(net8342));
 sg13g2_buf_4 fanout8343 (.X(net8343),
    .A(net8344));
 sg13g2_buf_8 fanout8344 (.A(_03834_),
    .X(net8344));
 sg13g2_buf_4 fanout8345 (.X(net8345),
    .A(net8348));
 sg13g2_buf_4 fanout8346 (.X(net8346),
    .A(net8348));
 sg13g2_buf_8 fanout8347 (.A(net8348),
    .X(net8347));
 sg13g2_buf_8 fanout8348 (.A(_03831_),
    .X(net8348));
 sg13g2_buf_4 fanout8349 (.X(net8349),
    .A(net8353));
 sg13g2_buf_4 fanout8350 (.X(net8350),
    .A(net8353));
 sg13g2_buf_2 fanout8351 (.A(net8352),
    .X(net8351));
 sg13g2_buf_4 fanout8352 (.X(net8352),
    .A(net8353));
 sg13g2_buf_2 fanout8353 (.A(net8360),
    .X(net8353));
 sg13g2_buf_4 fanout8354 (.X(net8354),
    .A(net8355));
 sg13g2_buf_2 fanout8355 (.A(net8356),
    .X(net8355));
 sg13g2_buf_4 fanout8356 (.X(net8356),
    .A(net8360));
 sg13g2_buf_2 fanout8357 (.A(net8359),
    .X(net8357));
 sg13g2_buf_2 fanout8358 (.A(net8359),
    .X(net8358));
 sg13g2_buf_2 fanout8359 (.A(net8360),
    .X(net8359));
 sg13g2_buf_2 fanout8360 (.A(_03823_),
    .X(net8360));
 sg13g2_buf_4 fanout8361 (.X(net8361),
    .A(net8366));
 sg13g2_buf_2 fanout8362 (.A(net8366),
    .X(net8362));
 sg13g2_buf_4 fanout8363 (.X(net8363),
    .A(net8365));
 sg13g2_buf_2 fanout8364 (.A(net8365),
    .X(net8364));
 sg13g2_buf_4 fanout8365 (.X(net8365),
    .A(net8366));
 sg13g2_buf_2 fanout8366 (.A(net8370),
    .X(net8366));
 sg13g2_buf_2 fanout8367 (.A(net8368),
    .X(net8367));
 sg13g2_buf_2 fanout8368 (.A(net8369),
    .X(net8368));
 sg13g2_buf_2 fanout8369 (.A(net8370),
    .X(net8369));
 sg13g2_buf_4 fanout8370 (.X(net8370),
    .A(_03822_));
 sg13g2_buf_2 fanout8371 (.A(net8372),
    .X(net8371));
 sg13g2_buf_2 fanout8372 (.A(_14129_),
    .X(net8372));
 sg13g2_buf_2 fanout8373 (.A(_13299_),
    .X(net8373));
 sg13g2_buf_4 fanout8374 (.X(net8374),
    .A(net8375));
 sg13g2_buf_2 fanout8375 (.A(_11760_),
    .X(net8375));
 sg13g2_buf_2 fanout8376 (.A(net8378),
    .X(net8376));
 sg13g2_buf_4 fanout8377 (.X(net8377),
    .A(net8378));
 sg13g2_buf_4 fanout8378 (.X(net8378),
    .A(_11760_));
 sg13g2_buf_4 fanout8379 (.X(net8379),
    .A(_11394_));
 sg13g2_buf_4 fanout8380 (.X(net8380),
    .A(_11294_));
 sg13g2_buf_4 fanout8381 (.X(net8381),
    .A(_11282_));
 sg13g2_buf_4 fanout8382 (.X(net8382),
    .A(_11238_));
 sg13g2_buf_2 fanout8383 (.A(net8388),
    .X(net8383));
 sg13g2_buf_2 fanout8384 (.A(net8385),
    .X(net8384));
 sg13g2_buf_1 fanout8385 (.A(net8388),
    .X(net8385));
 sg13g2_buf_2 fanout8386 (.A(net8387),
    .X(net8386));
 sg13g2_buf_2 fanout8387 (.A(net8388),
    .X(net8387));
 sg13g2_buf_4 fanout8388 (.X(net8388),
    .A(_11182_));
 sg13g2_buf_2 fanout8389 (.A(net8390),
    .X(net8389));
 sg13g2_buf_2 fanout8390 (.A(net8399),
    .X(net8390));
 sg13g2_buf_2 fanout8391 (.A(net8399),
    .X(net8391));
 sg13g2_buf_2 fanout8392 (.A(net8399),
    .X(net8392));
 sg13g2_buf_2 fanout8393 (.A(net8398),
    .X(net8393));
 sg13g2_buf_2 fanout8394 (.A(net8398),
    .X(net8394));
 sg13g2_buf_2 fanout8395 (.A(net8396),
    .X(net8395));
 sg13g2_buf_2 fanout8396 (.A(net8398),
    .X(net8396));
 sg13g2_buf_2 fanout8397 (.A(net8398),
    .X(net8397));
 sg13g2_buf_2 fanout8398 (.A(net8399),
    .X(net8398));
 sg13g2_buf_2 fanout8399 (.A(_11169_),
    .X(net8399));
 sg13g2_buf_4 fanout8400 (.X(net8400),
    .A(net8408));
 sg13g2_buf_2 fanout8401 (.A(net8402),
    .X(net8401));
 sg13g2_buf_2 fanout8402 (.A(net8403),
    .X(net8402));
 sg13g2_buf_2 fanout8403 (.A(net8408),
    .X(net8403));
 sg13g2_buf_2 fanout8404 (.A(net8407),
    .X(net8404));
 sg13g2_buf_1 fanout8405 (.A(net8407),
    .X(net8405));
 sg13g2_buf_2 fanout8406 (.A(net8407),
    .X(net8406));
 sg13g2_buf_2 fanout8407 (.A(net8408),
    .X(net8407));
 sg13g2_buf_4 fanout8408 (.X(net8408),
    .A(_11168_));
 sg13g2_buf_2 fanout8409 (.A(net8410),
    .X(net8409));
 sg13g2_buf_2 fanout8410 (.A(net8412),
    .X(net8410));
 sg13g2_buf_2 fanout8411 (.A(net8412),
    .X(net8411));
 sg13g2_buf_1 fanout8412 (.A(net8413),
    .X(net8412));
 sg13g2_buf_2 fanout8413 (.A(net8414),
    .X(net8413));
 sg13g2_buf_2 fanout8414 (.A(net8426),
    .X(net8414));
 sg13g2_buf_2 fanout8415 (.A(net8416),
    .X(net8415));
 sg13g2_buf_2 fanout8416 (.A(net8426),
    .X(net8416));
 sg13g2_buf_2 fanout8417 (.A(net8418),
    .X(net8417));
 sg13g2_buf_2 fanout8418 (.A(net8419),
    .X(net8418));
 sg13g2_buf_2 fanout8419 (.A(net8426),
    .X(net8419));
 sg13g2_buf_2 fanout8420 (.A(net8421),
    .X(net8420));
 sg13g2_buf_2 fanout8421 (.A(net8425),
    .X(net8421));
 sg13g2_buf_2 fanout8422 (.A(net8424),
    .X(net8422));
 sg13g2_buf_1 fanout8423 (.A(net8424),
    .X(net8423));
 sg13g2_buf_2 fanout8424 (.A(net8425),
    .X(net8424));
 sg13g2_buf_2 fanout8425 (.A(net8426),
    .X(net8425));
 sg13g2_buf_2 fanout8426 (.A(_11153_),
    .X(net8426));
 sg13g2_buf_4 fanout8427 (.X(net8427),
    .A(net8429));
 sg13g2_buf_2 fanout8428 (.A(net8429),
    .X(net8428));
 sg13g2_buf_4 fanout8429 (.X(net8429),
    .A(net8430));
 sg13g2_buf_4 fanout8430 (.X(net8430),
    .A(_11152_));
 sg13g2_buf_2 fanout8431 (.A(net8436),
    .X(net8431));
 sg13g2_buf_4 fanout8432 (.X(net8432),
    .A(net8433));
 sg13g2_buf_2 fanout8433 (.A(net8435),
    .X(net8433));
 sg13g2_buf_2 fanout8434 (.A(net8435),
    .X(net8434));
 sg13g2_buf_2 fanout8435 (.A(net8436),
    .X(net8435));
 sg13g2_buf_1 fanout8436 (.A(net8437),
    .X(net8436));
 sg13g2_buf_4 fanout8437 (.X(net8437),
    .A(_11137_));
 sg13g2_buf_4 fanout8438 (.X(net8438),
    .A(net8440));
 sg13g2_buf_4 fanout8439 (.X(net8439),
    .A(net8440));
 sg13g2_buf_2 fanout8440 (.A(net8441),
    .X(net8440));
 sg13g2_buf_4 fanout8441 (.X(net8441),
    .A(_11136_));
 sg13g2_buf_2 fanout8442 (.A(net8444),
    .X(net8442));
 sg13g2_buf_1 fanout8443 (.A(net8444),
    .X(net8443));
 sg13g2_buf_2 fanout8444 (.A(net8445),
    .X(net8444));
 sg13g2_buf_2 fanout8445 (.A(net8446),
    .X(net8445));
 sg13g2_buf_4 fanout8446 (.X(net8446),
    .A(_11125_));
 sg13g2_buf_2 fanout8447 (.A(net8449),
    .X(net8447));
 sg13g2_buf_2 fanout8448 (.A(net8449),
    .X(net8448));
 sg13g2_buf_2 fanout8449 (.A(net8450),
    .X(net8449));
 sg13g2_buf_4 fanout8450 (.X(net8450),
    .A(net8451));
 sg13g2_buf_4 fanout8451 (.X(net8451),
    .A(_11124_));
 sg13g2_buf_2 fanout8452 (.A(net8453),
    .X(net8452));
 sg13g2_buf_2 fanout8453 (.A(_07302_),
    .X(net8453));
 sg13g2_buf_4 fanout8454 (.X(net8454),
    .A(net8456));
 sg13g2_buf_2 fanout8455 (.A(net8456),
    .X(net8455));
 sg13g2_buf_4 fanout8456 (.X(net8456),
    .A(net8457));
 sg13g2_buf_4 fanout8457 (.X(net8457),
    .A(_05648_));
 sg13g2_buf_2 fanout8458 (.A(net8459),
    .X(net8458));
 sg13g2_buf_4 fanout8459 (.X(net8459),
    .A(net8461));
 sg13g2_buf_4 fanout8460 (.X(net8460),
    .A(net8461));
 sg13g2_buf_2 fanout8461 (.A(net8465),
    .X(net8461));
 sg13g2_buf_4 fanout8462 (.X(net8462),
    .A(net8464));
 sg13g2_buf_4 fanout8463 (.X(net8463),
    .A(net8464));
 sg13g2_buf_2 fanout8464 (.A(net8465),
    .X(net8464));
 sg13g2_buf_2 fanout8465 (.A(_05648_),
    .X(net8465));
 sg13g2_buf_2 fanout8466 (.A(net8467),
    .X(net8466));
 sg13g2_buf_1 fanout8467 (.A(net8468),
    .X(net8467));
 sg13g2_buf_1 fanout8468 (.A(net8469),
    .X(net8468));
 sg13g2_buf_2 fanout8469 (.A(net8471),
    .X(net8469));
 sg13g2_buf_4 fanout8470 (.X(net8470),
    .A(net8471));
 sg13g2_buf_2 fanout8471 (.A(_05647_),
    .X(net8471));
 sg13g2_buf_2 fanout8472 (.A(net8474),
    .X(net8472));
 sg13g2_buf_2 fanout8473 (.A(net8474),
    .X(net8473));
 sg13g2_buf_1 fanout8474 (.A(net8475),
    .X(net8474));
 sg13g2_buf_2 fanout8475 (.A(_05647_),
    .X(net8475));
 sg13g2_buf_2 fanout8476 (.A(net8477),
    .X(net8476));
 sg13g2_buf_2 fanout8477 (.A(net8481),
    .X(net8477));
 sg13g2_buf_2 fanout8478 (.A(net8479),
    .X(net8478));
 sg13g2_buf_2 fanout8479 (.A(net8481),
    .X(net8479));
 sg13g2_buf_2 fanout8480 (.A(net8481),
    .X(net8480));
 sg13g2_buf_2 fanout8481 (.A(net8482),
    .X(net8481));
 sg13g2_buf_4 fanout8482 (.X(net8482),
    .A(_04837_));
 sg13g2_buf_4 fanout8483 (.X(net8483),
    .A(net8484));
 sg13g2_buf_2 fanout8484 (.A(net8485),
    .X(net8484));
 sg13g2_buf_2 fanout8485 (.A(_04836_),
    .X(net8485));
 sg13g2_buf_4 fanout8486 (.X(net8486),
    .A(net8487));
 sg13g2_buf_4 fanout8487 (.X(net8487),
    .A(net8492));
 sg13g2_buf_2 fanout8488 (.A(net8489),
    .X(net8488));
 sg13g2_buf_2 fanout8489 (.A(net8491),
    .X(net8489));
 sg13g2_buf_2 fanout8490 (.A(net8491),
    .X(net8490));
 sg13g2_buf_2 fanout8491 (.A(net8492),
    .X(net8491));
 sg13g2_buf_4 fanout8492 (.X(net8492),
    .A(_03817_));
 sg13g2_buf_2 fanout8493 (.A(net8494),
    .X(net8493));
 sg13g2_buf_2 fanout8494 (.A(net8496),
    .X(net8494));
 sg13g2_buf_4 fanout8495 (.X(net8495),
    .A(net8496));
 sg13g2_buf_2 fanout8496 (.A(_13297_),
    .X(net8496));
 sg13g2_buf_2 fanout8497 (.A(_13296_),
    .X(net8497));
 sg13g2_buf_2 fanout8498 (.A(_13296_),
    .X(net8498));
 sg13g2_buf_2 fanout8499 (.A(net8500),
    .X(net8499));
 sg13g2_buf_2 fanout8500 (.A(_11746_),
    .X(net8500));
 sg13g2_buf_2 fanout8501 (.A(net8502),
    .X(net8501));
 sg13g2_buf_4 fanout8502 (.X(net8502),
    .A(_11746_));
 sg13g2_buf_2 fanout8503 (.A(net8504),
    .X(net8503));
 sg13g2_buf_2 fanout8504 (.A(_11746_),
    .X(net8504));
 sg13g2_buf_4 fanout8505 (.X(net8505),
    .A(_11250_));
 sg13g2_buf_4 fanout8506 (.X(net8506),
    .A(_11225_));
 sg13g2_buf_4 fanout8507 (.X(net8507),
    .A(_11212_));
 sg13g2_buf_2 fanout8508 (.A(net8509),
    .X(net8508));
 sg13g2_buf_1 fanout8509 (.A(net8510),
    .X(net8509));
 sg13g2_buf_2 fanout8510 (.A(net8518),
    .X(net8510));
 sg13g2_buf_2 fanout8511 (.A(net8512),
    .X(net8511));
 sg13g2_buf_1 fanout8512 (.A(net8513),
    .X(net8512));
 sg13g2_buf_2 fanout8513 (.A(net8518),
    .X(net8513));
 sg13g2_buf_2 fanout8514 (.A(net8518),
    .X(net8514));
 sg13g2_buf_2 fanout8515 (.A(net8516),
    .X(net8515));
 sg13g2_buf_2 fanout8516 (.A(net8517),
    .X(net8516));
 sg13g2_buf_1 fanout8517 (.A(net8518),
    .X(net8517));
 sg13g2_buf_2 fanout8518 (.A(net8519),
    .X(net8518));
 sg13g2_buf_2 fanout8519 (.A(_11181_),
    .X(net8519));
 sg13g2_buf_4 fanout8520 (.X(net8520),
    .A(_11109_));
 sg13g2_buf_4 fanout8521 (.X(net8521),
    .A(_11100_));
 sg13g2_buf_4 fanout8522 (.X(net8522),
    .A(_11090_));
 sg13g2_buf_2 fanout8523 (.A(_11060_),
    .X(net8523));
 sg13g2_buf_4 fanout8524 (.X(net8524),
    .A(net8525));
 sg13g2_buf_8 fanout8525 (.A(_10989_),
    .X(net8525));
 sg13g2_buf_2 fanout8526 (.A(net8528),
    .X(net8526));
 sg13g2_buf_4 fanout8527 (.X(net8527),
    .A(net8528));
 sg13g2_buf_4 fanout8528 (.X(net8528),
    .A(_10989_));
 sg13g2_buf_4 fanout8529 (.X(net8529),
    .A(_10965_));
 sg13g2_buf_4 fanout8530 (.X(net8530),
    .A(_08722_));
 sg13g2_buf_2 fanout8531 (.A(net8536),
    .X(net8531));
 sg13g2_buf_2 fanout8532 (.A(net8533),
    .X(net8532));
 sg13g2_buf_2 fanout8533 (.A(net8535),
    .X(net8533));
 sg13g2_buf_1 fanout8534 (.A(net8535),
    .X(net8534));
 sg13g2_buf_1 fanout8535 (.A(net8536),
    .X(net8535));
 sg13g2_buf_2 fanout8536 (.A(_07511_),
    .X(net8536));
 sg13g2_buf_4 fanout8537 (.X(net8537),
    .A(_07432_));
 sg13g2_buf_2 fanout8538 (.A(net8540),
    .X(net8538));
 sg13g2_buf_1 fanout8539 (.A(net8540),
    .X(net8539));
 sg13g2_buf_2 fanout8540 (.A(_06857_),
    .X(net8540));
 sg13g2_buf_2 fanout8541 (.A(net8542),
    .X(net8541));
 sg13g2_buf_2 fanout8542 (.A(_06856_),
    .X(net8542));
 sg13g2_buf_4 fanout8543 (.X(net8543),
    .A(_04611_));
 sg13g2_buf_4 fanout8544 (.X(net8544),
    .A(_02813_));
 sg13g2_buf_4 fanout8545 (.X(net8545),
    .A(_02808_));
 sg13g2_buf_4 fanout8546 (.X(net8546),
    .A(_02803_));
 sg13g2_buf_4 fanout8547 (.X(net8547),
    .A(_02799_));
 sg13g2_buf_4 fanout8548 (.X(net8548),
    .A(_14124_));
 sg13g2_buf_8 fanout8549 (.A(net8550),
    .X(net8549));
 sg13g2_buf_4 fanout8550 (.X(net8550),
    .A(_13998_));
 sg13g2_buf_2 fanout8551 (.A(_12562_),
    .X(net8551));
 sg13g2_buf_2 fanout8552 (.A(_12562_),
    .X(net8552));
 sg13g2_buf_2 fanout8553 (.A(net8554),
    .X(net8553));
 sg13g2_buf_2 fanout8554 (.A(net8555),
    .X(net8554));
 sg13g2_buf_2 fanout8555 (.A(_12562_),
    .X(net8555));
 sg13g2_buf_2 fanout8556 (.A(net8557),
    .X(net8556));
 sg13g2_buf_1 fanout8557 (.A(net8558),
    .X(net8557));
 sg13g2_buf_2 fanout8558 (.A(_12561_),
    .X(net8558));
 sg13g2_buf_2 fanout8559 (.A(net8561),
    .X(net8559));
 sg13g2_buf_2 fanout8560 (.A(net8561),
    .X(net8560));
 sg13g2_buf_2 fanout8561 (.A(_12561_),
    .X(net8561));
 sg13g2_buf_4 fanout8562 (.X(net8562),
    .A(_11175_));
 sg13g2_buf_2 fanout8563 (.A(_11175_),
    .X(net8563));
 sg13g2_buf_2 fanout8564 (.A(net8565),
    .X(net8564));
 sg13g2_buf_2 fanout8565 (.A(net8569),
    .X(net8565));
 sg13g2_buf_2 fanout8566 (.A(net8567),
    .X(net8566));
 sg13g2_buf_2 fanout8567 (.A(net8568),
    .X(net8567));
 sg13g2_buf_2 fanout8568 (.A(net8569),
    .X(net8568));
 sg13g2_buf_2 fanout8569 (.A(_10978_),
    .X(net8569));
 sg13g2_buf_2 fanout8570 (.A(net8571),
    .X(net8570));
 sg13g2_buf_2 fanout8571 (.A(net8572),
    .X(net8571));
 sg13g2_buf_4 fanout8572 (.X(net8572),
    .A(net8573));
 sg13g2_buf_2 fanout8573 (.A(net8574),
    .X(net8573));
 sg13g2_buf_4 fanout8574 (.X(net8574),
    .A(_10859_));
 sg13g2_buf_8 fanout8575 (.A(net8578),
    .X(net8575));
 sg13g2_buf_4 fanout8576 (.X(net8576),
    .A(net8578));
 sg13g2_buf_4 fanout8577 (.X(net8577),
    .A(net8578));
 sg13g2_buf_4 fanout8578 (.X(net8578),
    .A(_10859_));
 sg13g2_buf_4 fanout8579 (.X(net8579),
    .A(_08724_));
 sg13g2_buf_2 fanout8580 (.A(net8581),
    .X(net8580));
 sg13g2_buf_1 fanout8581 (.A(_07510_),
    .X(net8581));
 sg13g2_buf_2 fanout8582 (.A(_07186_),
    .X(net8582));
 sg13g2_buf_4 fanout8583 (.X(net8583),
    .A(_07001_));
 sg13g2_buf_4 fanout8584 (.X(net8584),
    .A(_06952_));
 sg13g2_buf_4 fanout8585 (.X(net8585),
    .A(net8590));
 sg13g2_buf_2 fanout8586 (.A(net8590),
    .X(net8586));
 sg13g2_buf_4 fanout8587 (.X(net8587),
    .A(net8588));
 sg13g2_buf_4 fanout8588 (.X(net8588),
    .A(net8589));
 sg13g2_buf_2 fanout8589 (.A(net8590),
    .X(net8589));
 sg13g2_buf_4 fanout8590 (.X(net8590),
    .A(_05756_));
 sg13g2_buf_4 fanout8591 (.X(net8591),
    .A(_04615_));
 sg13g2_buf_4 fanout8592 (.X(net8592),
    .A(_04613_));
 sg13g2_buf_4 fanout8593 (.X(net8593),
    .A(_04609_));
 sg13g2_buf_8 fanout8594 (.A(net8596),
    .X(net8594));
 sg13g2_buf_8 fanout8595 (.A(net8596),
    .X(net8595));
 sg13g2_buf_8 fanout8596 (.A(_02905_),
    .X(net8596));
 sg13g2_buf_16 fanout8597 (.X(net8597),
    .A(_02904_));
 sg13g2_buf_4 fanout8598 (.X(net8598),
    .A(_02904_));
 sg13g2_buf_4 fanout8599 (.X(net8599),
    .A(_02811_));
 sg13g2_buf_4 fanout8600 (.X(net8600),
    .A(_02806_));
 sg13g2_buf_2 fanout8601 (.A(net8602),
    .X(net8601));
 sg13g2_buf_1 fanout8602 (.A(net8603),
    .X(net8602));
 sg13g2_buf_2 fanout8603 (.A(_14273_),
    .X(net8603));
 sg13g2_buf_8 fanout8604 (.A(_14017_),
    .X(net8604));
 sg13g2_buf_2 fanout8605 (.A(_14017_),
    .X(net8605));
 sg13g2_buf_8 fanout8606 (.A(_14011_),
    .X(net8606));
 sg13g2_buf_2 fanout8607 (.A(_14011_),
    .X(net8607));
 sg13g2_buf_8 fanout8608 (.A(net8609),
    .X(net8608));
 sg13g2_buf_8 fanout8609 (.A(_14004_),
    .X(net8609));
 sg13g2_buf_8 fanout8610 (.A(_13992_),
    .X(net8610));
 sg13g2_buf_4 fanout8611 (.X(net8611),
    .A(_13992_));
 sg13g2_buf_8 fanout8612 (.A(_13986_),
    .X(net8612));
 sg13g2_buf_4 fanout8613 (.X(net8613),
    .A(_13986_));
 sg13g2_buf_4 fanout8614 (.X(net8614),
    .A(net8615));
 sg13g2_buf_4 fanout8615 (.X(net8615),
    .A(net8625));
 sg13g2_buf_2 fanout8616 (.A(net8625),
    .X(net8616));
 sg13g2_buf_4 fanout8617 (.X(net8617),
    .A(net8619));
 sg13g2_buf_2 fanout8618 (.A(net8619),
    .X(net8618));
 sg13g2_buf_2 fanout8619 (.A(net8624),
    .X(net8619));
 sg13g2_buf_2 fanout8620 (.A(net8621),
    .X(net8620));
 sg13g2_buf_2 fanout8621 (.A(net8622),
    .X(net8621));
 sg13g2_buf_2 fanout8622 (.A(net8623),
    .X(net8622));
 sg13g2_buf_2 fanout8623 (.A(net8624),
    .X(net8623));
 sg13g2_buf_2 fanout8624 (.A(net8625),
    .X(net8624));
 sg13g2_buf_4 fanout8625 (.X(net8625),
    .A(_13833_));
 sg13g2_buf_4 fanout8626 (.X(net8626),
    .A(_12560_));
 sg13g2_buf_2 fanout8627 (.A(net8629),
    .X(net8627));
 sg13g2_buf_2 fanout8628 (.A(net8629),
    .X(net8628));
 sg13g2_buf_2 fanout8629 (.A(_11733_),
    .X(net8629));
 sg13g2_buf_2 fanout8630 (.A(net8631),
    .X(net8630));
 sg13g2_buf_2 fanout8631 (.A(net8634),
    .X(net8631));
 sg13g2_buf_4 fanout8632 (.X(net8632),
    .A(net8633));
 sg13g2_buf_2 fanout8633 (.A(net8634),
    .X(net8633));
 sg13g2_buf_4 fanout8634 (.X(net8634),
    .A(_11733_));
 sg13g2_buf_2 fanout8635 (.A(net8636),
    .X(net8635));
 sg13g2_buf_2 fanout8636 (.A(net8637),
    .X(net8636));
 sg13g2_buf_4 fanout8637 (.X(net8637),
    .A(_11019_));
 sg13g2_buf_4 fanout8638 (.X(net8638),
    .A(net8639));
 sg13g2_buf_4 fanout8639 (.X(net8639),
    .A(net8640));
 sg13g2_buf_2 fanout8640 (.A(_11018_),
    .X(net8640));
 sg13g2_buf_2 fanout8641 (.A(_11013_),
    .X(net8641));
 sg13g2_buf_2 fanout8642 (.A(net8643),
    .X(net8642));
 sg13g2_buf_4 fanout8643 (.X(net8643),
    .A(_10996_));
 sg13g2_buf_2 fanout8644 (.A(net8645),
    .X(net8644));
 sg13g2_buf_1 fanout8645 (.A(net8646),
    .X(net8645));
 sg13g2_buf_2 fanout8646 (.A(_10995_),
    .X(net8646));
 sg13g2_buf_2 fanout8647 (.A(net8649),
    .X(net8647));
 sg13g2_buf_2 fanout8648 (.A(_10995_),
    .X(net8648));
 sg13g2_buf_2 fanout8649 (.A(_10995_),
    .X(net8649));
 sg13g2_buf_2 fanout8650 (.A(net8651),
    .X(net8650));
 sg13g2_buf_2 fanout8651 (.A(_10986_),
    .X(net8651));
 sg13g2_buf_2 fanout8652 (.A(net8653),
    .X(net8652));
 sg13g2_buf_2 fanout8653 (.A(net8654),
    .X(net8653));
 sg13g2_buf_2 fanout8654 (.A(_10986_),
    .X(net8654));
 sg13g2_buf_8 fanout8655 (.A(_10869_),
    .X(net8655));
 sg13g2_buf_4 fanout8656 (.X(net8656),
    .A(net8664));
 sg13g2_buf_2 fanout8657 (.A(net8663),
    .X(net8657));
 sg13g2_buf_1 fanout8658 (.A(net8663),
    .X(net8658));
 sg13g2_buf_4 fanout8659 (.X(net8659),
    .A(net8663));
 sg13g2_buf_2 fanout8660 (.A(net8661),
    .X(net8660));
 sg13g2_buf_2 fanout8661 (.A(net8663),
    .X(net8661));
 sg13g2_buf_2 fanout8662 (.A(net8663),
    .X(net8662));
 sg13g2_buf_4 fanout8663 (.X(net8663),
    .A(net8664));
 sg13g2_buf_2 fanout8664 (.A(_10868_),
    .X(net8664));
 sg13g2_buf_4 fanout8665 (.X(net8665),
    .A(net8666));
 sg13g2_buf_4 fanout8666 (.X(net8666),
    .A(net8667));
 sg13g2_buf_4 fanout8667 (.X(net8667),
    .A(_10857_));
 sg13g2_buf_2 fanout8668 (.A(net8670),
    .X(net8668));
 sg13g2_buf_1 fanout8669 (.A(net8670),
    .X(net8669));
 sg13g2_buf_2 fanout8670 (.A(_07176_),
    .X(net8670));
 sg13g2_buf_2 fanout8671 (.A(_06859_),
    .X(net8671));
 sg13g2_buf_2 fanout8672 (.A(_06859_),
    .X(net8672));
 sg13g2_buf_4 fanout8673 (.X(net8673),
    .A(_03818_));
 sg13g2_buf_8 fanout8674 (.A(_02895_),
    .X(net8674));
 sg13g2_buf_4 fanout8675 (.X(net8675),
    .A(_13238_));
 sg13g2_buf_1 fanout8676 (.A(_13238_),
    .X(net8676));
 sg13g2_buf_2 fanout8677 (.A(net8678),
    .X(net8677));
 sg13g2_buf_2 fanout8678 (.A(net8679),
    .X(net8678));
 sg13g2_buf_2 fanout8679 (.A(_11851_),
    .X(net8679));
 sg13g2_buf_2 fanout8680 (.A(net8682),
    .X(net8680));
 sg13g2_buf_4 fanout8681 (.X(net8681),
    .A(net8682));
 sg13g2_buf_4 fanout8682 (.X(net8682),
    .A(_11851_));
 sg13g2_buf_2 fanout8683 (.A(net8685),
    .X(net8683));
 sg13g2_buf_1 fanout8684 (.A(net8685),
    .X(net8684));
 sg13g2_buf_2 fanout8685 (.A(net8686),
    .X(net8685));
 sg13g2_buf_2 fanout8686 (.A(_11850_),
    .X(net8686));
 sg13g2_buf_2 fanout8687 (.A(net8688),
    .X(net8687));
 sg13g2_buf_1 fanout8688 (.A(net8689),
    .X(net8688));
 sg13g2_buf_2 fanout8689 (.A(_11850_),
    .X(net8689));
 sg13g2_buf_4 fanout8690 (.X(net8690),
    .A(_11740_));
 sg13g2_buf_2 fanout8691 (.A(net8695),
    .X(net8691));
 sg13g2_buf_2 fanout8692 (.A(net8693),
    .X(net8692));
 sg13g2_buf_1 fanout8693 (.A(net8694),
    .X(net8693));
 sg13g2_buf_2 fanout8694 (.A(net8695),
    .X(net8694));
 sg13g2_buf_4 fanout8695 (.X(net8695),
    .A(_11740_));
 sg13g2_buf_2 fanout8696 (.A(net8697),
    .X(net8696));
 sg13g2_buf_4 fanout8697 (.X(net8697),
    .A(_11739_));
 sg13g2_buf_2 fanout8698 (.A(net8700),
    .X(net8698));
 sg13g2_buf_2 fanout8699 (.A(net8700),
    .X(net8699));
 sg13g2_buf_4 fanout8700 (.X(net8700),
    .A(_11739_));
 sg13g2_buf_2 fanout8701 (.A(net8702),
    .X(net8701));
 sg13g2_buf_4 fanout8702 (.X(net8702),
    .A(_11735_));
 sg13g2_buf_2 fanout8703 (.A(net8705),
    .X(net8703));
 sg13g2_buf_2 fanout8704 (.A(net8705),
    .X(net8704));
 sg13g2_buf_4 fanout8705 (.X(net8705),
    .A(_11735_));
 sg13g2_buf_4 fanout8706 (.X(net8706),
    .A(net8707));
 sg13g2_buf_4 fanout8707 (.X(net8707),
    .A(_11734_));
 sg13g2_buf_4 fanout8708 (.X(net8708),
    .A(_11734_));
 sg13g2_buf_4 fanout8709 (.X(net8709),
    .A(_11064_));
 sg13g2_buf_2 fanout8710 (.A(_11064_),
    .X(net8710));
 sg13g2_buf_2 fanout8711 (.A(_11063_),
    .X(net8711));
 sg13g2_buf_4 fanout8712 (.X(net8712),
    .A(net8716));
 sg13g2_buf_2 fanout8713 (.A(net8714),
    .X(net8713));
 sg13g2_buf_2 fanout8714 (.A(net8715),
    .X(net8714));
 sg13g2_buf_2 fanout8715 (.A(net8716),
    .X(net8715));
 sg13g2_buf_4 fanout8716 (.X(net8716),
    .A(_10983_));
 sg13g2_buf_2 fanout8717 (.A(net8718),
    .X(net8717));
 sg13g2_buf_4 fanout8718 (.X(net8718),
    .A(net8719));
 sg13g2_buf_8 fanout8719 (.A(net8722),
    .X(net8719));
 sg13g2_buf_2 fanout8720 (.A(net8721),
    .X(net8720));
 sg13g2_buf_4 fanout8721 (.X(net8721),
    .A(net8722));
 sg13g2_buf_4 fanout8722 (.X(net8722),
    .A(_10982_));
 sg13g2_buf_4 fanout8723 (.X(net8723),
    .A(net8724));
 sg13g2_buf_4 fanout8724 (.X(net8724),
    .A(_10864_));
 sg13g2_buf_2 fanout8725 (.A(net8726),
    .X(net8725));
 sg13g2_buf_2 fanout8726 (.A(net8728),
    .X(net8726));
 sg13g2_buf_2 fanout8727 (.A(net8728),
    .X(net8727));
 sg13g2_buf_2 fanout8728 (.A(_10864_),
    .X(net8728));
 sg13g2_buf_2 fanout8729 (.A(net8732),
    .X(net8729));
 sg13g2_buf_2 fanout8730 (.A(net8731),
    .X(net8730));
 sg13g2_buf_2 fanout8731 (.A(net8732),
    .X(net8731));
 sg13g2_buf_2 fanout8732 (.A(_10845_),
    .X(net8732));
 sg13g2_buf_2 fanout8733 (.A(net8735),
    .X(net8733));
 sg13g2_buf_2 fanout8734 (.A(net8735),
    .X(net8734));
 sg13g2_buf_4 fanout8735 (.X(net8735),
    .A(net8737));
 sg13g2_buf_4 fanout8736 (.X(net8736),
    .A(net8737));
 sg13g2_buf_2 fanout8737 (.A(net8738),
    .X(net8737));
 sg13g2_buf_4 fanout8738 (.X(net8738),
    .A(_10845_));
 sg13g2_buf_4 fanout8739 (.X(net8739),
    .A(net8744));
 sg13g2_buf_4 fanout8740 (.X(net8740),
    .A(net8741));
 sg13g2_buf_2 fanout8741 (.A(net8742),
    .X(net8741));
 sg13g2_buf_2 fanout8742 (.A(net8743),
    .X(net8742));
 sg13g2_buf_4 fanout8743 (.X(net8743),
    .A(net8744));
 sg13g2_buf_4 fanout8744 (.X(net8744),
    .A(_10844_));
 sg13g2_buf_8 fanout8745 (.A(net8748),
    .X(net8745));
 sg13g2_buf_8 fanout8746 (.A(net8748),
    .X(net8746));
 sg13g2_buf_4 fanout8747 (.X(net8747),
    .A(net8748));
 sg13g2_buf_8 fanout8748 (.A(_09190_),
    .X(net8748));
 sg13g2_buf_2 fanout8749 (.A(net8750),
    .X(net8749));
 sg13g2_buf_4 fanout8750 (.X(net8750),
    .A(net8751));
 sg13g2_buf_2 fanout8751 (.A(net8755),
    .X(net8751));
 sg13g2_buf_4 fanout8752 (.X(net8752),
    .A(net8754));
 sg13g2_buf_2 fanout8753 (.A(net8754),
    .X(net8753));
 sg13g2_buf_2 fanout8754 (.A(net8755),
    .X(net8754));
 sg13g2_buf_2 fanout8755 (.A(net8768),
    .X(net8755));
 sg13g2_buf_4 fanout8756 (.X(net8756),
    .A(net8758));
 sg13g2_buf_2 fanout8757 (.A(net8758),
    .X(net8757));
 sg13g2_buf_2 fanout8758 (.A(net8768),
    .X(net8758));
 sg13g2_buf_4 fanout8759 (.X(net8759),
    .A(net8760));
 sg13g2_buf_2 fanout8760 (.A(net8768),
    .X(net8760));
 sg13g2_buf_4 fanout8761 (.X(net8761),
    .A(net8762));
 sg13g2_buf_4 fanout8762 (.X(net8762),
    .A(net8767));
 sg13g2_buf_4 fanout8763 (.X(net8763),
    .A(net8764));
 sg13g2_buf_4 fanout8764 (.X(net8764),
    .A(net8767));
 sg13g2_buf_4 fanout8765 (.X(net8765),
    .A(net8766));
 sg13g2_buf_4 fanout8766 (.X(net8766),
    .A(net8767));
 sg13g2_buf_2 fanout8767 (.A(net8768),
    .X(net8767));
 sg13g2_buf_8 fanout8768 (.A(_08544_),
    .X(net8768));
 sg13g2_buf_4 fanout8769 (.X(net8769),
    .A(net8778));
 sg13g2_buf_2 fanout8770 (.A(net8778),
    .X(net8770));
 sg13g2_buf_4 fanout8771 (.X(net8771),
    .A(net8772));
 sg13g2_buf_2 fanout8772 (.A(net8778),
    .X(net8772));
 sg13g2_buf_4 fanout8773 (.X(net8773),
    .A(net8778));
 sg13g2_buf_2 fanout8774 (.A(net8778),
    .X(net8774));
 sg13g2_buf_4 fanout8775 (.X(net8775),
    .A(net8777));
 sg13g2_buf_2 fanout8776 (.A(net8777),
    .X(net8776));
 sg13g2_buf_2 fanout8777 (.A(net8778),
    .X(net8777));
 sg13g2_buf_4 fanout8778 (.X(net8778),
    .A(_08544_));
 sg13g2_buf_4 fanout8779 (.X(net8779),
    .A(net8780));
 sg13g2_buf_2 fanout8780 (.A(net8795),
    .X(net8780));
 sg13g2_buf_4 fanout8781 (.X(net8781),
    .A(net8784));
 sg13g2_buf_2 fanout8782 (.A(net8784),
    .X(net8782));
 sg13g2_buf_2 fanout8783 (.A(net8784),
    .X(net8783));
 sg13g2_buf_2 fanout8784 (.A(net8795),
    .X(net8784));
 sg13g2_buf_4 fanout8785 (.X(net8785),
    .A(net8789));
 sg13g2_buf_2 fanout8786 (.A(net8789),
    .X(net8786));
 sg13g2_buf_4 fanout8787 (.X(net8787),
    .A(net8789));
 sg13g2_buf_2 fanout8788 (.A(net8789),
    .X(net8788));
 sg13g2_buf_2 fanout8789 (.A(net8795),
    .X(net8789));
 sg13g2_buf_4 fanout8790 (.X(net8790),
    .A(net8791));
 sg13g2_buf_4 fanout8791 (.X(net8791),
    .A(net8794));
 sg13g2_buf_4 fanout8792 (.X(net8792),
    .A(net8793));
 sg13g2_buf_4 fanout8793 (.X(net8793),
    .A(net8794));
 sg13g2_buf_2 fanout8794 (.A(net8795),
    .X(net8794));
 sg13g2_buf_4 fanout8795 (.X(net8795),
    .A(_08544_));
 sg13g2_buf_2 fanout8796 (.A(net8797),
    .X(net8796));
 sg13g2_buf_2 fanout8797 (.A(net8798),
    .X(net8797));
 sg13g2_buf_2 fanout8798 (.A(_06858_),
    .X(net8798));
 sg13g2_buf_4 fanout8799 (.X(net8799),
    .A(net8800));
 sg13g2_buf_2 fanout8800 (.A(net3401),
    .X(net8800));
 sg13g2_buf_4 fanout8801 (.X(net8801),
    .A(net8804));
 sg13g2_buf_4 fanout8802 (.X(net8802),
    .A(net8804));
 sg13g2_buf_2 fanout8803 (.A(net8804),
    .X(net8803));
 sg13g2_buf_4 fanout8804 (.X(net8804),
    .A(net8807));
 sg13g2_buf_4 fanout8805 (.X(net8805),
    .A(net8806));
 sg13g2_buf_8 fanout8806 (.A(net8807),
    .X(net8806));
 sg13g2_buf_4 fanout8807 (.X(net8807),
    .A(_04251_));
 sg13g2_buf_4 fanout8808 (.X(net8808),
    .A(net8810));
 sg13g2_buf_2 fanout8809 (.A(net8810),
    .X(net8809));
 sg13g2_buf_4 fanout8810 (.X(net8810),
    .A(net8818));
 sg13g2_buf_4 fanout8811 (.X(net8811),
    .A(net8818));
 sg13g2_buf_4 fanout8812 (.X(net8812),
    .A(net8818));
 sg13g2_buf_2 fanout8813 (.A(net8818),
    .X(net8813));
 sg13g2_buf_4 fanout8814 (.X(net8814),
    .A(net8817));
 sg13g2_buf_4 fanout8815 (.X(net8815),
    .A(net8817));
 sg13g2_buf_4 fanout8816 (.X(net8816),
    .A(net8817));
 sg13g2_buf_4 fanout8817 (.X(net8817),
    .A(net8818));
 sg13g2_buf_8 fanout8818 (.A(_02889_),
    .X(net8818));
 sg13g2_buf_2 fanout8819 (.A(_14120_),
    .X(net8819));
 sg13g2_buf_4 fanout8820 (.X(net8820),
    .A(net8821));
 sg13g2_buf_4 fanout8821 (.X(net8821),
    .A(net8822));
 sg13g2_buf_2 fanout8822 (.A(_13836_),
    .X(net8822));
 sg13g2_buf_4 fanout8823 (.X(net8823),
    .A(net8827));
 sg13g2_buf_2 fanout8824 (.A(net8827),
    .X(net8824));
 sg13g2_buf_4 fanout8825 (.X(net8825),
    .A(net8827));
 sg13g2_buf_2 fanout8826 (.A(net8827),
    .X(net8826));
 sg13g2_buf_2 fanout8827 (.A(_13836_),
    .X(net8827));
 sg13g2_buf_2 fanout8828 (.A(net8831),
    .X(net8828));
 sg13g2_buf_1 fanout8829 (.A(net8831),
    .X(net8829));
 sg13g2_buf_2 fanout8830 (.A(net8831),
    .X(net8830));
 sg13g2_buf_2 fanout8831 (.A(_13796_),
    .X(net8831));
 sg13g2_buf_4 fanout8832 (.X(net8832),
    .A(_13207_));
 sg13g2_buf_2 fanout8833 (.A(net8835),
    .X(net8833));
 sg13g2_buf_2 fanout8834 (.A(net8835),
    .X(net8834));
 sg13g2_buf_2 fanout8835 (.A(_13207_),
    .X(net8835));
 sg13g2_buf_2 fanout8836 (.A(net8837),
    .X(net8836));
 sg13g2_buf_2 fanout8837 (.A(_11736_),
    .X(net8837));
 sg13g2_buf_2 fanout8838 (.A(net8841),
    .X(net8838));
 sg13g2_buf_2 fanout8839 (.A(net8841),
    .X(net8839));
 sg13g2_buf_1 fanout8840 (.A(net8841),
    .X(net8840));
 sg13g2_buf_4 fanout8841 (.X(net8841),
    .A(_11736_));
 sg13g2_buf_4 fanout8842 (.X(net8842),
    .A(_10974_));
 sg13g2_buf_4 fanout8843 (.X(net8843),
    .A(_10974_));
 sg13g2_buf_2 fanout8844 (.A(net8845),
    .X(net8844));
 sg13g2_buf_2 fanout8845 (.A(net8846),
    .X(net8845));
 sg13g2_buf_4 fanout8846 (.X(net8846),
    .A(net8853));
 sg13g2_buf_2 fanout8847 (.A(net8848),
    .X(net8847));
 sg13g2_buf_2 fanout8848 (.A(net8849),
    .X(net8848));
 sg13g2_buf_2 fanout8849 (.A(net8853),
    .X(net8849));
 sg13g2_buf_2 fanout8850 (.A(net8851),
    .X(net8850));
 sg13g2_buf_2 fanout8851 (.A(net8852),
    .X(net8851));
 sg13g2_buf_2 fanout8852 (.A(net8853),
    .X(net8852));
 sg13g2_buf_8 fanout8853 (.A(_10973_),
    .X(net8853));
 sg13g2_buf_4 fanout8854 (.X(net8854),
    .A(net8855));
 sg13g2_buf_2 fanout8855 (.A(_10854_),
    .X(net8855));
 sg13g2_buf_4 fanout8856 (.X(net8856),
    .A(net8857));
 sg13g2_buf_2 fanout8857 (.A(net8858),
    .X(net8857));
 sg13g2_buf_2 fanout8858 (.A(net8859),
    .X(net8858));
 sg13g2_buf_4 fanout8859 (.X(net8859),
    .A(_10854_));
 sg13g2_buf_2 fanout8860 (.A(net8862),
    .X(net8860));
 sg13g2_buf_2 fanout8861 (.A(net8862),
    .X(net8861));
 sg13g2_buf_4 fanout8862 (.X(net8862),
    .A(net8871));
 sg13g2_buf_4 fanout8863 (.X(net8863),
    .A(net8865));
 sg13g2_buf_2 fanout8864 (.A(net8865),
    .X(net8864));
 sg13g2_buf_2 fanout8865 (.A(net8871),
    .X(net8865));
 sg13g2_buf_4 fanout8866 (.X(net8866),
    .A(net8867));
 sg13g2_buf_4 fanout8867 (.X(net8867),
    .A(net8868));
 sg13g2_buf_2 fanout8868 (.A(net8871),
    .X(net8868));
 sg13g2_buf_4 fanout8869 (.X(net8869),
    .A(net8870));
 sg13g2_buf_2 fanout8870 (.A(net8871),
    .X(net8870));
 sg13g2_buf_4 fanout8871 (.X(net8871),
    .A(net8906));
 sg13g2_buf_4 fanout8872 (.X(net8872),
    .A(net8873));
 sg13g2_buf_4 fanout8873 (.X(net8873),
    .A(net8877));
 sg13g2_buf_4 fanout8874 (.X(net8874),
    .A(net8875));
 sg13g2_buf_4 fanout8875 (.X(net8875),
    .A(net8877));
 sg13g2_buf_4 fanout8876 (.X(net8876),
    .A(net8877));
 sg13g2_buf_4 fanout8877 (.X(net8877),
    .A(net8906));
 sg13g2_buf_4 fanout8878 (.X(net8878),
    .A(net8887));
 sg13g2_buf_2 fanout8879 (.A(net8887),
    .X(net8879));
 sg13g2_buf_4 fanout8880 (.X(net8880),
    .A(net8881));
 sg13g2_buf_2 fanout8881 (.A(net8887),
    .X(net8881));
 sg13g2_buf_4 fanout8882 (.X(net8882),
    .A(net8887));
 sg13g2_buf_2 fanout8883 (.A(net8887),
    .X(net8883));
 sg13g2_buf_4 fanout8884 (.X(net8884),
    .A(net8886));
 sg13g2_buf_2 fanout8885 (.A(net8886),
    .X(net8885));
 sg13g2_buf_2 fanout8886 (.A(net8887),
    .X(net8886));
 sg13g2_buf_4 fanout8887 (.X(net8887),
    .A(net8906));
 sg13g2_buf_4 fanout8888 (.X(net8888),
    .A(net8889));
 sg13g2_buf_4 fanout8889 (.X(net8889),
    .A(net8894));
 sg13g2_buf_4 fanout8890 (.X(net8890),
    .A(net8893));
 sg13g2_buf_4 fanout8891 (.X(net8891),
    .A(net8893));
 sg13g2_buf_2 fanout8892 (.A(net8893),
    .X(net8892));
 sg13g2_buf_2 fanout8893 (.A(net8894),
    .X(net8893));
 sg13g2_buf_2 fanout8894 (.A(net8905),
    .X(net8894));
 sg13g2_buf_4 fanout8895 (.X(net8895),
    .A(net8899));
 sg13g2_buf_2 fanout8896 (.A(net8899),
    .X(net8896));
 sg13g2_buf_4 fanout8897 (.X(net8897),
    .A(net8899));
 sg13g2_buf_2 fanout8898 (.A(net8899),
    .X(net8898));
 sg13g2_buf_1 fanout8899 (.A(net8905),
    .X(net8899));
 sg13g2_buf_4 fanout8900 (.X(net8900),
    .A(net8902));
 sg13g2_buf_2 fanout8901 (.A(net8902),
    .X(net8901));
 sg13g2_buf_4 fanout8902 (.X(net8902),
    .A(net8905));
 sg13g2_buf_4 fanout8903 (.X(net8903),
    .A(net8904));
 sg13g2_buf_4 fanout8904 (.X(net8904),
    .A(net8905));
 sg13g2_buf_4 fanout8905 (.X(net8905),
    .A(net8906));
 sg13g2_buf_8 fanout8906 (.A(_08581_),
    .X(net8906));
 sg13g2_buf_4 fanout8907 (.X(net8907),
    .A(net8910));
 sg13g2_buf_4 fanout8908 (.X(net8908),
    .A(net8910));
 sg13g2_buf_8 fanout8909 (.A(net8910),
    .X(net8909));
 sg13g2_buf_8 fanout8910 (.A(net8916),
    .X(net8910));
 sg13g2_buf_8 fanout8911 (.A(net8916),
    .X(net8911));
 sg13g2_buf_4 fanout8912 (.X(net8912),
    .A(net8916));
 sg13g2_buf_4 fanout8913 (.X(net8913),
    .A(net8915));
 sg13g2_buf_4 fanout8914 (.X(net8914),
    .A(net8915));
 sg13g2_buf_8 fanout8915 (.A(net8916),
    .X(net8915));
 sg13g2_buf_8 fanout8916 (.A(_08543_),
    .X(net8916));
 sg13g2_buf_8 fanout8917 (.A(_08537_),
    .X(net8917));
 sg13g2_buf_4 fanout8918 (.X(net8918),
    .A(_08537_));
 sg13g2_buf_8 fanout8919 (.A(net8921),
    .X(net8919));
 sg13g2_buf_4 fanout8920 (.X(net8920),
    .A(net8921));
 sg13g2_buf_8 fanout8921 (.A(_08537_),
    .X(net8921));
 sg13g2_buf_8 fanout8922 (.A(net8923),
    .X(net8922));
 sg13g2_buf_8 fanout8923 (.A(net8928),
    .X(net8923));
 sg13g2_buf_2 fanout8924 (.A(net8928),
    .X(net8924));
 sg13g2_buf_8 fanout8925 (.A(net8928),
    .X(net8925));
 sg13g2_buf_8 fanout8926 (.A(net8927),
    .X(net8926));
 sg13g2_buf_8 fanout8927 (.A(net8928),
    .X(net8927));
 sg13g2_buf_8 fanout8928 (.A(_08536_),
    .X(net8928));
 sg13g2_buf_2 fanout8929 (.A(_07039_),
    .X(net8929));
 sg13g2_buf_1 fanout8930 (.A(_07039_),
    .X(net8930));
 sg13g2_buf_2 fanout8931 (.A(net8932),
    .X(net8931));
 sg13g2_buf_2 fanout8932 (.A(net8933),
    .X(net8932));
 sg13g2_buf_2 fanout8933 (.A(_07038_),
    .X(net8933));
 sg13g2_buf_2 fanout8934 (.A(_06961_),
    .X(net8934));
 sg13g2_buf_1 fanout8935 (.A(_06961_),
    .X(net8935));
 sg13g2_buf_4 fanout8936 (.X(net8936),
    .A(net8938));
 sg13g2_buf_2 fanout8937 (.A(net8938),
    .X(net8937));
 sg13g2_buf_2 fanout8938 (.A(_06960_),
    .X(net8938));
 sg13g2_buf_4 fanout8939 (.X(net8939),
    .A(_05026_));
 sg13g2_buf_2 fanout8940 (.A(net8941),
    .X(net8940));
 sg13g2_buf_2 fanout8941 (.A(net8942),
    .X(net8941));
 sg13g2_buf_2 fanout8942 (.A(net8944),
    .X(net8942));
 sg13g2_buf_4 fanout8943 (.X(net8943),
    .A(net8944));
 sg13g2_buf_2 fanout8944 (.A(_05025_),
    .X(net8944));
 sg13g2_buf_2 fanout8945 (.A(_04427_),
    .X(net8945));
 sg13g2_buf_4 fanout8946 (.X(net8946),
    .A(net8947));
 sg13g2_buf_4 fanout8947 (.X(net8947),
    .A(net8949));
 sg13g2_buf_4 fanout8948 (.X(net8948),
    .A(net8949));
 sg13g2_buf_4 fanout8949 (.X(net8949),
    .A(_02893_));
 sg13g2_buf_8 fanout8950 (.A(net8955),
    .X(net8950));
 sg13g2_buf_4 fanout8951 (.X(net8951),
    .A(net8955));
 sg13g2_buf_4 fanout8952 (.X(net8952),
    .A(net8953));
 sg13g2_buf_4 fanout8953 (.X(net8953),
    .A(net8955));
 sg13g2_buf_4 fanout8954 (.X(net8954),
    .A(net8955));
 sg13g2_buf_4 fanout8955 (.X(net8955),
    .A(_02893_));
 sg13g2_buf_4 fanout8956 (.X(net8956),
    .A(net8957));
 sg13g2_buf_2 fanout8957 (.A(_13835_),
    .X(net8957));
 sg13g2_buf_4 fanout8958 (.X(net8958),
    .A(net8959));
 sg13g2_buf_4 fanout8959 (.X(net8959),
    .A(_13834_));
 sg13g2_buf_4 fanout8960 (.X(net8960),
    .A(_12880_));
 sg13g2_buf_2 fanout8961 (.A(_12608_),
    .X(net8961));
 sg13g2_buf_8 fanout8962 (.A(_10915_),
    .X(net8962));
 sg13g2_buf_2 fanout8963 (.A(net8964),
    .X(net8963));
 sg13g2_buf_2 fanout8964 (.A(net8971),
    .X(net8964));
 sg13g2_buf_2 fanout8965 (.A(net8967),
    .X(net8965));
 sg13g2_buf_2 fanout8966 (.A(net8967),
    .X(net8966));
 sg13g2_buf_4 fanout8967 (.X(net8967),
    .A(net8971));
 sg13g2_buf_4 fanout8968 (.X(net8968),
    .A(net8970));
 sg13g2_buf_2 fanout8969 (.A(net8970),
    .X(net8969));
 sg13g2_buf_2 fanout8970 (.A(net8971),
    .X(net8970));
 sg13g2_buf_4 fanout8971 (.X(net8971),
    .A(net8972));
 sg13g2_buf_4 fanout8972 (.X(net8972),
    .A(_10913_));
 sg13g2_buf_2 fanout8973 (.A(_10853_),
    .X(net8973));
 sg13g2_buf_2 fanout8974 (.A(_10848_),
    .X(net8974));
 sg13g2_buf_2 fanout8975 (.A(net8976),
    .X(net8975));
 sg13g2_buf_2 fanout8976 (.A(_10840_),
    .X(net8976));
 sg13g2_buf_2 fanout8977 (.A(_10839_),
    .X(net8977));
 sg13g2_buf_4 fanout8978 (.X(net8978),
    .A(_10838_));
 sg13g2_buf_2 fanout8979 (.A(_10835_),
    .X(net8979));
 sg13g2_buf_2 fanout8980 (.A(_10833_),
    .X(net8980));
 sg13g2_buf_4 fanout8981 (.X(net8981),
    .A(_10674_));
 sg13g2_buf_2 fanout8982 (.A(_10674_),
    .X(net8982));
 sg13g2_buf_4 fanout8983 (.X(net8983),
    .A(_10607_));
 sg13g2_buf_4 fanout8984 (.X(net8984),
    .A(_10606_));
 sg13g2_buf_2 fanout8985 (.A(_10606_),
    .X(net8985));
 sg13g2_buf_4 fanout8986 (.X(net8986),
    .A(net8987));
 sg13g2_buf_4 fanout8987 (.X(net8987),
    .A(_10606_));
 sg13g2_buf_2 fanout8988 (.A(net8989),
    .X(net8988));
 sg13g2_buf_2 fanout8989 (.A(net8990),
    .X(net8989));
 sg13g2_buf_2 fanout8990 (.A(net8991),
    .X(net8990));
 sg13g2_buf_4 fanout8991 (.X(net8991),
    .A(_10605_));
 sg13g2_buf_2 fanout8992 (.A(net8993),
    .X(net8992));
 sg13g2_buf_4 fanout8993 (.X(net8993),
    .A(net8994));
 sg13g2_buf_4 fanout8994 (.X(net8994),
    .A(_10605_));
 sg13g2_buf_2 fanout8995 (.A(net8997),
    .X(net8995));
 sg13g2_buf_2 fanout8996 (.A(net8997),
    .X(net8996));
 sg13g2_buf_2 fanout8997 (.A(net8998),
    .X(net8997));
 sg13g2_buf_2 fanout8998 (.A(_10603_),
    .X(net8998));
 sg13g2_buf_2 fanout8999 (.A(net9000),
    .X(net8999));
 sg13g2_buf_2 fanout9000 (.A(_10603_),
    .X(net9000));
 sg13g2_buf_8 fanout9001 (.A(_10602_),
    .X(net9001));
 sg13g2_buf_2 fanout9002 (.A(net9003),
    .X(net9002));
 sg13g2_buf_4 fanout9003 (.X(net9003),
    .A(net9004));
 sg13g2_buf_4 fanout9004 (.X(net9004),
    .A(net9007));
 sg13g2_buf_4 fanout9005 (.X(net9005),
    .A(net9006));
 sg13g2_buf_4 fanout9006 (.X(net9006),
    .A(net9007));
 sg13g2_buf_2 fanout9007 (.A(net9015),
    .X(net9007));
 sg13g2_buf_4 fanout9008 (.X(net9008),
    .A(net9009));
 sg13g2_buf_4 fanout9009 (.X(net9009),
    .A(net9015));
 sg13g2_buf_2 fanout9010 (.A(net9011),
    .X(net9010));
 sg13g2_buf_2 fanout9011 (.A(net9012),
    .X(net9011));
 sg13g2_buf_2 fanout9012 (.A(net9015),
    .X(net9012));
 sg13g2_buf_4 fanout9013 (.X(net9013),
    .A(net9014));
 sg13g2_buf_4 fanout9014 (.X(net9014),
    .A(net9015));
 sg13g2_buf_4 fanout9015 (.X(net9015),
    .A(net9034));
 sg13g2_buf_4 fanout9016 (.X(net9016),
    .A(net9020));
 sg13g2_buf_4 fanout9017 (.X(net9017),
    .A(net9020));
 sg13g2_buf_2 fanout9018 (.A(net9019),
    .X(net9018));
 sg13g2_buf_4 fanout9019 (.X(net9019),
    .A(net9020));
 sg13g2_buf_2 fanout9020 (.A(net9021),
    .X(net9020));
 sg13g2_buf_4 fanout9021 (.X(net9021),
    .A(net9034));
 sg13g2_buf_4 fanout9022 (.X(net9022),
    .A(net9026));
 sg13g2_buf_2 fanout9023 (.A(net9025),
    .X(net9023));
 sg13g2_buf_2 fanout9024 (.A(net9025),
    .X(net9024));
 sg13g2_buf_4 fanout9025 (.X(net9025),
    .A(net9026));
 sg13g2_buf_4 fanout9026 (.X(net9026),
    .A(net9034));
 sg13g2_buf_4 fanout9027 (.X(net9027),
    .A(net9033));
 sg13g2_buf_2 fanout9028 (.A(net9033),
    .X(net9028));
 sg13g2_buf_4 fanout9029 (.X(net9029),
    .A(net9033));
 sg13g2_buf_2 fanout9030 (.A(net9032),
    .X(net9030));
 sg13g2_buf_4 fanout9031 (.X(net9031),
    .A(net9033));
 sg13g2_buf_2 fanout9032 (.A(net9033),
    .X(net9032));
 sg13g2_buf_4 fanout9033 (.X(net9033),
    .A(net9034));
 sg13g2_buf_4 fanout9034 (.X(net9034),
    .A(net9061));
 sg13g2_buf_2 fanout9035 (.A(net9036),
    .X(net9035));
 sg13g2_buf_2 fanout9036 (.A(net9037),
    .X(net9036));
 sg13g2_buf_4 fanout9037 (.X(net9037),
    .A(net9039));
 sg13g2_buf_4 fanout9038 (.X(net9038),
    .A(net9039));
 sg13g2_buf_2 fanout9039 (.A(net9053),
    .X(net9039));
 sg13g2_buf_4 fanout9040 (.X(net9040),
    .A(net9043));
 sg13g2_buf_2 fanout9041 (.A(net9042),
    .X(net9041));
 sg13g2_buf_2 fanout9042 (.A(net9043),
    .X(net9042));
 sg13g2_buf_2 fanout9043 (.A(net9053),
    .X(net9043));
 sg13g2_buf_2 fanout9044 (.A(net9045),
    .X(net9044));
 sg13g2_buf_4 fanout9045 (.X(net9045),
    .A(net9053));
 sg13g2_buf_2 fanout9046 (.A(net9049),
    .X(net9046));
 sg13g2_buf_2 fanout9047 (.A(net9049),
    .X(net9047));
 sg13g2_buf_2 fanout9048 (.A(net9049),
    .X(net9048));
 sg13g2_buf_2 fanout9049 (.A(net9053),
    .X(net9049));
 sg13g2_buf_2 fanout9050 (.A(net9051),
    .X(net9050));
 sg13g2_buf_4 fanout9051 (.X(net9051),
    .A(net9052));
 sg13g2_buf_4 fanout9052 (.X(net9052),
    .A(net9053));
 sg13g2_buf_8 fanout9053 (.A(net9061),
    .X(net9053));
 sg13g2_buf_4 fanout9054 (.X(net9054),
    .A(net9055));
 sg13g2_buf_4 fanout9055 (.X(net9055),
    .A(net9061));
 sg13g2_buf_4 fanout9056 (.X(net9056),
    .A(net9059));
 sg13g2_buf_2 fanout9057 (.A(net9058),
    .X(net9057));
 sg13g2_buf_4 fanout9058 (.X(net9058),
    .A(net9059));
 sg13g2_buf_2 fanout9059 (.A(net9060),
    .X(net9059));
 sg13g2_buf_4 fanout9060 (.X(net9060),
    .A(net9061));
 sg13g2_buf_8 fanout9061 (.A(_10593_),
    .X(net9061));
 sg13g2_buf_2 fanout9062 (.A(net9064),
    .X(net9062));
 sg13g2_buf_4 fanout9063 (.X(net9063),
    .A(net9064));
 sg13g2_buf_4 fanout9064 (.X(net9064),
    .A(_10513_));
 sg13g2_buf_2 fanout9065 (.A(net9066),
    .X(net9065));
 sg13g2_buf_2 fanout9066 (.A(_10512_),
    .X(net9066));
 sg13g2_buf_2 fanout9067 (.A(net9068),
    .X(net9067));
 sg13g2_buf_2 fanout9068 (.A(net9070),
    .X(net9068));
 sg13g2_buf_2 fanout9069 (.A(net9070),
    .X(net9069));
 sg13g2_buf_2 fanout9070 (.A(_10511_),
    .X(net9070));
 sg13g2_buf_2 fanout9071 (.A(net9073),
    .X(net9071));
 sg13g2_buf_4 fanout9072 (.X(net9072),
    .A(net9073));
 sg13g2_buf_2 fanout9073 (.A(_10510_),
    .X(net9073));
 sg13g2_buf_4 fanout9074 (.X(net9074),
    .A(net9075));
 sg13g2_buf_4 fanout9075 (.X(net9075),
    .A(net9076));
 sg13g2_buf_4 fanout9076 (.X(net9076),
    .A(_10509_));
 sg13g2_buf_4 fanout9077 (.X(net9077),
    .A(net9078));
 sg13g2_buf_4 fanout9078 (.X(net9078),
    .A(_10508_));
 sg13g2_buf_2 fanout9079 (.A(net9080),
    .X(net9079));
 sg13g2_buf_4 fanout9080 (.X(net9080),
    .A(net9091));
 sg13g2_buf_2 fanout9081 (.A(net9085),
    .X(net9081));
 sg13g2_buf_4 fanout9082 (.X(net9082),
    .A(net9084));
 sg13g2_buf_1 fanout9083 (.A(net9084),
    .X(net9083));
 sg13g2_buf_2 fanout9084 (.A(net9085),
    .X(net9084));
 sg13g2_buf_1 fanout9085 (.A(net9091),
    .X(net9085));
 sg13g2_buf_2 fanout9086 (.A(net9087),
    .X(net9086));
 sg13g2_buf_2 fanout9087 (.A(net9091),
    .X(net9087));
 sg13g2_buf_2 fanout9088 (.A(net9090),
    .X(net9088));
 sg13g2_buf_1 fanout9089 (.A(net9090),
    .X(net9089));
 sg13g2_buf_2 fanout9090 (.A(net9091),
    .X(net9090));
 sg13g2_buf_8 fanout9091 (.A(_10464_),
    .X(net9091));
 sg13g2_buf_4 fanout9092 (.X(net9092),
    .A(net9095));
 sg13g2_buf_2 fanout9093 (.A(net9094),
    .X(net9093));
 sg13g2_buf_4 fanout9094 (.X(net9094),
    .A(net9095));
 sg13g2_buf_1 fanout9095 (.A(_10464_),
    .X(net9095));
 sg13g2_buf_2 fanout9096 (.A(net9098),
    .X(net9096));
 sg13g2_buf_1 fanout9097 (.A(net9098),
    .X(net9097));
 sg13g2_buf_2 fanout9098 (.A(net9107),
    .X(net9098));
 sg13g2_buf_4 fanout9099 (.X(net9099),
    .A(net9107));
 sg13g2_buf_2 fanout9100 (.A(net9107),
    .X(net9100));
 sg13g2_buf_4 fanout9101 (.X(net9101),
    .A(net9102));
 sg13g2_buf_4 fanout9102 (.X(net9102),
    .A(net9106));
 sg13g2_buf_4 fanout9103 (.X(net9103),
    .A(net9104));
 sg13g2_buf_2 fanout9104 (.A(net9105),
    .X(net9104));
 sg13g2_buf_4 fanout9105 (.X(net9105),
    .A(net9106));
 sg13g2_buf_2 fanout9106 (.A(net9107),
    .X(net9106));
 sg13g2_buf_2 fanout9107 (.A(_10464_),
    .X(net9107));
 sg13g2_buf_8 fanout9108 (.A(_10463_),
    .X(net9108));
 sg13g2_buf_4 fanout9109 (.X(net9109),
    .A(_10463_));
 sg13g2_buf_8 fanout9110 (.A(_10463_),
    .X(net9110));
 sg13g2_buf_4 fanout9111 (.X(net9111),
    .A(_10461_));
 sg13g2_buf_4 fanout9112 (.X(net9112),
    .A(_10461_));
 sg13g2_buf_8 fanout9113 (.A(net9114),
    .X(net9113));
 sg13g2_buf_4 fanout9114 (.X(net9114),
    .A(net9115));
 sg13g2_buf_8 fanout9115 (.A(_10461_),
    .X(net9115));
 sg13g2_buf_2 fanout9116 (.A(net9118),
    .X(net9116));
 sg13g2_buf_2 fanout9117 (.A(net9118),
    .X(net9117));
 sg13g2_buf_4 fanout9118 (.X(net9118),
    .A(net9119));
 sg13g2_buf_2 fanout9119 (.A(net9121),
    .X(net9119));
 sg13g2_buf_4 fanout9120 (.X(net9120),
    .A(net9121));
 sg13g2_buf_2 fanout9121 (.A(net9133),
    .X(net9121));
 sg13g2_buf_2 fanout9122 (.A(net9123),
    .X(net9122));
 sg13g2_buf_4 fanout9123 (.X(net9123),
    .A(net9124));
 sg13g2_buf_2 fanout9124 (.A(net9126),
    .X(net9124));
 sg13g2_buf_4 fanout9125 (.X(net9125),
    .A(net9126));
 sg13g2_buf_2 fanout9126 (.A(net9133),
    .X(net9126));
 sg13g2_buf_2 fanout9127 (.A(net9128),
    .X(net9127));
 sg13g2_buf_4 fanout9128 (.X(net9128),
    .A(net9133));
 sg13g2_buf_2 fanout9129 (.A(net9132),
    .X(net9129));
 sg13g2_buf_2 fanout9130 (.A(net9132),
    .X(net9130));
 sg13g2_buf_2 fanout9131 (.A(net9132),
    .X(net9131));
 sg13g2_buf_4 fanout9132 (.X(net9132),
    .A(net9133));
 sg13g2_buf_8 fanout9133 (.A(_10460_),
    .X(net9133));
 sg13g2_buf_4 fanout9134 (.X(net9134),
    .A(net9140));
 sg13g2_buf_4 fanout9135 (.X(net9135),
    .A(net9140));
 sg13g2_buf_4 fanout9136 (.X(net9136),
    .A(net9140));
 sg13g2_buf_2 fanout9137 (.A(net9140),
    .X(net9137));
 sg13g2_buf_4 fanout9138 (.X(net9138),
    .A(net9139));
 sg13g2_buf_4 fanout9139 (.X(net9139),
    .A(net9140));
 sg13g2_buf_2 fanout9140 (.A(_10460_),
    .X(net9140));
 sg13g2_buf_4 fanout9141 (.X(net9141),
    .A(net9142));
 sg13g2_buf_2 fanout9142 (.A(net9157),
    .X(net9142));
 sg13g2_buf_4 fanout9143 (.X(net9143),
    .A(net9146));
 sg13g2_buf_2 fanout9144 (.A(net9146),
    .X(net9144));
 sg13g2_buf_4 fanout9145 (.X(net9145),
    .A(net9146));
 sg13g2_buf_2 fanout9146 (.A(net9157),
    .X(net9146));
 sg13g2_buf_4 fanout9147 (.X(net9147),
    .A(net9150));
 sg13g2_buf_4 fanout9148 (.X(net9148),
    .A(net9150));
 sg13g2_buf_2 fanout9149 (.A(net9150),
    .X(net9149));
 sg13g2_buf_2 fanout9150 (.A(net9157),
    .X(net9150));
 sg13g2_buf_2 fanout9151 (.A(net9152),
    .X(net9151));
 sg13g2_buf_4 fanout9152 (.X(net9152),
    .A(net9157));
 sg13g2_buf_4 fanout9153 (.X(net9153),
    .A(net9156));
 sg13g2_buf_2 fanout9154 (.A(net9156),
    .X(net9154));
 sg13g2_buf_2 fanout9155 (.A(net9156),
    .X(net9155));
 sg13g2_buf_2 fanout9156 (.A(net9157),
    .X(net9156));
 sg13g2_buf_4 fanout9157 (.X(net9157),
    .A(_10460_));
 sg13g2_buf_4 fanout9158 (.X(net9158),
    .A(net9162));
 sg13g2_buf_4 fanout9159 (.X(net9159),
    .A(net9162));
 sg13g2_buf_8 fanout9160 (.A(net9162),
    .X(net9160));
 sg13g2_buf_2 fanout9161 (.A(net9162),
    .X(net9161));
 sg13g2_buf_8 fanout9162 (.A(_10459_),
    .X(net9162));
 sg13g2_buf_4 fanout9163 (.X(net9163),
    .A(net9169));
 sg13g2_buf_4 fanout9164 (.X(net9164),
    .A(net9168));
 sg13g2_buf_4 fanout9165 (.X(net9165),
    .A(net9166));
 sg13g2_buf_4 fanout9166 (.X(net9166),
    .A(net9167));
 sg13g2_buf_4 fanout9167 (.X(net9167),
    .A(net9168));
 sg13g2_buf_2 fanout9168 (.A(net9169),
    .X(net9168));
 sg13g2_buf_4 fanout9169 (.X(net9169),
    .A(_10459_));
 sg13g2_buf_4 fanout9170 (.X(net9170),
    .A(net9171));
 sg13g2_buf_4 fanout9171 (.X(net9171),
    .A(_10396_));
 sg13g2_buf_4 fanout9172 (.X(net9172),
    .A(net9176));
 sg13g2_buf_2 fanout9173 (.A(net9176),
    .X(net9173));
 sg13g2_buf_4 fanout9174 (.X(net9174),
    .A(net9176));
 sg13g2_buf_2 fanout9175 (.A(net9176),
    .X(net9175));
 sg13g2_buf_2 fanout9176 (.A(_00003_),
    .X(net9176));
 sg13g2_buf_4 fanout9177 (.X(net9177),
    .A(net9178));
 sg13g2_buf_4 fanout9178 (.X(net9178),
    .A(_00002_));
 sg13g2_buf_4 fanout9179 (.X(net9179),
    .A(_00001_));
 sg13g2_buf_4 fanout9180 (.X(net9180),
    .A(_00001_));
 sg13g2_buf_2 fanout9181 (.A(net9182),
    .X(net9181));
 sg13g2_buf_4 fanout9182 (.X(net9182),
    .A(net9183));
 sg13g2_buf_4 fanout9183 (.X(net9183),
    .A(_00001_));
 sg13g2_buf_4 fanout9184 (.X(net9184),
    .A(net9186));
 sg13g2_buf_4 fanout9185 (.X(net9185),
    .A(net9187));
 sg13g2_buf_2 fanout9186 (.A(net9187),
    .X(net9186));
 sg13g2_buf_8 fanout9187 (.A(net9194),
    .X(net9187));
 sg13g2_buf_2 fanout9188 (.A(net9192),
    .X(net9188));
 sg13g2_buf_2 fanout9189 (.A(net9192),
    .X(net9189));
 sg13g2_buf_4 fanout9190 (.X(net9190),
    .A(net9192));
 sg13g2_buf_4 fanout9191 (.X(net9191),
    .A(net9192));
 sg13g2_buf_2 fanout9192 (.A(net9193),
    .X(net9192));
 sg13g2_buf_4 fanout9193 (.X(net9193),
    .A(net9194));
 sg13g2_buf_4 fanout9194 (.X(net9194),
    .A(_00000_));
 sg13g2_buf_4 fanout9195 (.X(net9195),
    .A(\soc_I.qqspi_I.state[5] ));
 sg13g2_buf_2 fanout9196 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[0] ),
    .X(net9196));
 sg13g2_buf_2 fanout9197 (.A(net9198),
    .X(net9197));
 sg13g2_buf_2 fanout9198 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[1] ),
    .X(net9198));
 sg13g2_buf_2 fanout9199 (.A(net9200),
    .X(net9199));
 sg13g2_buf_2 fanout9200 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[2] ),
    .X(net9200));
 sg13g2_buf_2 fanout9201 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[3] ),
    .X(net9201));
 sg13g2_buf_2 fanout9202 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[4] ),
    .X(net9202));
 sg13g2_buf_2 fanout9203 (.A(net9204),
    .X(net9203));
 sg13g2_buf_4 fanout9204 (.X(net9204),
    .A(\soc_I.kianv_I.control_unit_I.main_fsm_I.state[5] ));
 sg13g2_buf_2 fanout9205 (.A(net5512),
    .X(net9205));
 sg13g2_buf_2 fanout9206 (.A(net5527),
    .X(net9206));
 sg13g2_buf_2 fanout9207 (.A(net9209),
    .X(net9207));
 sg13g2_buf_2 fanout9208 (.A(net9209),
    .X(net9208));
 sg13g2_buf_2 fanout9209 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.state[1] ),
    .X(net9209));
 sg13g2_buf_4 fanout9210 (.X(net9210),
    .A(net9211));
 sg13g2_buf_2 fanout9211 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.state[1] ),
    .X(net9211));
 sg13g2_buf_2 fanout9212 (.A(net9213),
    .X(net9212));
 sg13g2_buf_4 fanout9213 (.X(net9213),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.state[1] ));
 sg13g2_buf_2 fanout9214 (.A(net9216),
    .X(net9214));
 sg13g2_buf_4 fanout9215 (.X(net9215),
    .A(net9217));
 sg13g2_buf_2 fanout9216 (.A(net9217),
    .X(net9216));
 sg13g2_buf_4 fanout9217 (.X(net9217),
    .A(net9223));
 sg13g2_buf_4 fanout9218 (.X(net9218),
    .A(net9223));
 sg13g2_buf_2 fanout9219 (.A(net9223),
    .X(net9219));
 sg13g2_buf_4 fanout9220 (.X(net9220),
    .A(net9222));
 sg13g2_buf_2 fanout9221 (.A(net9222),
    .X(net9221));
 sg13g2_buf_2 fanout9222 (.A(net9223),
    .X(net9222));
 sg13g2_buf_4 fanout9223 (.X(net9223),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.state[2] ));
 sg13g2_buf_2 fanout9224 (.A(net9225),
    .X(net9224));
 sg13g2_buf_1 fanout9225 (.A(net9231),
    .X(net9225));
 sg13g2_buf_2 fanout9226 (.A(net9231),
    .X(net9226));
 sg13g2_buf_2 fanout9227 (.A(net9231),
    .X(net9227));
 sg13g2_buf_2 fanout9228 (.A(net9230),
    .X(net9228));
 sg13g2_buf_2 fanout9229 (.A(net9230),
    .X(net9229));
 sg13g2_buf_2 fanout9230 (.A(net9231),
    .X(net9230));
 sg13g2_buf_4 fanout9231 (.X(net9231),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.div_state[1] ));
 sg13g2_buf_4 fanout9232 (.X(net9232),
    .A(net9236));
 sg13g2_buf_4 fanout9233 (.X(net9233),
    .A(net9234));
 sg13g2_buf_2 fanout9234 (.A(net9235),
    .X(net9234));
 sg13g2_buf_2 fanout9235 (.A(net9236),
    .X(net9235));
 sg13g2_buf_2 fanout9236 (.A(_00184_),
    .X(net9236));
 sg13g2_buf_2 fanout9237 (.A(net9239),
    .X(net9237));
 sg13g2_buf_2 fanout9238 (.A(net9239),
    .X(net9238));
 sg13g2_buf_4 fanout9239 (.X(net9239),
    .A(\soc_I.kianv_I.datapath_unit_I.div_I.div_state[2] ));
 sg13g2_buf_2 fanout9240 (.A(net9241),
    .X(net9240));
 sg13g2_buf_2 fanout9241 (.A(net9242),
    .X(net9241));
 sg13g2_buf_4 fanout9242 (.X(net9242),
    .A(\soc_I.rx_uart_i.data_rd ));
 sg13g2_buf_2 fanout9243 (.A(net9244),
    .X(net9243));
 sg13g2_buf_2 fanout9244 (.A(net9245),
    .X(net9244));
 sg13g2_buf_4 fanout9245 (.X(net9245),
    .A(net5521));
 sg13g2_buf_2 fanout9246 (.A(net9247),
    .X(net9246));
 sg13g2_buf_2 fanout9247 (.A(net9248),
    .X(net9247));
 sg13g2_buf_2 fanout9248 (.A(\soc_I.uart_tx_ready ),
    .X(net9248));
 sg13g2_buf_2 fanout9249 (.A(net9250),
    .X(net9249));
 sg13g2_buf_2 fanout9250 (.A(net9251),
    .X(net9250));
 sg13g2_buf_2 fanout9251 (.A(\soc_I.uart_tx_ready ),
    .X(net9251));
 sg13g2_buf_2 fanout9252 (.A(net9253),
    .X(net9252));
 sg13g2_buf_1 fanout9253 (.A(\soc_I.spi_div_ready ),
    .X(net9253));
 sg13g2_buf_4 fanout9254 (.X(net9254),
    .A(\soc_I.div_ready ));
 sg13g2_buf_2 fanout9255 (.A(net9257),
    .X(net9255));
 sg13g2_buf_2 fanout9256 (.A(net9257),
    .X(net9256));
 sg13g2_buf_2 fanout9257 (.A(\soc_I.qqspi_I.is_quad ),
    .X(net9257));
 sg13g2_buf_2 fanout9258 (.A(net9259),
    .X(net9258));
 sg13g2_buf_2 fanout9259 (.A(net9264),
    .X(net9259));
 sg13g2_buf_2 fanout9260 (.A(net9263),
    .X(net9260));
 sg13g2_buf_2 fanout9261 (.A(net9262),
    .X(net9261));
 sg13g2_buf_2 fanout9262 (.A(net9263),
    .X(net9262));
 sg13g2_buf_1 fanout9263 (.A(net9264),
    .X(net9263));
 sg13g2_buf_2 fanout9264 (.A(net9265),
    .X(net9264));
 sg13g2_buf_4 fanout9265 (.X(net9265),
    .A(\soc_I.qqspi_I.is_quad ));
 sg13g2_buf_2 fanout9266 (.A(net9267),
    .X(net9266));
 sg13g2_buf_2 fanout9267 (.A(net9268),
    .X(net9267));
 sg13g2_buf_2 fanout9268 (.A(net4817),
    .X(net9268));
 sg13g2_buf_2 fanout9269 (.A(net9271),
    .X(net9269));
 sg13g2_buf_2 fanout9270 (.A(net9271),
    .X(net9270));
 sg13g2_buf_2 fanout9271 (.A(\soc_I.qqspi_I.ready ),
    .X(net9271));
 sg13g2_buf_2 fanout9272 (.A(\soc_I.tx_uart_i.bit_idx[0] ),
    .X(net9272));
 sg13g2_buf_2 fanout9273 (.A(net5476),
    .X(net9273));
 sg13g2_buf_2 fanout9274 (.A(\soc_I.rx_uart_i.bit_idx[0] ),
    .X(net9274));
 sg13g2_buf_4 fanout9275 (.X(net9275),
    .A(net9276));
 sg13g2_buf_4 fanout9276 (.X(net9276),
    .A(net5528));
 sg13g2_buf_2 fanout9277 (.A(net9278),
    .X(net9277));
 sg13g2_buf_4 fanout9278 (.X(net9278),
    .A(net4681));
 sg13g2_buf_4 fanout9279 (.X(net9279),
    .A(net9281));
 sg13g2_buf_1 fanout9280 (.A(net9281),
    .X(net9280));
 sg13g2_buf_4 fanout9281 (.X(net9281),
    .A(net5352));
 sg13g2_buf_4 fanout9282 (.X(net9282),
    .A(\soc_I.rx_uart_i.fifo_i.din[4] ));
 sg13g2_buf_4 fanout9283 (.X(net9283),
    .A(\soc_I.rx_uart_i.fifo_i.din[4] ));
 sg13g2_buf_4 fanout9284 (.X(net9284),
    .A(net5493));
 sg13g2_buf_2 fanout9285 (.A(\soc_I.rx_uart_i.fifo_i.din[3] ),
    .X(net9285));
 sg13g2_buf_4 fanout9286 (.X(net9286),
    .A(net9287));
 sg13g2_buf_4 fanout9287 (.X(net9287),
    .A(net3981));
 sg13g2_buf_4 fanout9288 (.X(net9288),
    .A(net9289));
 sg13g2_buf_4 fanout9289 (.X(net9289),
    .A(\soc_I.rx_uart_i.fifo_i.din[1] ));
 sg13g2_buf_4 fanout9290 (.X(net9290),
    .A(net9293));
 sg13g2_buf_2 fanout9291 (.A(net9293),
    .X(net9291));
 sg13g2_buf_4 fanout9292 (.X(net9292),
    .A(net9293));
 sg13g2_buf_4 fanout9293 (.X(net9293),
    .A(\soc_I.clint_I.ready ));
 sg13g2_buf_2 fanout9294 (.A(net9295),
    .X(net9294));
 sg13g2_buf_2 fanout9295 (.A(net9296),
    .X(net9295));
 sg13g2_buf_4 fanout9296 (.X(net9296),
    .A(net9297));
 sg13g2_buf_8 fanout9297 (.A(net4985),
    .X(net9297));
 sg13g2_buf_4 fanout9298 (.X(net9298),
    .A(net9299));
 sg13g2_buf_4 fanout9299 (.X(net9299),
    .A(net9302));
 sg13g2_buf_4 fanout9300 (.X(net9300),
    .A(net9302));
 sg13g2_buf_2 fanout9301 (.A(net9302),
    .X(net9301));
 sg13g2_buf_2 fanout9302 (.A(net9336),
    .X(net9302));
 sg13g2_buf_2 fanout9303 (.A(net9304),
    .X(net9303));
 sg13g2_buf_2 fanout9304 (.A(net9305),
    .X(net9304));
 sg13g2_buf_2 fanout9305 (.A(net9306),
    .X(net9305));
 sg13g2_buf_2 fanout9306 (.A(net9336),
    .X(net9306));
 sg13g2_buf_2 fanout9307 (.A(net9309),
    .X(net9307));
 sg13g2_buf_2 fanout9308 (.A(net9314),
    .X(net9308));
 sg13g2_buf_1 fanout9309 (.A(net9314),
    .X(net9309));
 sg13g2_buf_2 fanout9310 (.A(net9311),
    .X(net9310));
 sg13g2_buf_2 fanout9311 (.A(net9314),
    .X(net9311));
 sg13g2_buf_2 fanout9312 (.A(net9313),
    .X(net9312));
 sg13g2_buf_4 fanout9313 (.X(net9313),
    .A(net9314));
 sg13g2_buf_2 fanout9314 (.A(net9336),
    .X(net9314));
 sg13g2_buf_4 fanout9315 (.X(net9315),
    .A(net9317));
 sg13g2_buf_1 fanout9316 (.A(net9317),
    .X(net9316));
 sg13g2_buf_2 fanout9317 (.A(net9336),
    .X(net9317));
 sg13g2_buf_2 fanout9318 (.A(net9319),
    .X(net9318));
 sg13g2_buf_4 fanout9319 (.X(net9319),
    .A(net9336));
 sg13g2_buf_2 fanout9320 (.A(net9322),
    .X(net9320));
 sg13g2_buf_1 fanout9321 (.A(net9322),
    .X(net9321));
 sg13g2_buf_4 fanout9322 (.X(net9322),
    .A(net9326));
 sg13g2_buf_4 fanout9323 (.X(net9323),
    .A(net9325));
 sg13g2_buf_2 fanout9324 (.A(net9325),
    .X(net9324));
 sg13g2_buf_2 fanout9325 (.A(net9326),
    .X(net9325));
 sg13g2_buf_4 fanout9326 (.X(net9326),
    .A(net9335));
 sg13g2_buf_4 fanout9327 (.X(net9327),
    .A(net9330));
 sg13g2_buf_4 fanout9328 (.X(net9328),
    .A(net9330));
 sg13g2_buf_1 fanout9329 (.A(net9330),
    .X(net9329));
 sg13g2_buf_2 fanout9330 (.A(net9335),
    .X(net9330));
 sg13g2_buf_2 fanout9331 (.A(net9332),
    .X(net9331));
 sg13g2_buf_2 fanout9332 (.A(net9333),
    .X(net9332));
 sg13g2_buf_2 fanout9333 (.A(net9335),
    .X(net9333));
 sg13g2_buf_4 fanout9334 (.X(net9334),
    .A(net9335));
 sg13g2_buf_2 fanout9335 (.A(net9336),
    .X(net9335));
 sg13g2_buf_8 fanout9336 (.A(net9420),
    .X(net9336));
 sg13g2_buf_4 fanout9337 (.X(net9337),
    .A(net9345));
 sg13g2_buf_2 fanout9338 (.A(net9345),
    .X(net9338));
 sg13g2_buf_4 fanout9339 (.X(net9339),
    .A(net9342));
 sg13g2_buf_2 fanout9340 (.A(net9341),
    .X(net9340));
 sg13g2_buf_2 fanout9341 (.A(net9342),
    .X(net9341));
 sg13g2_buf_4 fanout9342 (.X(net9342),
    .A(net9345));
 sg13g2_buf_4 fanout9343 (.X(net9343),
    .A(net9345));
 sg13g2_buf_4 fanout9344 (.X(net9344),
    .A(net9345));
 sg13g2_buf_2 fanout9345 (.A(net9420),
    .X(net9345));
 sg13g2_buf_4 fanout9346 (.X(net9346),
    .A(net9347));
 sg13g2_buf_2 fanout9347 (.A(net9353),
    .X(net9347));
 sg13g2_buf_4 fanout9348 (.X(net9348),
    .A(net9351));
 sg13g2_buf_4 fanout9349 (.X(net9349),
    .A(net9351));
 sg13g2_buf_2 fanout9350 (.A(net9351),
    .X(net9350));
 sg13g2_buf_2 fanout9351 (.A(net9353),
    .X(net9351));
 sg13g2_buf_2 fanout9352 (.A(net9353),
    .X(net9352));
 sg13g2_buf_2 fanout9353 (.A(net9369),
    .X(net9353));
 sg13g2_buf_4 fanout9354 (.X(net9354),
    .A(net9355));
 sg13g2_buf_4 fanout9355 (.X(net9355),
    .A(net9356));
 sg13g2_buf_4 fanout9356 (.X(net9356),
    .A(net9361));
 sg13g2_buf_4 fanout9357 (.X(net9357),
    .A(net9358));
 sg13g2_buf_2 fanout9358 (.A(net9361),
    .X(net9358));
 sg13g2_buf_4 fanout9359 (.X(net9359),
    .A(net9361));
 sg13g2_buf_2 fanout9360 (.A(net9361),
    .X(net9360));
 sg13g2_buf_2 fanout9361 (.A(net9369),
    .X(net9361));
 sg13g2_buf_4 fanout9362 (.X(net9362),
    .A(net9364));
 sg13g2_buf_4 fanout9363 (.X(net9363),
    .A(net9364));
 sg13g2_buf_4 fanout9364 (.X(net9364),
    .A(net9369));
 sg13g2_buf_4 fanout9365 (.X(net9365),
    .A(net9368));
 sg13g2_buf_4 fanout9366 (.X(net9366),
    .A(net9368));
 sg13g2_buf_1 fanout9367 (.A(net9368),
    .X(net9367));
 sg13g2_buf_2 fanout9368 (.A(net9369),
    .X(net9368));
 sg13g2_buf_2 fanout9369 (.A(net9420),
    .X(net9369));
 sg13g2_buf_4 fanout9370 (.X(net9370),
    .A(net9375));
 sg13g2_buf_1 fanout9371 (.A(net9375),
    .X(net9371));
 sg13g2_buf_4 fanout9372 (.X(net9372),
    .A(net9373));
 sg13g2_buf_4 fanout9373 (.X(net9373),
    .A(net9374));
 sg13g2_buf_4 fanout9374 (.X(net9374),
    .A(net9375));
 sg13g2_buf_2 fanout9375 (.A(net9380),
    .X(net9375));
 sg13g2_buf_4 fanout9376 (.X(net9376),
    .A(net9380));
 sg13g2_buf_2 fanout9377 (.A(net9380),
    .X(net9377));
 sg13g2_buf_4 fanout9378 (.X(net9378),
    .A(net9379));
 sg13g2_buf_2 fanout9379 (.A(net9380),
    .X(net9379));
 sg13g2_buf_2 fanout9380 (.A(net9407),
    .X(net9380));
 sg13g2_buf_4 fanout9381 (.X(net9381),
    .A(net9382));
 sg13g2_buf_4 fanout9382 (.X(net9382),
    .A(net9385));
 sg13g2_buf_4 fanout9383 (.X(net9383),
    .A(net9384));
 sg13g2_buf_4 fanout9384 (.X(net9384),
    .A(net9385));
 sg13g2_buf_2 fanout9385 (.A(net9391),
    .X(net9385));
 sg13g2_buf_4 fanout9386 (.X(net9386),
    .A(net9391));
 sg13g2_buf_4 fanout9387 (.X(net9387),
    .A(net9390));
 sg13g2_buf_2 fanout9388 (.A(net9390),
    .X(net9388));
 sg13g2_buf_4 fanout9389 (.X(net9389),
    .A(net9390));
 sg13g2_buf_2 fanout9390 (.A(net9391),
    .X(net9390));
 sg13g2_buf_4 fanout9391 (.X(net9391),
    .A(net9407));
 sg13g2_buf_4 fanout9392 (.X(net9392),
    .A(net9393));
 sg13g2_buf_2 fanout9393 (.A(net9394),
    .X(net9393));
 sg13g2_buf_2 fanout9394 (.A(net9395),
    .X(net9394));
 sg13g2_buf_2 fanout9395 (.A(net9396),
    .X(net9395));
 sg13g2_buf_4 fanout9396 (.X(net9396),
    .A(net9407));
 sg13g2_buf_4 fanout9397 (.X(net9397),
    .A(net9398));
 sg13g2_buf_4 fanout9398 (.X(net9398),
    .A(net9403));
 sg13g2_buf_4 fanout9399 (.X(net9399),
    .A(net9402));
 sg13g2_buf_2 fanout9400 (.A(net9402),
    .X(net9400));
 sg13g2_buf_4 fanout9401 (.X(net9401),
    .A(net9402));
 sg13g2_buf_2 fanout9402 (.A(net9403),
    .X(net9402));
 sg13g2_buf_2 fanout9403 (.A(net9407),
    .X(net9403));
 sg13g2_buf_4 fanout9404 (.X(net9404),
    .A(net9406));
 sg13g2_buf_2 fanout9405 (.A(net9406),
    .X(net9405));
 sg13g2_buf_4 fanout9406 (.X(net9406),
    .A(net9407));
 sg13g2_buf_8 fanout9407 (.A(net9419),
    .X(net9407));
 sg13g2_buf_2 fanout9408 (.A(net9409),
    .X(net9408));
 sg13g2_buf_2 fanout9409 (.A(net9413),
    .X(net9409));
 sg13g2_buf_4 fanout9410 (.X(net9410),
    .A(net9411));
 sg13g2_buf_4 fanout9411 (.X(net9411),
    .A(net9412));
 sg13g2_buf_2 fanout9412 (.A(net9413),
    .X(net9412));
 sg13g2_buf_4 fanout9413 (.X(net9413),
    .A(net9419));
 sg13g2_buf_2 fanout9414 (.A(net9415),
    .X(net9414));
 sg13g2_buf_1 fanout9415 (.A(net9416),
    .X(net9415));
 sg13g2_buf_4 fanout9416 (.X(net9416),
    .A(net9419));
 sg13g2_buf_2 fanout9417 (.A(net9418),
    .X(net9417));
 sg13g2_buf_4 fanout9418 (.X(net9418),
    .A(net9419));
 sg13g2_buf_8 fanout9419 (.A(net9420),
    .X(net9419));
 sg13g2_buf_8 fanout9420 (.A(\soc_I.clint_I.resetn ),
    .X(net9420));
 sg13g2_buf_2 fanout9421 (.A(\soc_I.kianv_I.datapath_unit_I.ADDR_I.q[1] ),
    .X(net9421));
 sg13g2_buf_2 fanout9422 (.A(\soc_I.kianv_I.datapath_unit_I.ADDR_I.q[1] ),
    .X(net9422));
 sg13g2_buf_2 fanout9423 (.A(net9424),
    .X(net9423));
 sg13g2_buf_2 fanout9424 (.A(net5503),
    .X(net9424));
 sg13g2_buf_2 fanout9425 (.A(net9426),
    .X(net9425));
 sg13g2_buf_2 fanout9426 (.A(net5487),
    .X(net9426));
 sg13g2_buf_4 fanout9427 (.X(net9427),
    .A(net9429));
 sg13g2_buf_1 fanout9428 (.A(net9429),
    .X(net9428));
 sg13g2_buf_2 fanout9429 (.A(\soc_I.kianv_I.Instr[29] ),
    .X(net9429));
 sg13g2_buf_4 fanout9430 (.X(net9430),
    .A(net5544));
 sg13g2_buf_4 fanout9431 (.X(net9431),
    .A(\soc_I.kianv_I.Instr[27] ));
 sg13g2_buf_4 fanout9432 (.X(net9432),
    .A(net9433));
 sg13g2_buf_2 fanout9433 (.A(net9435),
    .X(net9433));
 sg13g2_buf_8 fanout9434 (.A(net9435),
    .X(net9434));
 sg13g2_buf_8 fanout9435 (.A(\soc_I.kianv_I.Instr[24] ),
    .X(net9435));
 sg13g2_buf_4 fanout9436 (.X(net9436),
    .A(net9439));
 sg13g2_buf_4 fanout9437 (.X(net9437),
    .A(net9439));
 sg13g2_buf_8 fanout9438 (.A(net9439),
    .X(net9438));
 sg13g2_buf_8 fanout9439 (.A(\soc_I.kianv_I.Instr[24] ),
    .X(net9439));
 sg13g2_buf_4 fanout9440 (.X(net9440),
    .A(net9441));
 sg13g2_buf_4 fanout9441 (.X(net9441),
    .A(net9443));
 sg13g2_buf_8 fanout9442 (.A(net9443),
    .X(net9442));
 sg13g2_buf_8 fanout9443 (.A(\soc_I.kianv_I.Instr[23] ),
    .X(net9443));
 sg13g2_buf_8 fanout9444 (.A(net9450),
    .X(net9444));
 sg13g2_buf_4 fanout9445 (.X(net9445),
    .A(net9450));
 sg13g2_buf_4 fanout9446 (.X(net9446),
    .A(net9448));
 sg13g2_buf_4 fanout9447 (.X(net9447),
    .A(net9448));
 sg13g2_buf_2 fanout9448 (.A(net9450),
    .X(net9448));
 sg13g2_buf_4 fanout9449 (.X(net9449),
    .A(net9450));
 sg13g2_buf_8 fanout9450 (.A(\soc_I.kianv_I.Instr[23] ),
    .X(net9450));
 sg13g2_buf_4 fanout9451 (.X(net9451),
    .A(net9452));
 sg13g2_buf_2 fanout9452 (.A(net9454),
    .X(net9452));
 sg13g2_buf_4 fanout9453 (.X(net9453),
    .A(net9454));
 sg13g2_buf_2 fanout9454 (.A(net9461),
    .X(net9454));
 sg13g2_buf_4 fanout9455 (.X(net9455),
    .A(net9461));
 sg13g2_buf_2 fanout9456 (.A(net9461),
    .X(net9456));
 sg13g2_buf_4 fanout9457 (.X(net9457),
    .A(net9460));
 sg13g2_buf_4 fanout9458 (.X(net9458),
    .A(net9460));
 sg13g2_buf_2 fanout9459 (.A(net9460),
    .X(net9459));
 sg13g2_buf_2 fanout9460 (.A(net9461),
    .X(net9460));
 sg13g2_buf_4 fanout9461 (.X(net9461),
    .A(\soc_I.kianv_I.Instr[22] ));
 sg13g2_buf_4 fanout9462 (.X(net9462),
    .A(net9466));
 sg13g2_buf_2 fanout9463 (.A(net9466),
    .X(net9463));
 sg13g2_buf_2 fanout9464 (.A(net9466),
    .X(net9464));
 sg13g2_buf_2 fanout9465 (.A(net9466),
    .X(net9465));
 sg13g2_buf_2 fanout9466 (.A(\soc_I.kianv_I.Instr[22] ),
    .X(net9466));
 sg13g2_buf_4 fanout9467 (.X(net9467),
    .A(net9469));
 sg13g2_buf_4 fanout9468 (.X(net9468),
    .A(net9469));
 sg13g2_buf_4 fanout9469 (.X(net9469),
    .A(net9475));
 sg13g2_buf_4 fanout9470 (.X(net9470),
    .A(net9471));
 sg13g2_buf_4 fanout9471 (.X(net9471),
    .A(net9475));
 sg13g2_buf_4 fanout9472 (.X(net9472),
    .A(net9475));
 sg13g2_buf_2 fanout9473 (.A(net9474),
    .X(net9473));
 sg13g2_buf_4 fanout9474 (.X(net9474),
    .A(net9475));
 sg13g2_buf_4 fanout9475 (.X(net9475),
    .A(\soc_I.kianv_I.Instr[22] ));
 sg13g2_buf_4 fanout9476 (.X(net9476),
    .A(net9477));
 sg13g2_buf_4 fanout9477 (.X(net9477),
    .A(net9478));
 sg13g2_buf_2 fanout9478 (.A(net9484),
    .X(net9478));
 sg13g2_buf_4 fanout9479 (.X(net9479),
    .A(net9480));
 sg13g2_buf_4 fanout9480 (.X(net9480),
    .A(net9484));
 sg13g2_buf_4 fanout9481 (.X(net9481),
    .A(net9483));
 sg13g2_buf_2 fanout9482 (.A(net9483),
    .X(net9482));
 sg13g2_buf_4 fanout9483 (.X(net9483),
    .A(net9484));
 sg13g2_buf_8 fanout9484 (.A(\soc_I.kianv_I.Instr[21] ),
    .X(net9484));
 sg13g2_buf_4 fanout9485 (.X(net9485),
    .A(net9488));
 sg13g2_buf_4 fanout9486 (.X(net9486),
    .A(net9487));
 sg13g2_buf_4 fanout9487 (.X(net9487),
    .A(net9488));
 sg13g2_buf_8 fanout9488 (.A(\soc_I.kianv_I.Instr[21] ),
    .X(net9488));
 sg13g2_buf_4 fanout9489 (.X(net9489),
    .A(net9491));
 sg13g2_buf_4 fanout9490 (.X(net9490),
    .A(net9491));
 sg13g2_buf_4 fanout9491 (.X(net9491),
    .A(net9509));
 sg13g2_buf_4 fanout9492 (.X(net9492),
    .A(net9495));
 sg13g2_buf_4 fanout9493 (.X(net9493),
    .A(net9494));
 sg13g2_buf_2 fanout9494 (.A(net9495),
    .X(net9494));
 sg13g2_buf_2 fanout9495 (.A(net9509),
    .X(net9495));
 sg13g2_buf_4 fanout9496 (.X(net9496),
    .A(net9497));
 sg13g2_buf_4 fanout9497 (.X(net9497),
    .A(net9500));
 sg13g2_buf_4 fanout9498 (.X(net9498),
    .A(net9500));
 sg13g2_buf_4 fanout9499 (.X(net9499),
    .A(net9500));
 sg13g2_buf_2 fanout9500 (.A(net9509),
    .X(net9500));
 sg13g2_buf_4 fanout9501 (.X(net9501),
    .A(net9504));
 sg13g2_buf_4 fanout9502 (.X(net9502),
    .A(net9504));
 sg13g2_buf_2 fanout9503 (.A(net9504),
    .X(net9503));
 sg13g2_buf_2 fanout9504 (.A(net9509),
    .X(net9504));
 sg13g2_buf_4 fanout9505 (.X(net9505),
    .A(net9508));
 sg13g2_buf_2 fanout9506 (.A(net9508),
    .X(net9506));
 sg13g2_buf_4 fanout9507 (.X(net9507),
    .A(net9508));
 sg13g2_buf_2 fanout9508 (.A(net9509),
    .X(net9508));
 sg13g2_buf_8 fanout9509 (.A(\soc_I.kianv_I.Instr[21] ),
    .X(net9509));
 sg13g2_buf_4 fanout9510 (.X(net9510),
    .A(net9511));
 sg13g2_buf_4 fanout9511 (.X(net9511),
    .A(net9512));
 sg13g2_buf_2 fanout9512 (.A(net9524),
    .X(net9512));
 sg13g2_buf_4 fanout9513 (.X(net9513),
    .A(net9514));
 sg13g2_buf_4 fanout9514 (.X(net9514),
    .A(net9524));
 sg13g2_buf_4 fanout9515 (.X(net9515),
    .A(net9518));
 sg13g2_buf_2 fanout9516 (.A(net9518),
    .X(net9516));
 sg13g2_buf_4 fanout9517 (.X(net9517),
    .A(net9518));
 sg13g2_buf_2 fanout9518 (.A(net9524),
    .X(net9518));
 sg13g2_buf_4 fanout9519 (.X(net9519),
    .A(net9520));
 sg13g2_buf_4 fanout9520 (.X(net9520),
    .A(net9523));
 sg13g2_buf_4 fanout9521 (.X(net9521),
    .A(net9522));
 sg13g2_buf_8 fanout9522 (.A(net9523),
    .X(net9522));
 sg13g2_buf_4 fanout9523 (.X(net9523),
    .A(net9524));
 sg13g2_buf_8 fanout9524 (.A(\soc_I.kianv_I.Instr[20] ),
    .X(net9524));
 sg13g2_buf_4 fanout9525 (.X(net9525),
    .A(net9526));
 sg13g2_buf_2 fanout9526 (.A(net9531),
    .X(net9526));
 sg13g2_buf_4 fanout9527 (.X(net9527),
    .A(net9531));
 sg13g2_buf_4 fanout9528 (.X(net9528),
    .A(net9530));
 sg13g2_buf_1 fanout9529 (.A(net9530),
    .X(net9529));
 sg13g2_buf_4 fanout9530 (.X(net9530),
    .A(net9531));
 sg13g2_buf_2 fanout9531 (.A(net9545),
    .X(net9531));
 sg13g2_buf_4 fanout9532 (.X(net9532),
    .A(net9534));
 sg13g2_buf_2 fanout9533 (.A(net9534),
    .X(net9533));
 sg13g2_buf_2 fanout9534 (.A(net9545),
    .X(net9534));
 sg13g2_buf_4 fanout9535 (.X(net9535),
    .A(net9536));
 sg13g2_buf_4 fanout9536 (.X(net9536),
    .A(net9545));
 sg13g2_buf_4 fanout9537 (.X(net9537),
    .A(net9544));
 sg13g2_buf_4 fanout9538 (.X(net9538),
    .A(net9539));
 sg13g2_buf_4 fanout9539 (.X(net9539),
    .A(net9544));
 sg13g2_buf_4 fanout9540 (.X(net9540),
    .A(net9543));
 sg13g2_buf_2 fanout9541 (.A(net9543),
    .X(net9541));
 sg13g2_buf_4 fanout9542 (.X(net9542),
    .A(net9543));
 sg13g2_buf_4 fanout9543 (.X(net9543),
    .A(net9544));
 sg13g2_buf_2 fanout9544 (.A(net9545),
    .X(net9544));
 sg13g2_buf_8 fanout9545 (.A(\soc_I.kianv_I.Instr[20] ),
    .X(net9545));
 sg13g2_buf_8 fanout9546 (.A(net9547),
    .X(net9546));
 sg13g2_buf_8 fanout9547 (.A(net9552),
    .X(net9547));
 sg13g2_buf_4 fanout9548 (.X(net9548),
    .A(net9552));
 sg13g2_buf_2 fanout9549 (.A(net9552),
    .X(net9549));
 sg13g2_buf_8 fanout9550 (.A(net9551),
    .X(net9550));
 sg13g2_buf_8 fanout9551 (.A(net9552),
    .X(net9551));
 sg13g2_buf_8 fanout9552 (.A(net5460),
    .X(net9552));
 sg13g2_buf_4 fanout9553 (.X(net9553),
    .A(net9554));
 sg13g2_buf_8 fanout9554 (.A(net9556),
    .X(net9554));
 sg13g2_buf_8 fanout9555 (.A(net9556),
    .X(net9555));
 sg13g2_buf_8 fanout9556 (.A(net9563),
    .X(net9556));
 sg13g2_buf_4 fanout9557 (.X(net9557),
    .A(net9563));
 sg13g2_buf_2 fanout9558 (.A(net9563),
    .X(net9558));
 sg13g2_buf_4 fanout9559 (.X(net9559),
    .A(net9562));
 sg13g2_buf_4 fanout9560 (.X(net9560),
    .A(net9561));
 sg13g2_buf_4 fanout9561 (.X(net9561),
    .A(net9562));
 sg13g2_buf_4 fanout9562 (.X(net9562),
    .A(net9563));
 sg13g2_buf_8 fanout9563 (.A(\soc_I.kianv_I.Instr[18] ),
    .X(net9563));
 sg13g2_buf_4 fanout9564 (.X(net9564),
    .A(net9566));
 sg13g2_buf_4 fanout9565 (.X(net9565),
    .A(net9566));
 sg13g2_buf_4 fanout9566 (.X(net9566),
    .A(net9570));
 sg13g2_buf_4 fanout9567 (.X(net9567),
    .A(net9570));
 sg13g2_buf_4 fanout9568 (.X(net9568),
    .A(net9570));
 sg13g2_buf_4 fanout9569 (.X(net9569),
    .A(net9570));
 sg13g2_buf_8 fanout9570 (.A(\soc_I.kianv_I.Instr[17] ),
    .X(net9570));
 sg13g2_buf_4 fanout9571 (.X(net9571),
    .A(net9574));
 sg13g2_buf_4 fanout9572 (.X(net9572),
    .A(net9574));
 sg13g2_buf_2 fanout9573 (.A(net9574),
    .X(net9573));
 sg13g2_buf_4 fanout9574 (.X(net9574),
    .A(net9582));
 sg13g2_buf_4 fanout9575 (.X(net9575),
    .A(net9582));
 sg13g2_buf_2 fanout9576 (.A(net9582),
    .X(net9576));
 sg13g2_buf_4 fanout9577 (.X(net9577),
    .A(net9581));
 sg13g2_buf_4 fanout9578 (.X(net9578),
    .A(net9581));
 sg13g2_buf_2 fanout9579 (.A(net9580),
    .X(net9579));
 sg13g2_buf_4 fanout9580 (.X(net9580),
    .A(net9581));
 sg13g2_buf_4 fanout9581 (.X(net9581),
    .A(net9582));
 sg13g2_buf_8 fanout9582 (.A(\soc_I.kianv_I.Instr[17] ),
    .X(net9582));
 sg13g2_buf_4 fanout9583 (.X(net9583),
    .A(net9586));
 sg13g2_buf_2 fanout9584 (.A(net9586),
    .X(net9584));
 sg13g2_buf_4 fanout9585 (.X(net9585),
    .A(net9586));
 sg13g2_buf_2 fanout9586 (.A(net9587),
    .X(net9586));
 sg13g2_buf_2 fanout9587 (.A(net9607),
    .X(net9587));
 sg13g2_buf_4 fanout9588 (.X(net9588),
    .A(net9590));
 sg13g2_buf_2 fanout9589 (.A(net9590),
    .X(net9589));
 sg13g2_buf_4 fanout9590 (.X(net9590),
    .A(net9607));
 sg13g2_buf_4 fanout9591 (.X(net9591),
    .A(net9593));
 sg13g2_buf_4 fanout9592 (.X(net9592),
    .A(net9593));
 sg13g2_buf_4 fanout9593 (.X(net9593),
    .A(net9596));
 sg13g2_buf_4 fanout9594 (.X(net9594),
    .A(net9596));
 sg13g2_buf_2 fanout9595 (.A(net9596),
    .X(net9595));
 sg13g2_buf_2 fanout9596 (.A(net9607),
    .X(net9596));
 sg13g2_buf_4 fanout9597 (.X(net9597),
    .A(net9601));
 sg13g2_buf_2 fanout9598 (.A(net9601),
    .X(net9598));
 sg13g2_buf_4 fanout9599 (.X(net9599),
    .A(net9601));
 sg13g2_buf_2 fanout9600 (.A(net9601),
    .X(net9600));
 sg13g2_buf_2 fanout9601 (.A(net9607),
    .X(net9601));
 sg13g2_buf_4 fanout9602 (.X(net9602),
    .A(net9606));
 sg13g2_buf_2 fanout9603 (.A(net9606),
    .X(net9603));
 sg13g2_buf_4 fanout9604 (.X(net9604),
    .A(net9605));
 sg13g2_buf_2 fanout9605 (.A(net9606),
    .X(net9605));
 sg13g2_buf_4 fanout9606 (.X(net9606),
    .A(net9607));
 sg13g2_buf_8 fanout9607 (.A(\soc_I.kianv_I.Instr[16] ),
    .X(net9607));
 sg13g2_buf_4 fanout9608 (.X(net9608),
    .A(net9612));
 sg13g2_buf_2 fanout9609 (.A(net9612),
    .X(net9609));
 sg13g2_buf_4 fanout9610 (.X(net9610),
    .A(net9611));
 sg13g2_buf_4 fanout9611 (.X(net9611),
    .A(net9612));
 sg13g2_buf_2 fanout9612 (.A(net9641),
    .X(net9612));
 sg13g2_buf_4 fanout9613 (.X(net9613),
    .A(net9615));
 sg13g2_buf_4 fanout9614 (.X(net9614),
    .A(net9615));
 sg13g2_buf_2 fanout9615 (.A(net9641),
    .X(net9615));
 sg13g2_buf_4 fanout9616 (.X(net9616),
    .A(net9618));
 sg13g2_buf_2 fanout9617 (.A(net9618),
    .X(net9617));
 sg13g2_buf_2 fanout9618 (.A(net9641),
    .X(net9618));
 sg13g2_buf_4 fanout9619 (.X(net9619),
    .A(net9621));
 sg13g2_buf_2 fanout9620 (.A(net9621),
    .X(net9620));
 sg13g2_buf_2 fanout9621 (.A(net9622),
    .X(net9621));
 sg13g2_buf_2 fanout9622 (.A(net9640),
    .X(net9622));
 sg13g2_buf_4 fanout9623 (.X(net9623),
    .A(net9624));
 sg13g2_buf_4 fanout9624 (.X(net9624),
    .A(net9640));
 sg13g2_buf_4 fanout9625 (.X(net9625),
    .A(net9627));
 sg13g2_buf_4 fanout9626 (.X(net9626),
    .A(net9627));
 sg13g2_buf_2 fanout9627 (.A(net9640),
    .X(net9627));
 sg13g2_buf_4 fanout9628 (.X(net9628),
    .A(net9632));
 sg13g2_buf_4 fanout9629 (.X(net9629),
    .A(net9632));
 sg13g2_buf_4 fanout9630 (.X(net9630),
    .A(net9631));
 sg13g2_buf_4 fanout9631 (.X(net9631),
    .A(net9632));
 sg13g2_buf_2 fanout9632 (.A(net9640),
    .X(net9632));
 sg13g2_buf_4 fanout9633 (.X(net9633),
    .A(net9635));
 sg13g2_buf_4 fanout9634 (.X(net9634),
    .A(net9635));
 sg13g2_buf_2 fanout9635 (.A(net9639),
    .X(net9635));
 sg13g2_buf_4 fanout9636 (.X(net9636),
    .A(net9639));
 sg13g2_buf_2 fanout9637 (.A(net9639),
    .X(net9637));
 sg13g2_buf_4 fanout9638 (.X(net9638),
    .A(net9639));
 sg13g2_buf_2 fanout9639 (.A(net9640),
    .X(net9639));
 sg13g2_buf_4 fanout9640 (.X(net9640),
    .A(net9641));
 sg13g2_buf_4 fanout9641 (.X(net9641),
    .A(\soc_I.kianv_I.Instr[16] ));
 sg13g2_buf_8 fanout9642 (.A(net9645),
    .X(net9642));
 sg13g2_buf_4 fanout9643 (.X(net9643),
    .A(net9645));
 sg13g2_buf_4 fanout9644 (.X(net9644),
    .A(net9645));
 sg13g2_buf_2 fanout9645 (.A(net9646),
    .X(net9645));
 sg13g2_buf_2 fanout9646 (.A(net9664),
    .X(net9646));
 sg13g2_buf_8 fanout9647 (.A(net9649),
    .X(net9647));
 sg13g2_buf_4 fanout9648 (.X(net9648),
    .A(net9649));
 sg13g2_buf_4 fanout9649 (.X(net9649),
    .A(net9664));
 sg13g2_buf_4 fanout9650 (.X(net9650),
    .A(net9652));
 sg13g2_buf_4 fanout9651 (.X(net9651),
    .A(net9652));
 sg13g2_buf_4 fanout9652 (.X(net9652),
    .A(net9655));
 sg13g2_buf_4 fanout9653 (.X(net9653),
    .A(net9654));
 sg13g2_buf_2 fanout9654 (.A(net9655),
    .X(net9654));
 sg13g2_buf_2 fanout9655 (.A(net9664),
    .X(net9655));
 sg13g2_buf_4 fanout9656 (.X(net9656),
    .A(net9659));
 sg13g2_buf_4 fanout9657 (.X(net9657),
    .A(net9659));
 sg13g2_buf_2 fanout9658 (.A(net9659),
    .X(net9658));
 sg13g2_buf_4 fanout9659 (.X(net9659),
    .A(net9664));
 sg13g2_buf_8 fanout9660 (.A(net9663),
    .X(net9660));
 sg13g2_buf_4 fanout9661 (.X(net9661),
    .A(net9663));
 sg13g2_buf_8 fanout9662 (.A(net9663),
    .X(net9662));
 sg13g2_buf_4 fanout9663 (.X(net9663),
    .A(net9664));
 sg13g2_buf_4 fanout9664 (.X(net9664),
    .A(\soc_I.kianv_I.Instr[15] ));
 sg13g2_buf_4 fanout9665 (.X(net9665),
    .A(net9666));
 sg13g2_buf_4 fanout9666 (.X(net9666),
    .A(net9669));
 sg13g2_buf_4 fanout9667 (.X(net9667),
    .A(net9668));
 sg13g2_buf_4 fanout9668 (.X(net9668),
    .A(net9669));
 sg13g2_buf_2 fanout9669 (.A(net9697),
    .X(net9669));
 sg13g2_buf_8 fanout9670 (.A(net9672),
    .X(net9670));
 sg13g2_buf_4 fanout9671 (.X(net9671),
    .A(net9672));
 sg13g2_buf_4 fanout9672 (.X(net9672),
    .A(net9697));
 sg13g2_buf_8 fanout9673 (.A(net9675),
    .X(net9673));
 sg13g2_buf_4 fanout9674 (.X(net9674),
    .A(net9675));
 sg13g2_buf_2 fanout9675 (.A(net9697),
    .X(net9675));
 sg13g2_buf_4 fanout9676 (.X(net9676),
    .A(net9677));
 sg13g2_buf_4 fanout9677 (.X(net9677),
    .A(net9678));
 sg13g2_buf_4 fanout9678 (.X(net9678),
    .A(net9683));
 sg13g2_buf_4 fanout9679 (.X(net9679),
    .A(net9683));
 sg13g2_buf_4 fanout9680 (.X(net9680),
    .A(net9683));
 sg13g2_buf_8 fanout9681 (.A(net9682),
    .X(net9681));
 sg13g2_buf_4 fanout9682 (.X(net9682),
    .A(net9683));
 sg13g2_buf_2 fanout9683 (.A(net9697),
    .X(net9683));
 sg13g2_buf_8 fanout9684 (.A(net9685),
    .X(net9684));
 sg13g2_buf_4 fanout9685 (.X(net9685),
    .A(net9696));
 sg13g2_buf_8 fanout9686 (.A(net9696),
    .X(net9686));
 sg13g2_buf_8 fanout9687 (.A(net9696),
    .X(net9687));
 sg13g2_buf_4 fanout9688 (.X(net9688),
    .A(net9695));
 sg13g2_buf_2 fanout9689 (.A(net9695),
    .X(net9689));
 sg13g2_buf_4 fanout9690 (.X(net9690),
    .A(net9695));
 sg13g2_buf_4 fanout9691 (.X(net9691),
    .A(net9694));
 sg13g2_buf_8 fanout9692 (.A(net9694),
    .X(net9692));
 sg13g2_buf_4 fanout9693 (.X(net9693),
    .A(net9694));
 sg13g2_buf_2 fanout9694 (.A(net9695),
    .X(net9694));
 sg13g2_buf_2 fanout9695 (.A(net9696),
    .X(net9695));
 sg13g2_buf_4 fanout9696 (.X(net9696),
    .A(net9697));
 sg13g2_buf_8 fanout9697 (.A(\soc_I.kianv_I.Instr[15] ),
    .X(net9697));
 sg13g2_buf_4 fanout9698 (.X(net9698),
    .A(net9699));
 sg13g2_buf_4 fanout9699 (.X(net9699),
    .A(net5526));
 sg13g2_buf_4 fanout9700 (.X(net9700),
    .A(net5548));
 sg13g2_buf_4 fanout9701 (.X(net9701),
    .A(\soc_I.kianv_I.Instr[13] ));
 sg13g2_buf_4 fanout9702 (.X(net9702),
    .A(net9704));
 sg13g2_buf_4 fanout9703 (.X(net9703),
    .A(net9704));
 sg13g2_buf_2 fanout9704 (.A(net9705),
    .X(net9704));
 sg13g2_buf_4 fanout9705 (.X(net9705),
    .A(\soc_I.kianv_I.Instr[13] ));
 sg13g2_buf_4 fanout9706 (.X(net9706),
    .A(net9708));
 sg13g2_buf_4 fanout9707 (.X(net9707),
    .A(net5564));
 sg13g2_buf_2 fanout9708 (.A(\soc_I.kianv_I.Instr[12] ),
    .X(net9708));
 sg13g2_buf_4 fanout9709 (.X(net9709),
    .A(net5559));
 sg13g2_buf_2 fanout9710 (.A(net9711),
    .X(net9710));
 sg13g2_buf_2 fanout9711 (.A(\soc_I.kianv_I.Instr[10] ),
    .X(net9711));
 sg13g2_buf_4 fanout9712 (.X(net9712),
    .A(net5523));
 sg13g2_buf_2 fanout9713 (.A(net9714),
    .X(net9713));
 sg13g2_buf_1 fanout9714 (.A(net5491),
    .X(net9714));
 sg13g2_buf_2 fanout9715 (.A(net5494),
    .X(net9715));
 sg13g2_buf_2 fanout9716 (.A(net9717),
    .X(net9716));
 sg13g2_buf_2 fanout9717 (.A(net9718),
    .X(net9717));
 sg13g2_buf_1 fanout9718 (.A(net3890),
    .X(net9718));
 sg13g2_buf_4 fanout9719 (.X(net9719),
    .A(net9723));
 sg13g2_buf_2 fanout9720 (.A(net9721),
    .X(net9720));
 sg13g2_buf_2 fanout9721 (.A(net9722),
    .X(net9721));
 sg13g2_buf_2 fanout9722 (.A(net9723),
    .X(net9722));
 sg13g2_buf_2 fanout9723 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.bit_idx[4] ),
    .X(net9723));
 sg13g2_buf_2 fanout9724 (.A(net9726),
    .X(net9724));
 sg13g2_buf_1 fanout9725 (.A(net9726),
    .X(net9725));
 sg13g2_buf_2 fanout9726 (.A(net9730),
    .X(net9726));
 sg13g2_buf_2 fanout9727 (.A(net9728),
    .X(net9727));
 sg13g2_buf_2 fanout9728 (.A(net9729),
    .X(net9728));
 sg13g2_buf_2 fanout9729 (.A(net9730),
    .X(net9729));
 sg13g2_buf_2 fanout9730 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.bit_idx[4] ),
    .X(net9730));
 sg13g2_buf_4 fanout9731 (.X(net9731),
    .A(net9732));
 sg13g2_buf_2 fanout9732 (.A(_00254_),
    .X(net9732));
 sg13g2_buf_2 fanout9733 (.A(net9734),
    .X(net9733));
 sg13g2_buf_2 fanout9734 (.A(net9740),
    .X(net9734));
 sg13g2_buf_2 fanout9735 (.A(net9739),
    .X(net9735));
 sg13g2_buf_1 fanout9736 (.A(net9739),
    .X(net9736));
 sg13g2_buf_2 fanout9737 (.A(net9738),
    .X(net9737));
 sg13g2_buf_2 fanout9738 (.A(net9739),
    .X(net9738));
 sg13g2_buf_2 fanout9739 (.A(net9740),
    .X(net9739));
 sg13g2_buf_4 fanout9740 (.X(net9740),
    .A(net5469));
 sg13g2_buf_2 fanout9741 (.A(net9743),
    .X(net9741));
 sg13g2_buf_2 fanout9742 (.A(net9743),
    .X(net9742));
 sg13g2_buf_2 fanout9743 (.A(net9744),
    .X(net9743));
 sg13g2_buf_1 fanout9744 (.A(net5518),
    .X(net9744));
 sg13g2_buf_2 fanout9745 (.A(net9747),
    .X(net9745));
 sg13g2_buf_1 fanout9746 (.A(net9747),
    .X(net9746));
 sg13g2_buf_2 fanout9747 (.A(net9748),
    .X(net9747));
 sg13g2_buf_2 fanout9748 (.A(net9749),
    .X(net9748));
 sg13g2_buf_1 fanout9749 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.bit_idx[2] ),
    .X(net9749));
 sg13g2_buf_2 fanout9750 (.A(net9752),
    .X(net9750));
 sg13g2_buf_2 fanout9751 (.A(net9752),
    .X(net9751));
 sg13g2_buf_2 fanout9752 (.A(net9757),
    .X(net9752));
 sg13g2_buf_2 fanout9753 (.A(net9756),
    .X(net9753));
 sg13g2_buf_2 fanout9754 (.A(net9755),
    .X(net9754));
 sg13g2_buf_2 fanout9755 (.A(net9756),
    .X(net9755));
 sg13g2_buf_1 fanout9756 (.A(net9757),
    .X(net9756));
 sg13g2_buf_2 fanout9757 (.A(net9758),
    .X(net9757));
 sg13g2_buf_4 fanout9758 (.X(net9758),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.bit_idx[1] ));
 sg13g2_buf_2 fanout9759 (.A(net9763),
    .X(net9759));
 sg13g2_buf_1 fanout9760 (.A(net9763),
    .X(net9760));
 sg13g2_buf_2 fanout9761 (.A(net9762),
    .X(net9761));
 sg13g2_buf_2 fanout9762 (.A(net9763),
    .X(net9762));
 sg13g2_buf_1 fanout9763 (.A(net9768),
    .X(net9763));
 sg13g2_buf_2 fanout9764 (.A(net9766),
    .X(net9764));
 sg13g2_buf_2 fanout9765 (.A(net9766),
    .X(net9765));
 sg13g2_buf_2 fanout9766 (.A(net9767),
    .X(net9766));
 sg13g2_buf_4 fanout9767 (.X(net9767),
    .A(net9768));
 sg13g2_buf_4 fanout9768 (.X(net9768),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.bit_idx[0] ));
 sg13g2_buf_4 fanout9769 (.X(net9769),
    .A(\soc_I.kianv_I.datapath_unit_I.mul_I.bit_idx[0] ));
 sg13g2_buf_2 fanout9770 (.A(net9771),
    .X(net9770));
 sg13g2_buf_4 fanout9771 (.X(net9771),
    .A(net9780));
 sg13g2_buf_4 fanout9772 (.X(net9772),
    .A(net9774));
 sg13g2_buf_2 fanout9773 (.A(net9774),
    .X(net9773));
 sg13g2_buf_2 fanout9774 (.A(net9780),
    .X(net9774));
 sg13g2_buf_2 fanout9775 (.A(net9776),
    .X(net9775));
 sg13g2_buf_2 fanout9776 (.A(net9780),
    .X(net9776));
 sg13g2_buf_2 fanout9777 (.A(net9779),
    .X(net9777));
 sg13g2_buf_1 fanout9778 (.A(net9779),
    .X(net9778));
 sg13g2_buf_4 fanout9779 (.X(net9779),
    .A(net9780));
 sg13g2_buf_4 fanout9780 (.X(net9780),
    .A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_select ));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_4 input5 (.X(net5),
    .A(ui_in[3]));
 sg13g2_buf_2 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_buf_2 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_4 input11 (.X(net11),
    .A(uio_in[2]));
 sg13g2_buf_2 input12 (.A(uio_in[4]),
    .X(net12));
 sg13g2_buf_2 input13 (.A(uio_in[5]),
    .X(net13));
 sg13g2_tiehi _35931__14 (.L_HI(net14));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_leaf_49_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_2 clkbuf_leaf_50_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_2 clkbuf_leaf_51_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_2 clkbuf_leaf_52_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_2 clkbuf_leaf_53_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_2 clkbuf_leaf_54_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_2 clkbuf_leaf_55_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_2 clkbuf_leaf_56_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_2 clkbuf_leaf_57_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_2 clkbuf_leaf_58_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_2 clkbuf_leaf_59_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_2 clkbuf_leaf_60_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_2 clkbuf_leaf_61_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_2 clkbuf_leaf_62_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_2 clkbuf_leaf_63_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_2 clkbuf_leaf_64_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_2 clkbuf_leaf_65_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_2 clkbuf_leaf_66_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_2 clkbuf_leaf_67_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_2 clkbuf_leaf_68_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_2 clkbuf_leaf_69_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_2 clkbuf_leaf_70_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_2 clkbuf_leaf_71_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_2 clkbuf_leaf_72_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_2 clkbuf_leaf_73_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_2 clkbuf_leaf_74_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_2 clkbuf_leaf_75_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_2 clkbuf_leaf_76_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_2 clkbuf_leaf_77_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_2 clkbuf_leaf_78_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_2 clkbuf_leaf_79_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_2 clkbuf_leaf_80_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_2 clkbuf_leaf_81_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_2 clkbuf_leaf_82_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_2 clkbuf_leaf_83_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_2 clkbuf_leaf_84_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_2 clkbuf_leaf_85_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_2 clkbuf_leaf_86_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_2 clkbuf_leaf_87_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_2 clkbuf_leaf_88_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_2 clkbuf_leaf_89_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_2 clkbuf_leaf_90_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_2 clkbuf_leaf_91_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_2 clkbuf_leaf_92_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_2 clkbuf_leaf_93_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_2 clkbuf_leaf_94_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_2 clkbuf_leaf_95_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_2 clkbuf_leaf_96_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_2 clkbuf_leaf_97_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_2 clkbuf_leaf_98_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_2 clkbuf_leaf_99_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_2 clkbuf_leaf_100_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_2 clkbuf_leaf_101_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_2 clkbuf_leaf_102_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_2 clkbuf_leaf_103_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_2 clkbuf_leaf_104_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_2 clkbuf_leaf_105_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_2 clkbuf_leaf_106_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_2 clkbuf_leaf_107_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_2 clkbuf_leaf_108_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_2 clkbuf_leaf_109_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_2 clkbuf_leaf_110_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_110_clk));
 sg13g2_buf_2 clkbuf_leaf_111_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_111_clk));
 sg13g2_buf_2 clkbuf_leaf_112_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_112_clk));
 sg13g2_buf_2 clkbuf_leaf_113_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_113_clk));
 sg13g2_buf_2 clkbuf_leaf_114_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_114_clk));
 sg13g2_buf_2 clkbuf_leaf_115_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_115_clk));
 sg13g2_buf_2 clkbuf_leaf_116_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_116_clk));
 sg13g2_buf_2 clkbuf_leaf_117_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_117_clk));
 sg13g2_buf_2 clkbuf_leaf_118_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_118_clk));
 sg13g2_buf_2 clkbuf_leaf_119_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_119_clk));
 sg13g2_buf_2 clkbuf_leaf_120_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_120_clk));
 sg13g2_buf_2 clkbuf_leaf_121_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_121_clk));
 sg13g2_buf_2 clkbuf_leaf_122_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_122_clk));
 sg13g2_buf_2 clkbuf_leaf_123_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_123_clk));
 sg13g2_buf_2 clkbuf_leaf_124_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_124_clk));
 sg13g2_buf_2 clkbuf_leaf_125_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_125_clk));
 sg13g2_buf_2 clkbuf_leaf_126_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_126_clk));
 sg13g2_buf_2 clkbuf_leaf_127_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_127_clk));
 sg13g2_buf_2 clkbuf_leaf_128_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_128_clk));
 sg13g2_buf_2 clkbuf_leaf_129_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_129_clk));
 sg13g2_buf_2 clkbuf_leaf_130_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_130_clk));
 sg13g2_buf_2 clkbuf_leaf_131_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_131_clk));
 sg13g2_buf_2 clkbuf_leaf_132_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_132_clk));
 sg13g2_buf_2 clkbuf_leaf_133_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_133_clk));
 sg13g2_buf_2 clkbuf_leaf_134_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_134_clk));
 sg13g2_buf_2 clkbuf_leaf_135_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_135_clk));
 sg13g2_buf_2 clkbuf_leaf_136_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_136_clk));
 sg13g2_buf_2 clkbuf_leaf_137_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_137_clk));
 sg13g2_buf_2 clkbuf_leaf_138_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_138_clk));
 sg13g2_buf_2 clkbuf_leaf_139_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_139_clk));
 sg13g2_buf_2 clkbuf_leaf_140_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_140_clk));
 sg13g2_buf_2 clkbuf_leaf_141_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_141_clk));
 sg13g2_buf_2 clkbuf_leaf_142_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_142_clk));
 sg13g2_buf_2 clkbuf_leaf_143_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_143_clk));
 sg13g2_buf_2 clkbuf_leaf_144_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_144_clk));
 sg13g2_buf_2 clkbuf_leaf_145_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_145_clk));
 sg13g2_buf_2 clkbuf_leaf_146_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_146_clk));
 sg13g2_buf_2 clkbuf_leaf_147_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_147_clk));
 sg13g2_buf_2 clkbuf_leaf_148_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_148_clk));
 sg13g2_buf_2 clkbuf_leaf_149_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_149_clk));
 sg13g2_buf_2 clkbuf_leaf_150_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_150_clk));
 sg13g2_buf_2 clkbuf_leaf_151_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_151_clk));
 sg13g2_buf_2 clkbuf_leaf_152_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_152_clk));
 sg13g2_buf_2 clkbuf_leaf_153_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_153_clk));
 sg13g2_buf_2 clkbuf_leaf_154_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_154_clk));
 sg13g2_buf_2 clkbuf_leaf_155_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_155_clk));
 sg13g2_buf_2 clkbuf_leaf_156_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_156_clk));
 sg13g2_buf_2 clkbuf_leaf_157_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_157_clk));
 sg13g2_buf_2 clkbuf_leaf_158_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_158_clk));
 sg13g2_buf_2 clkbuf_leaf_159_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_159_clk));
 sg13g2_buf_2 clkbuf_leaf_160_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_160_clk));
 sg13g2_buf_2 clkbuf_leaf_161_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_161_clk));
 sg13g2_buf_2 clkbuf_leaf_162_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_162_clk));
 sg13g2_buf_2 clkbuf_leaf_163_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_163_clk));
 sg13g2_buf_2 clkbuf_leaf_164_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_164_clk));
 sg13g2_buf_2 clkbuf_leaf_165_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_165_clk));
 sg13g2_buf_2 clkbuf_leaf_166_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_166_clk));
 sg13g2_buf_2 clkbuf_leaf_167_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_167_clk));
 sg13g2_buf_2 clkbuf_leaf_168_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_168_clk));
 sg13g2_buf_2 clkbuf_leaf_169_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_169_clk));
 sg13g2_buf_2 clkbuf_leaf_170_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_170_clk));
 sg13g2_buf_2 clkbuf_leaf_171_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_171_clk));
 sg13g2_buf_2 clkbuf_leaf_172_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_172_clk));
 sg13g2_buf_2 clkbuf_leaf_173_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_173_clk));
 sg13g2_buf_2 clkbuf_leaf_174_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_174_clk));
 sg13g2_buf_2 clkbuf_leaf_175_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_175_clk));
 sg13g2_buf_2 clkbuf_leaf_176_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_176_clk));
 sg13g2_buf_2 clkbuf_leaf_177_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_177_clk));
 sg13g2_buf_2 clkbuf_leaf_178_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_178_clk));
 sg13g2_buf_2 clkbuf_leaf_179_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_179_clk));
 sg13g2_buf_2 clkbuf_leaf_180_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_180_clk));
 sg13g2_buf_2 clkbuf_leaf_181_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_181_clk));
 sg13g2_buf_2 clkbuf_leaf_182_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_182_clk));
 sg13g2_buf_2 clkbuf_leaf_183_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_183_clk));
 sg13g2_buf_2 clkbuf_leaf_184_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_184_clk));
 sg13g2_buf_2 clkbuf_leaf_185_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_185_clk));
 sg13g2_buf_2 clkbuf_leaf_186_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_186_clk));
 sg13g2_buf_2 clkbuf_leaf_187_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_187_clk));
 sg13g2_buf_2 clkbuf_leaf_188_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_188_clk));
 sg13g2_buf_2 clkbuf_leaf_189_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_189_clk));
 sg13g2_buf_2 clkbuf_leaf_190_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_190_clk));
 sg13g2_buf_2 clkbuf_leaf_191_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_191_clk));
 sg13g2_buf_2 clkbuf_leaf_192_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_192_clk));
 sg13g2_buf_2 clkbuf_leaf_193_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_193_clk));
 sg13g2_buf_2 clkbuf_leaf_194_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_194_clk));
 sg13g2_buf_2 clkbuf_leaf_195_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_195_clk));
 sg13g2_buf_2 clkbuf_leaf_196_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_196_clk));
 sg13g2_buf_2 clkbuf_leaf_197_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_197_clk));
 sg13g2_buf_2 clkbuf_leaf_198_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_198_clk));
 sg13g2_buf_2 clkbuf_leaf_199_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_199_clk));
 sg13g2_buf_2 clkbuf_leaf_200_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_200_clk));
 sg13g2_buf_2 clkbuf_leaf_201_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_201_clk));
 sg13g2_buf_2 clkbuf_leaf_202_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_202_clk));
 sg13g2_buf_2 clkbuf_leaf_203_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_203_clk));
 sg13g2_buf_2 clkbuf_leaf_204_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_204_clk));
 sg13g2_buf_2 clkbuf_leaf_205_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_205_clk));
 sg13g2_buf_2 clkbuf_leaf_206_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_206_clk));
 sg13g2_buf_2 clkbuf_leaf_207_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_207_clk));
 sg13g2_buf_2 clkbuf_leaf_208_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_208_clk));
 sg13g2_buf_2 clkbuf_leaf_209_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_209_clk));
 sg13g2_buf_2 clkbuf_leaf_210_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_210_clk));
 sg13g2_buf_2 clkbuf_leaf_211_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_211_clk));
 sg13g2_buf_2 clkbuf_leaf_212_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_212_clk));
 sg13g2_buf_2 clkbuf_leaf_213_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_213_clk));
 sg13g2_buf_2 clkbuf_leaf_214_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_214_clk));
 sg13g2_buf_2 clkbuf_leaf_215_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_215_clk));
 sg13g2_buf_2 clkbuf_leaf_216_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_216_clk));
 sg13g2_buf_2 clkbuf_leaf_217_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_217_clk));
 sg13g2_buf_2 clkbuf_leaf_218_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_218_clk));
 sg13g2_buf_2 clkbuf_leaf_219_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_219_clk));
 sg13g2_buf_2 clkbuf_leaf_220_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_220_clk));
 sg13g2_buf_2 clkbuf_leaf_221_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_221_clk));
 sg13g2_buf_2 clkbuf_leaf_222_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_222_clk));
 sg13g2_buf_2 clkbuf_leaf_223_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_223_clk));
 sg13g2_buf_2 clkbuf_leaf_224_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_224_clk));
 sg13g2_buf_2 clkbuf_leaf_225_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_225_clk));
 sg13g2_buf_2 clkbuf_leaf_226_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_226_clk));
 sg13g2_buf_2 clkbuf_leaf_227_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_227_clk));
 sg13g2_buf_2 clkbuf_leaf_228_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_228_clk));
 sg13g2_buf_2 clkbuf_leaf_229_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_229_clk));
 sg13g2_buf_2 clkbuf_leaf_230_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_230_clk));
 sg13g2_buf_2 clkbuf_leaf_231_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_231_clk));
 sg13g2_buf_2 clkbuf_leaf_232_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_232_clk));
 sg13g2_buf_2 clkbuf_leaf_233_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_233_clk));
 sg13g2_buf_2 clkbuf_leaf_234_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_234_clk));
 sg13g2_buf_2 clkbuf_leaf_235_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_235_clk));
 sg13g2_buf_2 clkbuf_leaf_236_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_236_clk));
 sg13g2_buf_2 clkbuf_leaf_237_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_237_clk));
 sg13g2_buf_2 clkbuf_leaf_238_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_238_clk));
 sg13g2_buf_2 clkbuf_leaf_239_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_239_clk));
 sg13g2_buf_2 clkbuf_leaf_240_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_240_clk));
 sg13g2_buf_2 clkbuf_leaf_241_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_241_clk));
 sg13g2_buf_2 clkbuf_leaf_242_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_242_clk));
 sg13g2_buf_2 clkbuf_leaf_243_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_243_clk));
 sg13g2_buf_2 clkbuf_leaf_244_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_244_clk));
 sg13g2_buf_2 clkbuf_leaf_245_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_245_clk));
 sg13g2_buf_2 clkbuf_leaf_246_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_246_clk));
 sg13g2_buf_2 clkbuf_leaf_247_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_247_clk));
 sg13g2_buf_2 clkbuf_leaf_248_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_248_clk));
 sg13g2_buf_2 clkbuf_leaf_249_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_249_clk));
 sg13g2_buf_2 clkbuf_leaf_250_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_250_clk));
 sg13g2_buf_2 clkbuf_leaf_251_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_251_clk));
 sg13g2_buf_2 clkbuf_leaf_252_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_252_clk));
 sg13g2_buf_2 clkbuf_leaf_253_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_253_clk));
 sg13g2_buf_2 clkbuf_leaf_254_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_254_clk));
 sg13g2_buf_2 clkbuf_leaf_255_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_255_clk));
 sg13g2_buf_2 clkbuf_leaf_256_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_256_clk));
 sg13g2_buf_2 clkbuf_leaf_257_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_257_clk));
 sg13g2_buf_2 clkbuf_leaf_258_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_258_clk));
 sg13g2_buf_2 clkbuf_leaf_259_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_259_clk));
 sg13g2_buf_2 clkbuf_leaf_260_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_260_clk));
 sg13g2_buf_2 clkbuf_leaf_261_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_261_clk));
 sg13g2_buf_2 clkbuf_leaf_262_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_262_clk));
 sg13g2_buf_2 clkbuf_leaf_263_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_263_clk));
 sg13g2_buf_2 clkbuf_leaf_264_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_264_clk));
 sg13g2_buf_2 clkbuf_leaf_265_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_265_clk));
 sg13g2_buf_2 clkbuf_leaf_266_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_266_clk));
 sg13g2_buf_2 clkbuf_leaf_267_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_267_clk));
 sg13g2_buf_2 clkbuf_leaf_268_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_268_clk));
 sg13g2_buf_2 clkbuf_leaf_269_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_269_clk));
 sg13g2_buf_2 clkbuf_leaf_270_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_270_clk));
 sg13g2_buf_2 clkbuf_leaf_271_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_271_clk));
 sg13g2_buf_2 clkbuf_leaf_272_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_272_clk));
 sg13g2_buf_2 clkbuf_leaf_273_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_273_clk));
 sg13g2_buf_2 clkbuf_leaf_274_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_274_clk));
 sg13g2_buf_2 clkbuf_leaf_275_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_275_clk));
 sg13g2_buf_2 clkbuf_leaf_276_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_276_clk));
 sg13g2_buf_2 clkbuf_leaf_277_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_277_clk));
 sg13g2_buf_2 clkbuf_leaf_278_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_278_clk));
 sg13g2_buf_2 clkbuf_leaf_279_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_279_clk));
 sg13g2_buf_2 clkbuf_leaf_280_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_280_clk));
 sg13g2_buf_2 clkbuf_leaf_281_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_281_clk));
 sg13g2_buf_2 clkbuf_leaf_282_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_282_clk));
 sg13g2_buf_2 clkbuf_leaf_283_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_283_clk));
 sg13g2_buf_2 clkbuf_leaf_284_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_284_clk));
 sg13g2_buf_2 clkbuf_leaf_285_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_285_clk));
 sg13g2_buf_2 clkbuf_leaf_286_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_286_clk));
 sg13g2_buf_2 clkbuf_leaf_287_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_287_clk));
 sg13g2_buf_2 clkbuf_leaf_288_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_288_clk));
 sg13g2_buf_2 clkbuf_leaf_289_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_289_clk));
 sg13g2_buf_2 clkbuf_leaf_290_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_290_clk));
 sg13g2_buf_2 clkbuf_leaf_291_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_291_clk));
 sg13g2_buf_2 clkbuf_leaf_292_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_292_clk));
 sg13g2_buf_2 clkbuf_leaf_293_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_293_clk));
 sg13g2_buf_2 clkbuf_leaf_294_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_294_clk));
 sg13g2_buf_2 clkbuf_leaf_295_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_295_clk));
 sg13g2_buf_2 clkbuf_leaf_296_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_296_clk));
 sg13g2_buf_2 clkbuf_leaf_297_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_297_clk));
 sg13g2_buf_2 clkbuf_leaf_298_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_298_clk));
 sg13g2_buf_2 clkbuf_leaf_299_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_299_clk));
 sg13g2_buf_2 clkbuf_leaf_300_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_300_clk));
 sg13g2_buf_2 clkbuf_leaf_301_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_301_clk));
 sg13g2_buf_2 clkbuf_leaf_302_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_302_clk));
 sg13g2_buf_2 clkbuf_leaf_303_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_303_clk));
 sg13g2_buf_2 clkbuf_leaf_304_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_304_clk));
 sg13g2_buf_2 clkbuf_leaf_305_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_305_clk));
 sg13g2_buf_2 clkbuf_leaf_306_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_306_clk));
 sg13g2_buf_2 clkbuf_leaf_307_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_307_clk));
 sg13g2_buf_2 clkbuf_leaf_308_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_308_clk));
 sg13g2_buf_2 clkbuf_leaf_309_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_309_clk));
 sg13g2_buf_2 clkbuf_leaf_310_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_310_clk));
 sg13g2_buf_2 clkbuf_leaf_311_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_311_clk));
 sg13g2_buf_2 clkbuf_leaf_312_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_312_clk));
 sg13g2_buf_2 clkbuf_leaf_313_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_313_clk));
 sg13g2_buf_2 clkbuf_leaf_314_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_314_clk));
 sg13g2_buf_2 clkbuf_leaf_315_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_315_clk));
 sg13g2_buf_2 clkbuf_leaf_316_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_316_clk));
 sg13g2_buf_2 clkbuf_leaf_317_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_317_clk));
 sg13g2_buf_2 clkbuf_leaf_318_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_318_clk));
 sg13g2_buf_2 clkbuf_leaf_319_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_319_clk));
 sg13g2_buf_2 clkbuf_leaf_320_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_320_clk));
 sg13g2_buf_2 clkbuf_leaf_321_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_321_clk));
 sg13g2_buf_2 clkbuf_leaf_322_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_322_clk));
 sg13g2_buf_2 clkbuf_leaf_323_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_323_clk));
 sg13g2_buf_2 clkbuf_leaf_324_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_324_clk));
 sg13g2_buf_2 clkbuf_leaf_325_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_325_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_2_0_0_clk (.A(clknet_0_clk),
    .X(clknet_2_0_0_clk));
 sg13g2_buf_2 clkbuf_2_1_0_clk (.A(clknet_0_clk),
    .X(clknet_2_1_0_clk));
 sg13g2_buf_2 clkbuf_2_2_0_clk (.A(clknet_0_clk),
    .X(clknet_2_2_0_clk));
 sg13g2_buf_2 clkbuf_2_3_0_clk (.A(clknet_0_clk),
    .X(clknet_2_3_0_clk));
 sg13g2_buf_2 clkbuf_5_0_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_0_0_clk));
 sg13g2_buf_2 clkbuf_5_1_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_1_0_clk));
 sg13g2_buf_2 clkbuf_5_2_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_2_0_clk));
 sg13g2_buf_2 clkbuf_5_3_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_3_0_clk));
 sg13g2_buf_2 clkbuf_5_4_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_4_0_clk));
 sg13g2_buf_2 clkbuf_5_5_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_5_0_clk));
 sg13g2_buf_2 clkbuf_5_6_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_6_0_clk));
 sg13g2_buf_2 clkbuf_5_7_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_7_0_clk));
 sg13g2_buf_2 clkbuf_5_8_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_8_0_clk));
 sg13g2_buf_2 clkbuf_5_9_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_9_0_clk));
 sg13g2_buf_2 clkbuf_5_10_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_10_0_clk));
 sg13g2_buf_2 clkbuf_5_11_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_11_0_clk));
 sg13g2_buf_2 clkbuf_5_12_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_12_0_clk));
 sg13g2_buf_2 clkbuf_5_13_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_13_0_clk));
 sg13g2_buf_2 clkbuf_5_14_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_14_0_clk));
 sg13g2_buf_2 clkbuf_5_15_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_15_0_clk));
 sg13g2_buf_2 clkbuf_5_16_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_16_0_clk));
 sg13g2_buf_2 clkbuf_5_17_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_17_0_clk));
 sg13g2_buf_2 clkbuf_5_18_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_18_0_clk));
 sg13g2_buf_2 clkbuf_5_19_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_19_0_clk));
 sg13g2_buf_2 clkbuf_5_20_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_20_0_clk));
 sg13g2_buf_2 clkbuf_5_21_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_21_0_clk));
 sg13g2_buf_2 clkbuf_5_22_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_22_0_clk));
 sg13g2_buf_2 clkbuf_5_23_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_23_0_clk));
 sg13g2_buf_2 clkbuf_5_24_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_24_0_clk));
 sg13g2_buf_2 clkbuf_5_25_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_25_0_clk));
 sg13g2_buf_2 clkbuf_5_26_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_26_0_clk));
 sg13g2_buf_2 clkbuf_5_27_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_27_0_clk));
 sg13g2_buf_2 clkbuf_5_28_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_28_0_clk));
 sg13g2_buf_2 clkbuf_5_29_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_29_0_clk));
 sg13g2_buf_2 clkbuf_5_30_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_30_0_clk));
 sg13g2_buf_2 clkbuf_5_31_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_31_0_clk));
 sg13g2_buf_2 clkbuf_6_0__f_clk (.A(clknet_5_0_0_clk),
    .X(clknet_6_0__leaf_clk));
 sg13g2_buf_2 clkbuf_6_1__f_clk (.A(clknet_5_0_0_clk),
    .X(clknet_6_1__leaf_clk));
 sg13g2_buf_2 clkbuf_6_2__f_clk (.A(clknet_5_1_0_clk),
    .X(clknet_6_2__leaf_clk));
 sg13g2_buf_2 clkbuf_6_3__f_clk (.A(clknet_5_1_0_clk),
    .X(clknet_6_3__leaf_clk));
 sg13g2_buf_2 clkbuf_6_4__f_clk (.A(clknet_5_2_0_clk),
    .X(clknet_6_4__leaf_clk));
 sg13g2_buf_2 clkbuf_6_5__f_clk (.A(clknet_5_2_0_clk),
    .X(clknet_6_5__leaf_clk));
 sg13g2_buf_2 clkbuf_6_6__f_clk (.A(clknet_5_3_0_clk),
    .X(clknet_6_6__leaf_clk));
 sg13g2_buf_2 clkbuf_6_7__f_clk (.A(clknet_5_3_0_clk),
    .X(clknet_6_7__leaf_clk));
 sg13g2_buf_2 clkbuf_6_8__f_clk (.A(clknet_5_4_0_clk),
    .X(clknet_6_8__leaf_clk));
 sg13g2_buf_2 clkbuf_6_9__f_clk (.A(clknet_5_4_0_clk),
    .X(clknet_6_9__leaf_clk));
 sg13g2_buf_2 clkbuf_6_10__f_clk (.A(clknet_5_5_0_clk),
    .X(clknet_6_10__leaf_clk));
 sg13g2_buf_2 clkbuf_6_11__f_clk (.A(clknet_5_5_0_clk),
    .X(clknet_6_11__leaf_clk));
 sg13g2_buf_2 clkbuf_6_12__f_clk (.A(clknet_5_6_0_clk),
    .X(clknet_6_12__leaf_clk));
 sg13g2_buf_2 clkbuf_6_13__f_clk (.A(clknet_5_6_0_clk),
    .X(clknet_6_13__leaf_clk));
 sg13g2_buf_2 clkbuf_6_14__f_clk (.A(clknet_5_7_0_clk),
    .X(clknet_6_14__leaf_clk));
 sg13g2_buf_2 clkbuf_6_15__f_clk (.A(clknet_5_7_0_clk),
    .X(clknet_6_15__leaf_clk));
 sg13g2_buf_2 clkbuf_6_16__f_clk (.A(clknet_5_8_0_clk),
    .X(clknet_6_16__leaf_clk));
 sg13g2_buf_2 clkbuf_6_17__f_clk (.A(clknet_5_8_0_clk),
    .X(clknet_6_17__leaf_clk));
 sg13g2_buf_2 clkbuf_6_18__f_clk (.A(clknet_5_9_0_clk),
    .X(clknet_6_18__leaf_clk));
 sg13g2_buf_2 clkbuf_6_19__f_clk (.A(clknet_5_9_0_clk),
    .X(clknet_6_19__leaf_clk));
 sg13g2_buf_2 clkbuf_6_20__f_clk (.A(clknet_5_10_0_clk),
    .X(clknet_6_20__leaf_clk));
 sg13g2_buf_2 clkbuf_6_21__f_clk (.A(clknet_5_10_0_clk),
    .X(clknet_6_21__leaf_clk));
 sg13g2_buf_2 clkbuf_6_22__f_clk (.A(clknet_5_11_0_clk),
    .X(clknet_6_22__leaf_clk));
 sg13g2_buf_2 clkbuf_6_23__f_clk (.A(clknet_5_11_0_clk),
    .X(clknet_6_23__leaf_clk));
 sg13g2_buf_2 clkbuf_6_24__f_clk (.A(clknet_5_12_0_clk),
    .X(clknet_6_24__leaf_clk));
 sg13g2_buf_2 clkbuf_6_25__f_clk (.A(clknet_5_12_0_clk),
    .X(clknet_6_25__leaf_clk));
 sg13g2_buf_2 clkbuf_6_26__f_clk (.A(clknet_5_13_0_clk),
    .X(clknet_6_26__leaf_clk));
 sg13g2_buf_2 clkbuf_6_27__f_clk (.A(clknet_5_13_0_clk),
    .X(clknet_6_27__leaf_clk));
 sg13g2_buf_2 clkbuf_6_28__f_clk (.A(clknet_5_14_0_clk),
    .X(clknet_6_28__leaf_clk));
 sg13g2_buf_2 clkbuf_6_29__f_clk (.A(clknet_5_14_0_clk),
    .X(clknet_6_29__leaf_clk));
 sg13g2_buf_2 clkbuf_6_30__f_clk (.A(clknet_5_15_0_clk),
    .X(clknet_6_30__leaf_clk));
 sg13g2_buf_2 clkbuf_6_31__f_clk (.A(clknet_5_15_0_clk),
    .X(clknet_6_31__leaf_clk));
 sg13g2_buf_2 clkbuf_6_32__f_clk (.A(clknet_5_16_0_clk),
    .X(clknet_6_32__leaf_clk));
 sg13g2_buf_2 clkbuf_6_33__f_clk (.A(clknet_5_16_0_clk),
    .X(clknet_6_33__leaf_clk));
 sg13g2_buf_2 clkbuf_6_34__f_clk (.A(clknet_5_17_0_clk),
    .X(clknet_6_34__leaf_clk));
 sg13g2_buf_2 clkbuf_6_35__f_clk (.A(clknet_5_17_0_clk),
    .X(clknet_6_35__leaf_clk));
 sg13g2_buf_2 clkbuf_6_36__f_clk (.A(clknet_5_18_0_clk),
    .X(clknet_6_36__leaf_clk));
 sg13g2_buf_2 clkbuf_6_37__f_clk (.A(clknet_5_18_0_clk),
    .X(clknet_6_37__leaf_clk));
 sg13g2_buf_2 clkbuf_6_38__f_clk (.A(clknet_5_19_0_clk),
    .X(clknet_6_38__leaf_clk));
 sg13g2_buf_2 clkbuf_6_39__f_clk (.A(clknet_5_19_0_clk),
    .X(clknet_6_39__leaf_clk));
 sg13g2_buf_2 clkbuf_6_40__f_clk (.A(clknet_5_20_0_clk),
    .X(clknet_6_40__leaf_clk));
 sg13g2_buf_2 clkbuf_6_41__f_clk (.A(clknet_5_20_0_clk),
    .X(clknet_6_41__leaf_clk));
 sg13g2_buf_2 clkbuf_6_42__f_clk (.A(clknet_5_21_0_clk),
    .X(clknet_6_42__leaf_clk));
 sg13g2_buf_2 clkbuf_6_43__f_clk (.A(clknet_5_21_0_clk),
    .X(clknet_6_43__leaf_clk));
 sg13g2_buf_2 clkbuf_6_44__f_clk (.A(clknet_5_22_0_clk),
    .X(clknet_6_44__leaf_clk));
 sg13g2_buf_2 clkbuf_6_45__f_clk (.A(clknet_5_22_0_clk),
    .X(clknet_6_45__leaf_clk));
 sg13g2_buf_2 clkbuf_6_46__f_clk (.A(clknet_5_23_0_clk),
    .X(clknet_6_46__leaf_clk));
 sg13g2_buf_2 clkbuf_6_47__f_clk (.A(clknet_5_23_0_clk),
    .X(clknet_6_47__leaf_clk));
 sg13g2_buf_2 clkbuf_6_48__f_clk (.A(clknet_5_24_0_clk),
    .X(clknet_6_48__leaf_clk));
 sg13g2_buf_2 clkbuf_6_49__f_clk (.A(clknet_5_24_0_clk),
    .X(clknet_6_49__leaf_clk));
 sg13g2_buf_2 clkbuf_6_50__f_clk (.A(clknet_5_25_0_clk),
    .X(clknet_6_50__leaf_clk));
 sg13g2_buf_2 clkbuf_6_51__f_clk (.A(clknet_5_25_0_clk),
    .X(clknet_6_51__leaf_clk));
 sg13g2_buf_2 clkbuf_6_52__f_clk (.A(clknet_5_26_0_clk),
    .X(clknet_6_52__leaf_clk));
 sg13g2_buf_2 clkbuf_6_53__f_clk (.A(clknet_5_26_0_clk),
    .X(clknet_6_53__leaf_clk));
 sg13g2_buf_2 clkbuf_6_54__f_clk (.A(clknet_5_27_0_clk),
    .X(clknet_6_54__leaf_clk));
 sg13g2_buf_2 clkbuf_6_55__f_clk (.A(clknet_5_27_0_clk),
    .X(clknet_6_55__leaf_clk));
 sg13g2_buf_2 clkbuf_6_56__f_clk (.A(clknet_5_28_0_clk),
    .X(clknet_6_56__leaf_clk));
 sg13g2_buf_2 clkbuf_6_57__f_clk (.A(clknet_5_28_0_clk),
    .X(clknet_6_57__leaf_clk));
 sg13g2_buf_2 clkbuf_6_58__f_clk (.A(clknet_5_29_0_clk),
    .X(clknet_6_58__leaf_clk));
 sg13g2_buf_2 clkbuf_6_59__f_clk (.A(clknet_5_29_0_clk),
    .X(clknet_6_59__leaf_clk));
 sg13g2_buf_2 clkbuf_6_60__f_clk (.A(clknet_5_30_0_clk),
    .X(clknet_6_60__leaf_clk));
 sg13g2_buf_2 clkbuf_6_61__f_clk (.A(clknet_5_30_0_clk),
    .X(clknet_6_61__leaf_clk));
 sg13g2_buf_2 clkbuf_6_62__f_clk (.A(clknet_5_31_0_clk),
    .X(clknet_6_62__leaf_clk));
 sg13g2_buf_2 clkbuf_6_63__f_clk (.A(clknet_5_31_0_clk),
    .X(clknet_6_63__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_6_1__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_6_9__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_6_17__leaf_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_6_33__leaf_clk));
 sg13g2_buf_2 clkload4 (.A(clknet_6_41__leaf_clk));
 sg13g2_buf_2 clkload5 (.A(clknet_6_49__leaf_clk));
 sg13g2_inv_2 clkload6 (.A(clknet_leaf_325_clk));
 sg13g2_inv_4 clkload7 (.A(clknet_leaf_179_clk));
 sg13g2_inv_4 clkload8 (.A(clknet_leaf_142_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_leaf_138_clk));
 sg13g2_inv_4 clkload10 (.A(clknet_leaf_146_clk));
 sg13g2_inv_4 clkload11 (.A(clknet_leaf_166_clk));
 sg13g2_inv_4 clkload12 (.A(clknet_leaf_164_clk));
 sg13g2_inv_4 clkload13 (.A(clknet_leaf_161_clk));
 sg13g2_inv_4 clkload14 (.A(clknet_leaf_178_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_00301_),
    .X(net2598));
 sg13g2_dlygate4sd3_1 hold2 (.A(_01763_),
    .X(net2599));
 sg13g2_dlygate4sd3_1 hold3 (.A(_00304_),
    .X(net2600));
 sg13g2_dlygate4sd3_1 hold4 (.A(_00283_),
    .X(net2601));
 sg13g2_dlygate4sd3_1 hold5 (.A(_02141_),
    .X(net2602));
 sg13g2_dlygate4sd3_1 hold6 (.A(_00303_),
    .X(net2603));
 sg13g2_dlygate4sd3_1 hold7 (.A(_00299_),
    .X(net2604));
 sg13g2_dlygate4sd3_1 hold8 (.A(_01859_),
    .X(net2605));
 sg13g2_dlygate4sd3_1 hold9 (.A(_00298_),
    .X(net2606));
 sg13g2_dlygate4sd3_1 hold10 (.A(_01863_),
    .X(net2607));
 sg13g2_dlygate4sd3_1 hold11 (.A(_00297_),
    .X(net2608));
 sg13g2_dlygate4sd3_1 hold12 (.A(_01873_),
    .X(net2609));
 sg13g2_dlygate4sd3_1 hold13 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][31] ),
    .X(net2610));
 sg13g2_dlygate4sd3_1 hold14 (.A(\soc_I.rx_uart_i.return_state[0] ),
    .X(net2611));
 sg13g2_dlygate4sd3_1 hold15 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][9] ),
    .X(net2612));
 sg13g2_dlygate4sd3_1 hold16 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][25] ),
    .X(net2613));
 sg13g2_dlygate4sd3_1 hold17 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][6] ),
    .X(net2614));
 sg13g2_dlygate4sd3_1 hold18 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][15] ),
    .X(net2615));
 sg13g2_dlygate4sd3_1 hold19 (.A(_00284_),
    .X(net2616));
 sg13g2_dlygate4sd3_1 hold20 (.A(_02142_),
    .X(net2617));
 sg13g2_dlygate4sd3_1 hold21 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][19] ),
    .X(net2618));
 sg13g2_dlygate4sd3_1 hold22 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][16] ),
    .X(net2619));
 sg13g2_dlygate4sd3_1 hold23 (.A(\soc_I.rx_uart_i.fifo_i.ram[8][0] ),
    .X(net2620));
 sg13g2_dlygate4sd3_1 hold24 (.A(_07433_),
    .X(net2621));
 sg13g2_dlygate4sd3_1 hold25 (.A(_02100_),
    .X(net2622));
 sg13g2_dlygate4sd3_1 hold26 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][3] ),
    .X(net2623));
 sg13g2_dlygate4sd3_1 hold27 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][15] ),
    .X(net2624));
 sg13g2_dlygate4sd3_1 hold28 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][23] ),
    .X(net2625));
 sg13g2_dlygate4sd3_1 hold29 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][14] ),
    .X(net2626));
 sg13g2_dlygate4sd3_1 hold30 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][20] ),
    .X(net2627));
 sg13g2_dlygate4sd3_1 hold31 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][5] ),
    .X(net2628));
 sg13g2_dlygate4sd3_1 hold32 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][13] ),
    .X(net2629));
 sg13g2_dlygate4sd3_1 hold33 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[5] ),
    .X(net2630));
 sg13g2_dlygate4sd3_1 hold34 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[4] ),
    .X(net2631));
 sg13g2_dlygate4sd3_1 hold35 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][17] ),
    .X(net2632));
 sg13g2_dlygate4sd3_1 hold36 (.A(\soc_I.rx_uart_i.wait_states[16] ),
    .X(net2633));
 sg13g2_dlygate4sd3_1 hold37 (.A(_01858_),
    .X(net2634));
 sg13g2_dlygate4sd3_1 hold38 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[4] ),
    .X(net2635));
 sg13g2_dlygate4sd3_1 hold39 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][1] ),
    .X(net2636));
 sg13g2_dlygate4sd3_1 hold40 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][1] ),
    .X(net2637));
 sg13g2_dlygate4sd3_1 hold41 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[20] ),
    .X(net2638));
 sg13g2_dlygate4sd3_1 hold42 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][8] ),
    .X(net2639));
 sg13g2_dlygate4sd3_1 hold43 (.A(\soc_I.qqspi_I.rdata[15] ),
    .X(net2640));
 sg13g2_dlygate4sd3_1 hold44 (.A(_01811_),
    .X(net2641));
 sg13g2_dlygate4sd3_1 hold45 (.A(\soc_I.rx_uart_i.fifo_i.ram[7][0] ),
    .X(net2642));
 sg13g2_dlygate4sd3_1 hold46 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[29] ),
    .X(net2643));
 sg13g2_dlygate4sd3_1 hold47 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][14] ),
    .X(net2644));
 sg13g2_dlygate4sd3_1 hold48 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][0] ),
    .X(net2645));
 sg13g2_dlygate4sd3_1 hold49 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][28] ),
    .X(net2646));
 sg13g2_dlygate4sd3_1 hold50 (.A(\soc_I.rx_uart_i.fifo_i.ram[12][0] ),
    .X(net2647));
 sg13g2_dlygate4sd3_1 hold51 (.A(_02809_),
    .X(net2648));
 sg13g2_dlygate4sd3_1 hold52 (.A(_00654_),
    .X(net2649));
 sg13g2_dlygate4sd3_1 hold53 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[26] ),
    .X(net2650));
 sg13g2_dlygate4sd3_1 hold54 (.A(\soc_I.rx_uart_i.fifo_i.ram[3][0] ),
    .X(net2651));
 sg13g2_dlygate4sd3_1 hold55 (.A(\soc_I.rx_uart_i.fifo_i.ram[4][0] ),
    .X(net2652));
 sg13g2_dlygate4sd3_1 hold56 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][28] ),
    .X(net2653));
 sg13g2_dlygate4sd3_1 hold57 (.A(\soc_I.qqspi_I.rdata[11] ),
    .X(net2654));
 sg13g2_dlygate4sd3_1 hold58 (.A(_01807_),
    .X(net2655));
 sg13g2_dlygate4sd3_1 hold59 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[11] ),
    .X(net2656));
 sg13g2_dlygate4sd3_1 hold60 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][13] ),
    .X(net2657));
 sg13g2_dlygate4sd3_1 hold61 (.A(\soc_I.rx_uart_i.fifo_i.ram[0][0] ),
    .X(net2658));
 sg13g2_dlygate4sd3_1 hold62 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][26] ),
    .X(net2659));
 sg13g2_dlygate4sd3_1 hold63 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[23] ),
    .X(net2660));
 sg13g2_dlygate4sd3_1 hold64 (.A(\soc_I.rx_uart_i.fifo_i.ram[2][0] ),
    .X(net2661));
 sg13g2_dlygate4sd3_1 hold65 (.A(_01081_),
    .X(net2662));
 sg13g2_dlygate4sd3_1 hold66 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[9] ),
    .X(net2663));
 sg13g2_dlygate4sd3_1 hold67 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[31] ),
    .X(net2664));
 sg13g2_dlygate4sd3_1 hold68 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[28] ),
    .X(net2665));
 sg13g2_dlygate4sd3_1 hold69 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][11] ),
    .X(net2666));
 sg13g2_dlygate4sd3_1 hold70 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[21] ),
    .X(net2667));
 sg13g2_dlygate4sd3_1 hold71 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[22] ),
    .X(net2668));
 sg13g2_dlygate4sd3_1 hold72 (.A(\soc_I.qqspi_I.rdata[25] ),
    .X(net2669));
 sg13g2_dlygate4sd3_1 hold73 (.A(_01821_),
    .X(net2670));
 sg13g2_dlygate4sd3_1 hold74 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][24] ),
    .X(net2671));
 sg13g2_dlygate4sd3_1 hold75 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][19] ),
    .X(net2672));
 sg13g2_dlygate4sd3_1 hold76 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][2] ),
    .X(net2673));
 sg13g2_dlygate4sd3_1 hold77 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][24] ),
    .X(net2674));
 sg13g2_dlygate4sd3_1 hold78 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][16] ),
    .X(net2675));
 sg13g2_dlygate4sd3_1 hold79 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][19] ),
    .X(net2676));
 sg13g2_dlygate4sd3_1 hold80 (.A(\soc_I.qqspi_I.rdata[2] ),
    .X(net2677));
 sg13g2_dlygate4sd3_1 hold81 (.A(_01798_),
    .X(net2678));
 sg13g2_dlygate4sd3_1 hold82 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][0] ),
    .X(net2679));
 sg13g2_dlygate4sd3_1 hold83 (.A(_00305_),
    .X(net2680));
 sg13g2_dlygate4sd3_1 hold84 (.A(_01137_),
    .X(net2681));
 sg13g2_dlygate4sd3_1 hold85 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][30] ),
    .X(net2682));
 sg13g2_dlygate4sd3_1 hold86 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[28] ),
    .X(net2683));
 sg13g2_dlygate4sd3_1 hold87 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][20] ),
    .X(net2684));
 sg13g2_dlygate4sd3_1 hold88 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][9] ),
    .X(net2685));
 sg13g2_dlygate4sd3_1 hold89 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][1] ),
    .X(net2686));
 sg13g2_dlygate4sd3_1 hold90 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[18] ),
    .X(net2687));
 sg13g2_dlygate4sd3_1 hold91 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][21] ),
    .X(net2688));
 sg13g2_dlygate4sd3_1 hold92 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][21] ),
    .X(net2689));
 sg13g2_dlygate4sd3_1 hold93 (.A(\soc_I.qqspi_I.rdata[27] ),
    .X(net2690));
 sg13g2_dlygate4sd3_1 hold94 (.A(_01823_),
    .X(net2691));
 sg13g2_dlygate4sd3_1 hold95 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][29] ),
    .X(net2692));
 sg13g2_dlygate4sd3_1 hold96 (.A(\soc_I.qqspi_I.rdata[28] ),
    .X(net2693));
 sg13g2_dlygate4sd3_1 hold97 (.A(_01824_),
    .X(net2694));
 sg13g2_dlygate4sd3_1 hold98 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][20] ),
    .X(net2695));
 sg13g2_dlygate4sd3_1 hold99 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[12] ),
    .X(net2696));
 sg13g2_dlygate4sd3_1 hold100 (.A(\soc_I.qqspi_I.rdata[6] ),
    .X(net2697));
 sg13g2_dlygate4sd3_1 hold101 (.A(_01802_),
    .X(net2698));
 sg13g2_dlygate4sd3_1 hold102 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][20] ),
    .X(net2699));
 sg13g2_dlygate4sd3_1 hold103 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][30] ),
    .X(net2700));
 sg13g2_dlygate4sd3_1 hold104 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][14] ),
    .X(net2701));
 sg13g2_dlygate4sd3_1 hold105 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][22] ),
    .X(net2702));
 sg13g2_dlygate4sd3_1 hold106 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[25] ),
    .X(net2703));
 sg13g2_dlygate4sd3_1 hold107 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][2] ),
    .X(net2704));
 sg13g2_dlygate4sd3_1 hold108 (.A(\soc_I.qqspi_I.rdata[16] ),
    .X(net2705));
 sg13g2_dlygate4sd3_1 hold109 (.A(_01812_),
    .X(net2706));
 sg13g2_dlygate4sd3_1 hold110 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][18] ),
    .X(net2707));
 sg13g2_dlygate4sd3_1 hold111 (.A(\soc_I.rx_uart_i.fifo_i.ram[5][0] ),
    .X(net2708));
 sg13g2_dlygate4sd3_1 hold112 (.A(\soc_I.rx_uart_i.fifo_i.ram[11][0] ),
    .X(net2709));
 sg13g2_dlygate4sd3_1 hold113 (.A(_02807_),
    .X(net2710));
 sg13g2_dlygate4sd3_1 hold114 (.A(_00646_),
    .X(net2711));
 sg13g2_dlygate4sd3_1 hold115 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][25] ),
    .X(net2712));
 sg13g2_dlygate4sd3_1 hold116 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][28] ),
    .X(net2713));
 sg13g2_dlygate4sd3_1 hold117 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][17] ),
    .X(net2714));
 sg13g2_dlygate4sd3_1 hold118 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[9] ),
    .X(net2715));
 sg13g2_dlygate4sd3_1 hold119 (.A(\soc_I.rx_uart_i.fifo_i.ram[1][0] ),
    .X(net2716));
 sg13g2_dlygate4sd3_1 hold120 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][21] ),
    .X(net2717));
 sg13g2_dlygate4sd3_1 hold121 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][24] ),
    .X(net2718));
 sg13g2_dlygate4sd3_1 hold122 (.A(\soc_I.qqspi_I.rdata[19] ),
    .X(net2719));
 sg13g2_dlygate4sd3_1 hold123 (.A(_01815_),
    .X(net2720));
 sg13g2_dlygate4sd3_1 hold124 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][20] ),
    .X(net2721));
 sg13g2_dlygate4sd3_1 hold125 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][7] ),
    .X(net2722));
 sg13g2_dlygate4sd3_1 hold126 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][23] ),
    .X(net2723));
 sg13g2_dlygate4sd3_1 hold127 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][23] ),
    .X(net2724));
 sg13g2_dlygate4sd3_1 hold128 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[7] ),
    .X(net2725));
 sg13g2_dlygate4sd3_1 hold129 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[30] ),
    .X(net2726));
 sg13g2_dlygate4sd3_1 hold130 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][22] ),
    .X(net2727));
 sg13g2_dlygate4sd3_1 hold131 (.A(\soc_I.rx_uart_i.rx_in_sync[0] ),
    .X(net2728));
 sg13g2_dlygate4sd3_1 hold132 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][14] ),
    .X(net2729));
 sg13g2_dlygate4sd3_1 hold133 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][8] ),
    .X(net2730));
 sg13g2_dlygate4sd3_1 hold134 (.A(\soc_I.rx_uart_i.fifo_i.ram[14][2] ),
    .X(net2731));
 sg13g2_dlygate4sd3_1 hold135 (.A(_00672_),
    .X(net2732));
 sg13g2_dlygate4sd3_1 hold136 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][13] ),
    .X(net2733));
 sg13g2_dlygate4sd3_1 hold137 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][20] ),
    .X(net2734));
 sg13g2_dlygate4sd3_1 hold138 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][12] ),
    .X(net2735));
 sg13g2_dlygate4sd3_1 hold139 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[11] ),
    .X(net2736));
 sg13g2_dlygate4sd3_1 hold140 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][24] ),
    .X(net2737));
 sg13g2_dlygate4sd3_1 hold141 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][11] ),
    .X(net2738));
 sg13g2_dlygate4sd3_1 hold142 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[30] ),
    .X(net2739));
 sg13g2_dlygate4sd3_1 hold143 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[14] ),
    .X(net2740));
 sg13g2_dlygate4sd3_1 hold144 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[16] ),
    .X(net2741));
 sg13g2_dlygate4sd3_1 hold145 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][21] ),
    .X(net2742));
 sg13g2_dlygate4sd3_1 hold146 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][5] ),
    .X(net2743));
 sg13g2_dlygate4sd3_1 hold147 (.A(\soc_I.rx_uart_i.fifo_i.ram[10][0] ),
    .X(net2744));
 sg13g2_dlygate4sd3_1 hold148 (.A(_00638_),
    .X(net2745));
 sg13g2_dlygate4sd3_1 hold149 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[27] ),
    .X(net2746));
 sg13g2_dlygate4sd3_1 hold150 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][4] ),
    .X(net2747));
 sg13g2_dlygate4sd3_1 hold151 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][27] ),
    .X(net2748));
 sg13g2_dlygate4sd3_1 hold152 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][0] ),
    .X(net2749));
 sg13g2_dlygate4sd3_1 hold153 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][12] ),
    .X(net2750));
 sg13g2_dlygate4sd3_1 hold154 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[8] ),
    .X(net2751));
 sg13g2_dlygate4sd3_1 hold155 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][28] ),
    .X(net2752));
 sg13g2_dlygate4sd3_1 hold156 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][17] ),
    .X(net2753));
 sg13g2_dlygate4sd3_1 hold157 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][12] ),
    .X(net2754));
 sg13g2_dlygate4sd3_1 hold158 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[29] ),
    .X(net2755));
 sg13g2_dlygate4sd3_1 hold159 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][4] ),
    .X(net2756));
 sg13g2_dlygate4sd3_1 hold160 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][10] ),
    .X(net2757));
 sg13g2_dlygate4sd3_1 hold161 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][5] ),
    .X(net2758));
 sg13g2_dlygate4sd3_1 hold162 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[18] ),
    .X(net2759));
 sg13g2_dlygate4sd3_1 hold163 (.A(\soc_I.rx_uart_i.fifo_i.ram[15][0] ),
    .X(net2760));
 sg13g2_dlygate4sd3_1 hold164 (.A(_01097_),
    .X(net2761));
 sg13g2_dlygate4sd3_1 hold165 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][9] ),
    .X(net2762));
 sg13g2_dlygate4sd3_1 hold166 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][25] ),
    .X(net2763));
 sg13g2_dlygate4sd3_1 hold167 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][13] ),
    .X(net2764));
 sg13g2_dlygate4sd3_1 hold168 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][7] ),
    .X(net2765));
 sg13g2_dlygate4sd3_1 hold169 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][19] ),
    .X(net2766));
 sg13g2_dlygate4sd3_1 hold170 (.A(\soc_I.qqspi_I.rdata[21] ),
    .X(net2767));
 sg13g2_dlygate4sd3_1 hold171 (.A(_01817_),
    .X(net2768));
 sg13g2_dlygate4sd3_1 hold172 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][0] ),
    .X(net2769));
 sg13g2_dlygate4sd3_1 hold173 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][4] ),
    .X(net2770));
 sg13g2_dlygate4sd3_1 hold174 (.A(\soc_I.rx_uart_i.fifo_i.ram[14][5] ),
    .X(net2771));
 sg13g2_dlygate4sd3_1 hold175 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[24] ),
    .X(net2772));
 sg13g2_dlygate4sd3_1 hold176 (.A(\soc_I.qqspi_I.rdata[30] ),
    .X(net2773));
 sg13g2_dlygate4sd3_1 hold177 (.A(_01826_),
    .X(net2774));
 sg13g2_dlygate4sd3_1 hold178 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][17] ),
    .X(net2775));
 sg13g2_dlygate4sd3_1 hold179 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][17] ),
    .X(net2776));
 sg13g2_dlygate4sd3_1 hold180 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[17] ),
    .X(net2777));
 sg13g2_dlygate4sd3_1 hold181 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][14] ),
    .X(net2778));
 sg13g2_dlygate4sd3_1 hold182 (.A(\soc_I.qqspi_I.rdata[26] ),
    .X(net2779));
 sg13g2_dlygate4sd3_1 hold183 (.A(_01822_),
    .X(net2780));
 sg13g2_dlygate4sd3_1 hold184 (.A(\soc_I.qqspi_I.rdata[18] ),
    .X(net2781));
 sg13g2_dlygate4sd3_1 hold185 (.A(_01814_),
    .X(net2782));
 sg13g2_dlygate4sd3_1 hold186 (.A(\soc_I.qqspi_I.rdata[5] ),
    .X(net2783));
 sg13g2_dlygate4sd3_1 hold187 (.A(_01801_),
    .X(net2784));
 sg13g2_dlygate4sd3_1 hold188 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][4] ),
    .X(net2785));
 sg13g2_dlygate4sd3_1 hold189 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][8] ),
    .X(net2786));
 sg13g2_dlygate4sd3_1 hold190 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][2] ),
    .X(net2787));
 sg13g2_dlygate4sd3_1 hold191 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][6] ),
    .X(net2788));
 sg13g2_dlygate4sd3_1 hold192 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][30] ),
    .X(net2789));
 sg13g2_dlygate4sd3_1 hold193 (.A(\soc_I.qqspi_I.rdata[31] ),
    .X(net2790));
 sg13g2_dlygate4sd3_1 hold194 (.A(_01827_),
    .X(net2791));
 sg13g2_dlygate4sd3_1 hold195 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][28] ),
    .X(net2792));
 sg13g2_dlygate4sd3_1 hold196 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][28] ),
    .X(net2793));
 sg13g2_dlygate4sd3_1 hold197 (.A(\soc_I.rst_cnt[0] ),
    .X(net2794));
 sg13g2_dlygate4sd3_1 hold198 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][31] ),
    .X(net2795));
 sg13g2_dlygate4sd3_1 hold199 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][18] ),
    .X(net2796));
 sg13g2_dlygate4sd3_1 hold200 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][9] ),
    .X(net2797));
 sg13g2_dlygate4sd3_1 hold201 (.A(\soc_I.rx_uart_i.fifo_i.ram[9][0] ),
    .X(net2798));
 sg13g2_dlygate4sd3_1 hold202 (.A(_07002_),
    .X(net2799));
 sg13g2_dlygate4sd3_1 hold203 (.A(_01884_),
    .X(net2800));
 sg13g2_dlygate4sd3_1 hold204 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][27] ),
    .X(net2801));
 sg13g2_dlygate4sd3_1 hold205 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[8] ),
    .X(net2802));
 sg13g2_dlygate4sd3_1 hold206 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[15] ),
    .X(net2803));
 sg13g2_dlygate4sd3_1 hold207 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][7] ),
    .X(net2804));
 sg13g2_dlygate4sd3_1 hold208 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[6] ),
    .X(net2805));
 sg13g2_dlygate4sd3_1 hold209 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][18] ),
    .X(net2806));
 sg13g2_dlygate4sd3_1 hold210 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[1] ),
    .X(net2807));
 sg13g2_dlygate4sd3_1 hold211 (.A(_04426_),
    .X(net2808));
 sg13g2_dlygate4sd3_1 hold212 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][27] ),
    .X(net2809));
 sg13g2_dlygate4sd3_1 hold213 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][8] ),
    .X(net2810));
 sg13g2_dlygate4sd3_1 hold214 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][13] ),
    .X(net2811));
 sg13g2_dlygate4sd3_1 hold215 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][4] ),
    .X(net2812));
 sg13g2_dlygate4sd3_1 hold216 (.A(\soc_I.qqspi_I.rdata[4] ),
    .X(net2813));
 sg13g2_dlygate4sd3_1 hold217 (.A(_01800_),
    .X(net2814));
 sg13g2_dlygate4sd3_1 hold218 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[25] ),
    .X(net2815));
 sg13g2_dlygate4sd3_1 hold219 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][5] ),
    .X(net2816));
 sg13g2_dlygate4sd3_1 hold220 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][31] ),
    .X(net2817));
 sg13g2_dlygate4sd3_1 hold221 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[19] ),
    .X(net2818));
 sg13g2_dlygate4sd3_1 hold222 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][10] ),
    .X(net2819));
 sg13g2_dlygate4sd3_1 hold223 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][9] ),
    .X(net2820));
 sg13g2_dlygate4sd3_1 hold224 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][28] ),
    .X(net2821));
 sg13g2_dlygate4sd3_1 hold225 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][14] ),
    .X(net2822));
 sg13g2_dlygate4sd3_1 hold226 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][6] ),
    .X(net2823));
 sg13g2_dlygate4sd3_1 hold227 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][28] ),
    .X(net2824));
 sg13g2_dlygate4sd3_1 hold228 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][11] ),
    .X(net2825));
 sg13g2_dlygate4sd3_1 hold229 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][17] ),
    .X(net2826));
 sg13g2_dlygate4sd3_1 hold230 (.A(_00727_),
    .X(net2827));
 sg13g2_dlygate4sd3_1 hold231 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[28] ),
    .X(net2828));
 sg13g2_dlygate4sd3_1 hold232 (.A(_05568_),
    .X(net2829));
 sg13g2_dlygate4sd3_1 hold233 (.A(_01293_),
    .X(net2830));
 sg13g2_dlygate4sd3_1 hold234 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][15] ),
    .X(net2831));
 sg13g2_dlygate4sd3_1 hold235 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][1] ),
    .X(net2832));
 sg13g2_dlygate4sd3_1 hold236 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][9] ),
    .X(net2833));
 sg13g2_dlygate4sd3_1 hold237 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][25] ),
    .X(net2834));
 sg13g2_dlygate4sd3_1 hold238 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][12] ),
    .X(net2835));
 sg13g2_dlygate4sd3_1 hold239 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][22] ),
    .X(net2836));
 sg13g2_dlygate4sd3_1 hold240 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][26] ),
    .X(net2837));
 sg13g2_dlygate4sd3_1 hold241 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][18] ),
    .X(net2838));
 sg13g2_dlygate4sd3_1 hold242 (.A(\soc_I.spi0_I.sio0_si_mosi ),
    .X(net2839));
 sg13g2_dlygate4sd3_1 hold243 (.A(_01753_),
    .X(net2840));
 sg13g2_dlygate4sd3_1 hold244 (.A(\soc_I.rx_uart_i.fifo_i.ram[6][0] ),
    .X(net2841));
 sg13g2_dlygate4sd3_1 hold245 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][12] ),
    .X(net2842));
 sg13g2_dlygate4sd3_1 hold246 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][13] ),
    .X(net2843));
 sg13g2_dlygate4sd3_1 hold247 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][21] ),
    .X(net2844));
 sg13g2_dlygate4sd3_1 hold248 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][5] ),
    .X(net2845));
 sg13g2_dlygate4sd3_1 hold249 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][31] ),
    .X(net2846));
 sg13g2_dlygate4sd3_1 hold250 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][0] ),
    .X(net2847));
 sg13g2_dlygate4sd3_1 hold251 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][25] ),
    .X(net2848));
 sg13g2_dlygate4sd3_1 hold252 (.A(\soc_I.qqspi_I.rdata[1] ),
    .X(net2849));
 sg13g2_dlygate4sd3_1 hold253 (.A(_01797_),
    .X(net2850));
 sg13g2_dlygate4sd3_1 hold254 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][11] ),
    .X(net2851));
 sg13g2_dlygate4sd3_1 hold255 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][31] ),
    .X(net2852));
 sg13g2_dlygate4sd3_1 hold256 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][14] ),
    .X(net2853));
 sg13g2_dlygate4sd3_1 hold257 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[24] ),
    .X(net2854));
 sg13g2_dlygate4sd3_1 hold258 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][15] ),
    .X(net2855));
 sg13g2_dlygate4sd3_1 hold259 (.A(\soc_I.qqspi_I.rdata[29] ),
    .X(net2856));
 sg13g2_dlygate4sd3_1 hold260 (.A(_01825_),
    .X(net2857));
 sg13g2_dlygate4sd3_1 hold261 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][7] ),
    .X(net2858));
 sg13g2_dlygate4sd3_1 hold262 (.A(\soc_I.qqspi_I.rdata[0] ),
    .X(net2859));
 sg13g2_dlygate4sd3_1 hold263 (.A(_01796_),
    .X(net2860));
 sg13g2_dlygate4sd3_1 hold264 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][9] ),
    .X(net2861));
 sg13g2_dlygate4sd3_1 hold265 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][9] ),
    .X(net2862));
 sg13g2_dlygate4sd3_1 hold266 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][14] ),
    .X(net2863));
 sg13g2_dlygate4sd3_1 hold267 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][10] ),
    .X(net2864));
 sg13g2_dlygate4sd3_1 hold268 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][12] ),
    .X(net2865));
 sg13g2_dlygate4sd3_1 hold269 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][17] ),
    .X(net2866));
 sg13g2_dlygate4sd3_1 hold270 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][8] ),
    .X(net2867));
 sg13g2_dlygate4sd3_1 hold271 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][2] ),
    .X(net2868));
 sg13g2_dlygate4sd3_1 hold272 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.bit_idx[1] ),
    .X(net2869));
 sg13g2_dlygate4sd3_1 hold273 (.A(_05632_),
    .X(net2870));
 sg13g2_dlygate4sd3_1 hold274 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][20] ),
    .X(net2871));
 sg13g2_dlygate4sd3_1 hold275 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][1] ),
    .X(net2872));
 sg13g2_dlygate4sd3_1 hold276 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][11] ),
    .X(net2873));
 sg13g2_dlygate4sd3_1 hold277 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][19] ),
    .X(net2874));
 sg13g2_dlygate4sd3_1 hold278 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][20] ),
    .X(net2875));
 sg13g2_dlygate4sd3_1 hold279 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][14] ),
    .X(net2876));
 sg13g2_dlygate4sd3_1 hold280 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][30] ),
    .X(net2877));
 sg13g2_dlygate4sd3_1 hold281 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][9] ),
    .X(net2878));
 sg13g2_dlygate4sd3_1 hold282 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][12] ),
    .X(net2879));
 sg13g2_dlygate4sd3_1 hold283 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][23] ),
    .X(net2880));
 sg13g2_dlygate4sd3_1 hold284 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][5] ),
    .X(net2881));
 sg13g2_dlygate4sd3_1 hold285 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][1] ),
    .X(net2882));
 sg13g2_dlygate4sd3_1 hold286 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][25] ),
    .X(net2883));
 sg13g2_dlygate4sd3_1 hold287 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][26] ),
    .X(net2884));
 sg13g2_dlygate4sd3_1 hold288 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][17] ),
    .X(net2885));
 sg13g2_dlygate4sd3_1 hold289 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][10] ),
    .X(net2886));
 sg13g2_dlygate4sd3_1 hold290 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][11] ),
    .X(net2887));
 sg13g2_dlygate4sd3_1 hold291 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][12] ),
    .X(net2888));
 sg13g2_dlygate4sd3_1 hold292 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][17] ),
    .X(net2889));
 sg13g2_dlygate4sd3_1 hold293 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][31] ),
    .X(net2890));
 sg13g2_dlygate4sd3_1 hold294 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][19] ),
    .X(net2891));
 sg13g2_dlygate4sd3_1 hold295 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][26] ),
    .X(net2892));
 sg13g2_dlygate4sd3_1 hold296 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][18] ),
    .X(net2893));
 sg13g2_dlygate4sd3_1 hold297 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][7] ),
    .X(net2894));
 sg13g2_dlygate4sd3_1 hold298 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][15] ),
    .X(net2895));
 sg13g2_dlygate4sd3_1 hold299 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][20] ),
    .X(net2896));
 sg13g2_dlygate4sd3_1 hold300 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][17] ),
    .X(net2897));
 sg13g2_dlygate4sd3_1 hold301 (.A(_02730_),
    .X(net2898));
 sg13g2_dlygate4sd3_1 hold302 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][13] ),
    .X(net2899));
 sg13g2_dlygate4sd3_1 hold303 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][22] ),
    .X(net2900));
 sg13g2_dlygate4sd3_1 hold304 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[13] ),
    .X(net2901));
 sg13g2_dlygate4sd3_1 hold305 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][2] ),
    .X(net2902));
 sg13g2_dlygate4sd3_1 hold306 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][31] ),
    .X(net2903));
 sg13g2_dlygate4sd3_1 hold307 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][20] ),
    .X(net2904));
 sg13g2_dlygate4sd3_1 hold308 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][10] ),
    .X(net2905));
 sg13g2_dlygate4sd3_1 hold309 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][1] ),
    .X(net2906));
 sg13g2_dlygate4sd3_1 hold310 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][8] ),
    .X(net2907));
 sg13g2_dlygate4sd3_1 hold311 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][21] ),
    .X(net2908));
 sg13g2_dlygate4sd3_1 hold312 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][18] ),
    .X(net2909));
 sg13g2_dlygate4sd3_1 hold313 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][0] ),
    .X(net2910));
 sg13g2_dlygate4sd3_1 hold314 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][6] ),
    .X(net2911));
 sg13g2_dlygate4sd3_1 hold315 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][24] ),
    .X(net2912));
 sg13g2_dlygate4sd3_1 hold316 (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[8] ),
    .X(net2913));
 sg13g2_dlygate4sd3_1 hold317 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][31] ),
    .X(net2914));
 sg13g2_dlygate4sd3_1 hold318 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][1] ),
    .X(net2915));
 sg13g2_dlygate4sd3_1 hold319 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][3] ),
    .X(net2916));
 sg13g2_dlygate4sd3_1 hold320 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][6] ),
    .X(net2917));
 sg13g2_dlygate4sd3_1 hold321 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][28] ),
    .X(net2918));
 sg13g2_dlygate4sd3_1 hold322 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][5] ),
    .X(net2919));
 sg13g2_dlygate4sd3_1 hold323 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][22] ),
    .X(net2920));
 sg13g2_dlygate4sd3_1 hold324 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][21] ),
    .X(net2921));
 sg13g2_dlygate4sd3_1 hold325 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][18] ),
    .X(net2922));
 sg13g2_dlygate4sd3_1 hold326 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][2] ),
    .X(net2923));
 sg13g2_dlygate4sd3_1 hold327 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][30] ),
    .X(net2924));
 sg13g2_dlygate4sd3_1 hold328 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][29] ),
    .X(net2925));
 sg13g2_dlygate4sd3_1 hold329 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][22] ),
    .X(net2926));
 sg13g2_dlygate4sd3_1 hold330 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][16] ),
    .X(net2927));
 sg13g2_dlygate4sd3_1 hold331 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][7] ),
    .X(net2928));
 sg13g2_dlygate4sd3_1 hold332 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][19] ),
    .X(net2929));
 sg13g2_dlygate4sd3_1 hold333 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][12] ),
    .X(net2930));
 sg13g2_dlygate4sd3_1 hold334 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][10] ),
    .X(net2931));
 sg13g2_dlygate4sd3_1 hold335 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][29] ),
    .X(net2932));
 sg13g2_dlygate4sd3_1 hold336 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][17] ),
    .X(net2933));
 sg13g2_dlygate4sd3_1 hold337 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][0] ),
    .X(net2934));
 sg13g2_dlygate4sd3_1 hold338 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][22] ),
    .X(net2935));
 sg13g2_dlygate4sd3_1 hold339 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][6] ),
    .X(net2936));
 sg13g2_dlygate4sd3_1 hold340 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][20] ),
    .X(net2937));
 sg13g2_dlygate4sd3_1 hold341 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][26] ),
    .X(net2938));
 sg13g2_dlygate4sd3_1 hold342 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][12] ),
    .X(net2939));
 sg13g2_dlygate4sd3_1 hold343 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][1] ),
    .X(net2940));
 sg13g2_dlygate4sd3_1 hold344 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][12] ),
    .X(net2941));
 sg13g2_dlygate4sd3_1 hold345 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][9] ),
    .X(net2942));
 sg13g2_dlygate4sd3_1 hold346 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][16] ),
    .X(net2943));
 sg13g2_dlygate4sd3_1 hold347 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][9] ),
    .X(net2944));
 sg13g2_dlygate4sd3_1 hold348 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][28] ),
    .X(net2945));
 sg13g2_dlygate4sd3_1 hold349 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][13] ),
    .X(net2946));
 sg13g2_dlygate4sd3_1 hold350 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][0] ),
    .X(net2947));
 sg13g2_dlygate4sd3_1 hold351 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][3] ),
    .X(net2948));
 sg13g2_dlygate4sd3_1 hold352 (.A(\soc_I.qqspi_I.rdata[7] ),
    .X(net2949));
 sg13g2_dlygate4sd3_1 hold353 (.A(_01803_),
    .X(net2950));
 sg13g2_dlygate4sd3_1 hold354 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][17] ),
    .X(net2951));
 sg13g2_dlygate4sd3_1 hold355 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][17] ),
    .X(net2952));
 sg13g2_dlygate4sd3_1 hold356 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][18] ),
    .X(net2953));
 sg13g2_dlygate4sd3_1 hold357 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][10] ),
    .X(net2954));
 sg13g2_dlygate4sd3_1 hold358 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][2] ),
    .X(net2955));
 sg13g2_dlygate4sd3_1 hold359 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][11] ),
    .X(net2956));
 sg13g2_dlygate4sd3_1 hold360 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][2] ),
    .X(net2957));
 sg13g2_dlygate4sd3_1 hold361 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][24] ),
    .X(net2958));
 sg13g2_dlygate4sd3_1 hold362 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][4] ),
    .X(net2959));
 sg13g2_dlygate4sd3_1 hold363 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][28] ),
    .X(net2960));
 sg13g2_dlygate4sd3_1 hold364 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][8] ),
    .X(net2961));
 sg13g2_dlygate4sd3_1 hold365 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][0] ),
    .X(net2962));
 sg13g2_dlygate4sd3_1 hold366 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][5] ),
    .X(net2963));
 sg13g2_dlygate4sd3_1 hold367 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][5] ),
    .X(net2964));
 sg13g2_dlygate4sd3_1 hold368 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][27] ),
    .X(net2965));
 sg13g2_dlygate4sd3_1 hold369 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][15] ),
    .X(net2966));
 sg13g2_dlygate4sd3_1 hold370 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][0] ),
    .X(net2967));
 sg13g2_dlygate4sd3_1 hold371 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][1] ),
    .X(net2968));
 sg13g2_dlygate4sd3_1 hold372 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][2] ),
    .X(net2969));
 sg13g2_dlygate4sd3_1 hold373 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][3] ),
    .X(net2970));
 sg13g2_dlygate4sd3_1 hold374 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][10] ),
    .X(net2971));
 sg13g2_dlygate4sd3_1 hold375 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][8] ),
    .X(net2972));
 sg13g2_dlygate4sd3_1 hold376 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][10] ),
    .X(net2973));
 sg13g2_dlygate4sd3_1 hold377 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][17] ),
    .X(net2974));
 sg13g2_dlygate4sd3_1 hold378 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][1] ),
    .X(net2975));
 sg13g2_dlygate4sd3_1 hold379 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][28] ),
    .X(net2976));
 sg13g2_dlygate4sd3_1 hold380 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][17] ),
    .X(net2977));
 sg13g2_dlygate4sd3_1 hold381 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][9] ),
    .X(net2978));
 sg13g2_dlygate4sd3_1 hold382 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][22] ),
    .X(net2979));
 sg13g2_dlygate4sd3_1 hold383 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][10] ),
    .X(net2980));
 sg13g2_dlygate4sd3_1 hold384 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][9] ),
    .X(net2981));
 sg13g2_dlygate4sd3_1 hold385 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][5] ),
    .X(net2982));
 sg13g2_dlygate4sd3_1 hold386 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][2] ),
    .X(net2983));
 sg13g2_dlygate4sd3_1 hold387 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][10] ),
    .X(net2984));
 sg13g2_dlygate4sd3_1 hold388 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][10] ),
    .X(net2985));
 sg13g2_dlygate4sd3_1 hold389 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][9] ),
    .X(net2986));
 sg13g2_dlygate4sd3_1 hold390 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][21] ),
    .X(net2987));
 sg13g2_dlygate4sd3_1 hold391 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][19] ),
    .X(net2988));
 sg13g2_dlygate4sd3_1 hold392 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][16] ),
    .X(net2989));
 sg13g2_dlygate4sd3_1 hold393 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][6] ),
    .X(net2990));
 sg13g2_dlygate4sd3_1 hold394 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][28] ),
    .X(net2991));
 sg13g2_dlygate4sd3_1 hold395 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][15] ),
    .X(net2992));
 sg13g2_dlygate4sd3_1 hold396 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][23] ),
    .X(net2993));
 sg13g2_dlygate4sd3_1 hold397 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][6] ),
    .X(net2994));
 sg13g2_dlygate4sd3_1 hold398 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][9] ),
    .X(net2995));
 sg13g2_dlygate4sd3_1 hold399 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][0] ),
    .X(net2996));
 sg13g2_dlygate4sd3_1 hold400 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][21] ),
    .X(net2997));
 sg13g2_dlygate4sd3_1 hold401 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][25] ),
    .X(net2998));
 sg13g2_dlygate4sd3_1 hold402 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][29] ),
    .X(net2999));
 sg13g2_dlygate4sd3_1 hold403 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][10] ),
    .X(net3000));
 sg13g2_dlygate4sd3_1 hold404 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][11] ),
    .X(net3001));
 sg13g2_dlygate4sd3_1 hold405 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][31] ),
    .X(net3002));
 sg13g2_dlygate4sd3_1 hold406 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][22] ),
    .X(net3003));
 sg13g2_dlygate4sd3_1 hold407 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][9] ),
    .X(net3004));
 sg13g2_dlygate4sd3_1 hold408 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][10] ),
    .X(net3005));
 sg13g2_dlygate4sd3_1 hold409 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][2] ),
    .X(net3006));
 sg13g2_dlygate4sd3_1 hold410 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][20] ),
    .X(net3007));
 sg13g2_dlygate4sd3_1 hold411 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][2] ),
    .X(net3008));
 sg13g2_dlygate4sd3_1 hold412 (.A(\soc_I.rx_uart_i.return_state[1] ),
    .X(net3009));
 sg13g2_dlygate4sd3_1 hold413 (.A(_02139_),
    .X(net3010));
 sg13g2_dlygate4sd3_1 hold414 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][13] ),
    .X(net3011));
 sg13g2_dlygate4sd3_1 hold415 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][15] ),
    .X(net3012));
 sg13g2_dlygate4sd3_1 hold416 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][24] ),
    .X(net3013));
 sg13g2_dlygate4sd3_1 hold417 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][22] ),
    .X(net3014));
 sg13g2_dlygate4sd3_1 hold418 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][17] ),
    .X(net3015));
 sg13g2_dlygate4sd3_1 hold419 (.A(\soc_I.tx_uart_i.wait_states[8] ),
    .X(net3016));
 sg13g2_dlygate4sd3_1 hold420 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][22] ),
    .X(net3017));
 sg13g2_dlygate4sd3_1 hold421 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][10] ),
    .X(net3018));
 sg13g2_dlygate4sd3_1 hold422 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][29] ),
    .X(net3019));
 sg13g2_dlygate4sd3_1 hold423 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][13] ),
    .X(net3020));
 sg13g2_dlygate4sd3_1 hold424 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][16] ),
    .X(net3021));
 sg13g2_dlygate4sd3_1 hold425 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][2] ),
    .X(net3022));
 sg13g2_dlygate4sd3_1 hold426 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][26] ),
    .X(net3023));
 sg13g2_dlygate4sd3_1 hold427 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][23] ),
    .X(net3024));
 sg13g2_dlygate4sd3_1 hold428 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][9] ),
    .X(net3025));
 sg13g2_dlygate4sd3_1 hold429 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][6] ),
    .X(net3026));
 sg13g2_dlygate4sd3_1 hold430 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][26] ),
    .X(net3027));
 sg13g2_dlygate4sd3_1 hold431 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][3] ),
    .X(net3028));
 sg13g2_dlygate4sd3_1 hold432 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][29] ),
    .X(net3029));
 sg13g2_dlygate4sd3_1 hold433 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][29] ),
    .X(net3030));
 sg13g2_dlygate4sd3_1 hold434 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][25] ),
    .X(net3031));
 sg13g2_dlygate4sd3_1 hold435 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][16] ),
    .X(net3032));
 sg13g2_dlygate4sd3_1 hold436 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][10] ),
    .X(net3033));
 sg13g2_dlygate4sd3_1 hold437 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][19] ),
    .X(net3034));
 sg13g2_dlygate4sd3_1 hold438 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][27] ),
    .X(net3035));
 sg13g2_dlygate4sd3_1 hold439 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][19] ),
    .X(net3036));
 sg13g2_dlygate4sd3_1 hold440 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[0] ),
    .X(net3037));
 sg13g2_dlygate4sd3_1 hold441 (.A(_04425_),
    .X(net3038));
 sg13g2_dlygate4sd3_1 hold442 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][7] ),
    .X(net3039));
 sg13g2_dlygate4sd3_1 hold443 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][20] ),
    .X(net3040));
 sg13g2_dlygate4sd3_1 hold444 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][29] ),
    .X(net3041));
 sg13g2_dlygate4sd3_1 hold445 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][18] ),
    .X(net3042));
 sg13g2_dlygate4sd3_1 hold446 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][8] ),
    .X(net3043));
 sg13g2_dlygate4sd3_1 hold447 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][11] ),
    .X(net3044));
 sg13g2_dlygate4sd3_1 hold448 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][0] ),
    .X(net3045));
 sg13g2_dlygate4sd3_1 hold449 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][10] ),
    .X(net3046));
 sg13g2_dlygate4sd3_1 hold450 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][20] ),
    .X(net3047));
 sg13g2_dlygate4sd3_1 hold451 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][8] ),
    .X(net3048));
 sg13g2_dlygate4sd3_1 hold452 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][9] ),
    .X(net3049));
 sg13g2_dlygate4sd3_1 hold453 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][31] ),
    .X(net3050));
 sg13g2_dlygate4sd3_1 hold454 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][3] ),
    .X(net3051));
 sg13g2_dlygate4sd3_1 hold455 (.A(_00011_),
    .X(net3052));
 sg13g2_dlygate4sd3_1 hold456 (.A(_01984_),
    .X(net3053));
 sg13g2_dlygate4sd3_1 hold457 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][22] ),
    .X(net3054));
 sg13g2_dlygate4sd3_1 hold458 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][0] ),
    .X(net3055));
 sg13g2_dlygate4sd3_1 hold459 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][16] ),
    .X(net3056));
 sg13g2_dlygate4sd3_1 hold460 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][8] ),
    .X(net3057));
 sg13g2_dlygate4sd3_1 hold461 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][26] ),
    .X(net3058));
 sg13g2_dlygate4sd3_1 hold462 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][30] ),
    .X(net3059));
 sg13g2_dlygate4sd3_1 hold463 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][29] ),
    .X(net3060));
 sg13g2_dlygate4sd3_1 hold464 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][0] ),
    .X(net3061));
 sg13g2_dlygate4sd3_1 hold465 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][5] ),
    .X(net3062));
 sg13g2_dlygate4sd3_1 hold466 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][31] ),
    .X(net3063));
 sg13g2_dlygate4sd3_1 hold467 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][8] ),
    .X(net3064));
 sg13g2_dlygate4sd3_1 hold468 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][5] ),
    .X(net3065));
 sg13g2_dlygate4sd3_1 hold469 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][4] ),
    .X(net3066));
 sg13g2_dlygate4sd3_1 hold470 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][9] ),
    .X(net3067));
 sg13g2_dlygate4sd3_1 hold471 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][6] ),
    .X(net3068));
 sg13g2_dlygate4sd3_1 hold472 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][7] ),
    .X(net3069));
 sg13g2_dlygate4sd3_1 hold473 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][6] ),
    .X(net3070));
 sg13g2_dlygate4sd3_1 hold474 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][25] ),
    .X(net3071));
 sg13g2_dlygate4sd3_1 hold475 (.A(sio3_o),
    .X(net3072));
 sg13g2_dlygate4sd3_1 hold476 (.A(_07300_),
    .X(net3073));
 sg13g2_dlygate4sd3_1 hold477 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][9] ),
    .X(net3074));
 sg13g2_dlygate4sd3_1 hold478 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][15] ),
    .X(net3075));
 sg13g2_dlygate4sd3_1 hold479 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][22] ),
    .X(net3076));
 sg13g2_dlygate4sd3_1 hold480 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][31] ),
    .X(net3077));
 sg13g2_dlygate4sd3_1 hold481 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][21] ),
    .X(net3078));
 sg13g2_dlygate4sd3_1 hold482 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][24] ),
    .X(net3079));
 sg13g2_dlygate4sd3_1 hold483 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][21] ),
    .X(net3080));
 sg13g2_dlygate4sd3_1 hold484 (.A(_01913_),
    .X(net3081));
 sg13g2_dlygate4sd3_1 hold485 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][22] ),
    .X(net3082));
 sg13g2_dlygate4sd3_1 hold486 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][17] ),
    .X(net3083));
 sg13g2_dlygate4sd3_1 hold487 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][25] ),
    .X(net3084));
 sg13g2_dlygate4sd3_1 hold488 (.A(\soc_I.qqspi_I.rdata[22] ),
    .X(net3085));
 sg13g2_dlygate4sd3_1 hold489 (.A(_01818_),
    .X(net3086));
 sg13g2_dlygate4sd3_1 hold490 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][16] ),
    .X(net3087));
 sg13g2_dlygate4sd3_1 hold491 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][30] ),
    .X(net3088));
 sg13g2_dlygate4sd3_1 hold492 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][17] ),
    .X(net3089));
 sg13g2_dlygate4sd3_1 hold493 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][3] ),
    .X(net3090));
 sg13g2_dlygate4sd3_1 hold494 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][31] ),
    .X(net3091));
 sg13g2_dlygate4sd3_1 hold495 (.A(\soc_I.qqspi_I.rdata[24] ),
    .X(net3092));
 sg13g2_dlygate4sd3_1 hold496 (.A(_01820_),
    .X(net3093));
 sg13g2_dlygate4sd3_1 hold497 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][7] ),
    .X(net3094));
 sg13g2_dlygate4sd3_1 hold498 (.A(_00300_),
    .X(net3095));
 sg13g2_dlygate4sd3_1 hold499 (.A(_01839_),
    .X(net3096));
 sg13g2_dlygate4sd3_1 hold500 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][14] ),
    .X(net3097));
 sg13g2_dlygate4sd3_1 hold501 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[10] ),
    .X(net3098));
 sg13g2_dlygate4sd3_1 hold502 (.A(_01147_),
    .X(net3099));
 sg13g2_dlygate4sd3_1 hold503 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][18] ),
    .X(net3100));
 sg13g2_dlygate4sd3_1 hold504 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][3] ),
    .X(net3101));
 sg13g2_dlygate4sd3_1 hold505 (.A(sio2_o),
    .X(net3102));
 sg13g2_dlygate4sd3_1 hold506 (.A(_07299_),
    .X(net3103));
 sg13g2_dlygate4sd3_1 hold507 (.A(\soc_I.qqspi_I.state[4] ),
    .X(net3104));
 sg13g2_dlygate4sd3_1 hold508 (.A(_12569_),
    .X(net3105));
 sg13g2_dlygate4sd3_1 hold509 (.A(_00008_),
    .X(net3106));
 sg13g2_dlygate4sd3_1 hold510 (.A(\soc_I.tx_uart_i.wait_states[7] ),
    .X(net3107));
 sg13g2_dlygate4sd3_1 hold511 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][21] ),
    .X(net3108));
 sg13g2_dlygate4sd3_1 hold512 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][6] ),
    .X(net3109));
 sg13g2_dlygate4sd3_1 hold513 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][27] ),
    .X(net3110));
 sg13g2_dlygate4sd3_1 hold514 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][5] ),
    .X(net3111));
 sg13g2_dlygate4sd3_1 hold515 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][16] ),
    .X(net3112));
 sg13g2_dlygate4sd3_1 hold516 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][22] ),
    .X(net3113));
 sg13g2_dlygate4sd3_1 hold517 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][0] ),
    .X(net3114));
 sg13g2_dlygate4sd3_1 hold518 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][29] ),
    .X(net3115));
 sg13g2_dlygate4sd3_1 hold519 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][30] ),
    .X(net3116));
 sg13g2_dlygate4sd3_1 hold520 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][21] ),
    .X(net3117));
 sg13g2_dlygate4sd3_1 hold521 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][21] ),
    .X(net3118));
 sg13g2_dlygate4sd3_1 hold522 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][1] ),
    .X(net3119));
 sg13g2_dlygate4sd3_1 hold523 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][9] ),
    .X(net3120));
 sg13g2_dlygate4sd3_1 hold524 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][11] ),
    .X(net3121));
 sg13g2_dlygate4sd3_1 hold525 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][0] ),
    .X(net3122));
 sg13g2_dlygate4sd3_1 hold526 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][25] ),
    .X(net3123));
 sg13g2_dlygate4sd3_1 hold527 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][19] ),
    .X(net3124));
 sg13g2_dlygate4sd3_1 hold528 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][24] ),
    .X(net3125));
 sg13g2_dlygate4sd3_1 hold529 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][30] ),
    .X(net3126));
 sg13g2_dlygate4sd3_1 hold530 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][8] ),
    .X(net3127));
 sg13g2_dlygate4sd3_1 hold531 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][4] ),
    .X(net3128));
 sg13g2_dlygate4sd3_1 hold532 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][28] ),
    .X(net3129));
 sg13g2_dlygate4sd3_1 hold533 (.A(\soc_I.rx_uart_i.fifo_i.ram[13][4] ),
    .X(net3130));
 sg13g2_dlygate4sd3_1 hold534 (.A(_00666_),
    .X(net3131));
 sg13g2_dlygate4sd3_1 hold535 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][19] ),
    .X(net3132));
 sg13g2_dlygate4sd3_1 hold536 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][18] ),
    .X(net3133));
 sg13g2_dlygate4sd3_1 hold537 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][5] ),
    .X(net3134));
 sg13g2_dlygate4sd3_1 hold538 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][10] ),
    .X(net3135));
 sg13g2_dlygate4sd3_1 hold539 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][25] ),
    .X(net3136));
 sg13g2_dlygate4sd3_1 hold540 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][29] ),
    .X(net3137));
 sg13g2_dlygate4sd3_1 hold541 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][1] ),
    .X(net3138));
 sg13g2_dlygate4sd3_1 hold542 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][29] ),
    .X(net3139));
 sg13g2_dlygate4sd3_1 hold543 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][5] ),
    .X(net3140));
 sg13g2_dlygate4sd3_1 hold544 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][7] ),
    .X(net3141));
 sg13g2_dlygate4sd3_1 hold545 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][3] ),
    .X(net3142));
 sg13g2_dlygate4sd3_1 hold546 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][25] ),
    .X(net3143));
 sg13g2_dlygate4sd3_1 hold547 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][15] ),
    .X(net3144));
 sg13g2_dlygate4sd3_1 hold548 (.A(\soc_I.qqspi_I.rdata[13] ),
    .X(net3145));
 sg13g2_dlygate4sd3_1 hold549 (.A(_01809_),
    .X(net3146));
 sg13g2_dlygate4sd3_1 hold550 (.A(\soc_I.rx_uart_i.fifo_i.rd_ptr[3] ),
    .X(net3147));
 sg13g2_dlygate4sd3_1 hold551 (.A(_02780_),
    .X(net3148));
 sg13g2_dlygate4sd3_1 hold552 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][30] ),
    .X(net3149));
 sg13g2_dlygate4sd3_1 hold553 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][6] ),
    .X(net3150));
 sg13g2_dlygate4sd3_1 hold554 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][27] ),
    .X(net3151));
 sg13g2_dlygate4sd3_1 hold555 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][27] ),
    .X(net3152));
 sg13g2_dlygate4sd3_1 hold556 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][13] ),
    .X(net3153));
 sg13g2_dlygate4sd3_1 hold557 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][25] ),
    .X(net3154));
 sg13g2_dlygate4sd3_1 hold558 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][14] ),
    .X(net3155));
 sg13g2_dlygate4sd3_1 hold559 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][10] ),
    .X(net3156));
 sg13g2_dlygate4sd3_1 hold560 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][1] ),
    .X(net3157));
 sg13g2_dlygate4sd3_1 hold561 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][2] ),
    .X(net3158));
 sg13g2_dlygate4sd3_1 hold562 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][13] ),
    .X(net3159));
 sg13g2_dlygate4sd3_1 hold563 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][24] ),
    .X(net3160));
 sg13g2_dlygate4sd3_1 hold564 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][26] ),
    .X(net3161));
 sg13g2_dlygate4sd3_1 hold565 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][5] ),
    .X(net3162));
 sg13g2_dlygate4sd3_1 hold566 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][9] ),
    .X(net3163));
 sg13g2_dlygate4sd3_1 hold567 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][6] ),
    .X(net3164));
 sg13g2_dlygate4sd3_1 hold568 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][13] ),
    .X(net3165));
 sg13g2_dlygate4sd3_1 hold569 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][10] ),
    .X(net3166));
 sg13g2_dlygate4sd3_1 hold570 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][10] ),
    .X(net3167));
 sg13g2_dlygate4sd3_1 hold571 (.A(\soc_I.rx_uart_i.fifo_i.ram[13][7] ),
    .X(net3168));
 sg13g2_dlygate4sd3_1 hold572 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][19] ),
    .X(net3169));
 sg13g2_dlygate4sd3_1 hold573 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][14] ),
    .X(net3170));
 sg13g2_dlygate4sd3_1 hold574 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][23] ),
    .X(net3171));
 sg13g2_dlygate4sd3_1 hold575 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][9] ),
    .X(net3172));
 sg13g2_dlygate4sd3_1 hold576 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][30] ),
    .X(net3173));
 sg13g2_dlygate4sd3_1 hold577 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][29] ),
    .X(net3174));
 sg13g2_dlygate4sd3_1 hold578 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][31] ),
    .X(net3175));
 sg13g2_dlygate4sd3_1 hold579 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][15] ),
    .X(net3176));
 sg13g2_dlygate4sd3_1 hold580 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][13] ),
    .X(net3177));
 sg13g2_dlygate4sd3_1 hold581 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][3] ),
    .X(net3178));
 sg13g2_dlygate4sd3_1 hold582 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][28] ),
    .X(net3179));
 sg13g2_dlygate4sd3_1 hold583 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][21] ),
    .X(net3180));
 sg13g2_dlygate4sd3_1 hold584 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][0] ),
    .X(net3181));
 sg13g2_dlygate4sd3_1 hold585 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][28] ),
    .X(net3182));
 sg13g2_dlygate4sd3_1 hold586 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][6] ),
    .X(net3183));
 sg13g2_dlygate4sd3_1 hold587 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][30] ),
    .X(net3184));
 sg13g2_dlygate4sd3_1 hold588 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][3] ),
    .X(net3185));
 sg13g2_dlygate4sd3_1 hold589 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][26] ),
    .X(net3186));
 sg13g2_dlygate4sd3_1 hold590 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][6] ),
    .X(net3187));
 sg13g2_dlygate4sd3_1 hold591 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][23] ),
    .X(net3188));
 sg13g2_dlygate4sd3_1 hold592 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][23] ),
    .X(net3189));
 sg13g2_dlygate4sd3_1 hold593 (.A(\soc_I.spi0_I.xfer_cycles[3] ),
    .X(net3190));
 sg13g2_dlygate4sd3_1 hold594 (.A(_01749_),
    .X(net3191));
 sg13g2_dlygate4sd3_1 hold595 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][14] ),
    .X(net3192));
 sg13g2_dlygate4sd3_1 hold596 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[62] ),
    .X(net3193));
 sg13g2_dlygate4sd3_1 hold597 (.A(_01199_),
    .X(net3194));
 sg13g2_dlygate4sd3_1 hold598 (.A(\soc_I.rx_uart_i.fifo_i.ram[13][2] ),
    .X(net3195));
 sg13g2_dlygate4sd3_1 hold599 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][16] ),
    .X(net3196));
 sg13g2_dlygate4sd3_1 hold600 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][22] ),
    .X(net3197));
 sg13g2_dlygate4sd3_1 hold601 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][0] ),
    .X(net3198));
 sg13g2_dlygate4sd3_1 hold602 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][2] ),
    .X(net3199));
 sg13g2_dlygate4sd3_1 hold603 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][3] ),
    .X(net3200));
 sg13g2_dlygate4sd3_1 hold604 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][22] ),
    .X(net3201));
 sg13g2_dlygate4sd3_1 hold605 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][23] ),
    .X(net3202));
 sg13g2_dlygate4sd3_1 hold606 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][0] ),
    .X(net3203));
 sg13g2_dlygate4sd3_1 hold607 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][10] ),
    .X(net3204));
 sg13g2_dlygate4sd3_1 hold608 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[58] ),
    .X(net3205));
 sg13g2_dlygate4sd3_1 hold609 (.A(_05618_),
    .X(net3206));
 sg13g2_dlygate4sd3_1 hold610 (.A(_01323_),
    .X(net3207));
 sg13g2_dlygate4sd3_1 hold611 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][13] ),
    .X(net3208));
 sg13g2_dlygate4sd3_1 hold612 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][17] ),
    .X(net3209));
 sg13g2_dlygate4sd3_1 hold613 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][23] ),
    .X(net3210));
 sg13g2_dlygate4sd3_1 hold614 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][1] ),
    .X(net3211));
 sg13g2_dlygate4sd3_1 hold615 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][0] ),
    .X(net3212));
 sg13g2_dlygate4sd3_1 hold616 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][22] ),
    .X(net3213));
 sg13g2_dlygate4sd3_1 hold617 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][8] ),
    .X(net3214));
 sg13g2_dlygate4sd3_1 hold618 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[10] ),
    .X(net3215));
 sg13g2_dlygate4sd3_1 hold619 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][31] ),
    .X(net3216));
 sg13g2_dlygate4sd3_1 hold620 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][26] ),
    .X(net3217));
 sg13g2_dlygate4sd3_1 hold621 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][30] ),
    .X(net3218));
 sg13g2_dlygate4sd3_1 hold622 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[14] ),
    .X(net3219));
 sg13g2_dlygate4sd3_1 hold623 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][29] ),
    .X(net3220));
 sg13g2_dlygate4sd3_1 hold624 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][31] ),
    .X(net3221));
 sg13g2_dlygate4sd3_1 hold625 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][1] ),
    .X(net3222));
 sg13g2_dlygate4sd3_1 hold626 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][18] ),
    .X(net3223));
 sg13g2_dlygate4sd3_1 hold627 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][18] ),
    .X(net3224));
 sg13g2_dlygate4sd3_1 hold628 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][5] ),
    .X(net3225));
 sg13g2_dlygate4sd3_1 hold629 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][11] ),
    .X(net3226));
 sg13g2_dlygate4sd3_1 hold630 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][13] ),
    .X(net3227));
 sg13g2_dlygate4sd3_1 hold631 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][22] ),
    .X(net3228));
 sg13g2_dlygate4sd3_1 hold632 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[5] ),
    .X(net3229));
 sg13g2_dlygate4sd3_1 hold633 (.A(_02203_),
    .X(net3230));
 sg13g2_dlygate4sd3_1 hold634 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][29] ),
    .X(net3231));
 sg13g2_dlygate4sd3_1 hold635 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][2] ),
    .X(net3232));
 sg13g2_dlygate4sd3_1 hold636 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][19] ),
    .X(net3233));
 sg13g2_dlygate4sd3_1 hold637 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][4] ),
    .X(net3234));
 sg13g2_dlygate4sd3_1 hold638 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][12] ),
    .X(net3235));
 sg13g2_dlygate4sd3_1 hold639 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[17] ),
    .X(net3236));
 sg13g2_dlygate4sd3_1 hold640 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][25] ),
    .X(net3237));
 sg13g2_dlygate4sd3_1 hold641 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][5] ),
    .X(net3238));
 sg13g2_dlygate4sd3_1 hold642 (.A(\soc_I.tx_uart_i.wait_states[3] ),
    .X(net3239));
 sg13g2_dlygate4sd3_1 hold643 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][2] ),
    .X(net3240));
 sg13g2_dlygate4sd3_1 hold644 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][5] ),
    .X(net3241));
 sg13g2_dlygate4sd3_1 hold645 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][24] ),
    .X(net3242));
 sg13g2_dlygate4sd3_1 hold646 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][9] ),
    .X(net3243));
 sg13g2_dlygate4sd3_1 hold647 (.A(\soc_I.tx_uart_i.wait_states[2] ),
    .X(net3244));
 sg13g2_dlygate4sd3_1 hold648 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][7] ),
    .X(net3245));
 sg13g2_dlygate4sd3_1 hold649 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][28] ),
    .X(net3246));
 sg13g2_dlygate4sd3_1 hold650 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][13] ),
    .X(net3247));
 sg13g2_dlygate4sd3_1 hold651 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][16] ),
    .X(net3248));
 sg13g2_dlygate4sd3_1 hold652 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][9] ),
    .X(net3249));
 sg13g2_dlygate4sd3_1 hold653 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][11] ),
    .X(net3250));
 sg13g2_dlygate4sd3_1 hold654 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][23] ),
    .X(net3251));
 sg13g2_dlygate4sd3_1 hold655 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][23] ),
    .X(net3252));
 sg13g2_dlygate4sd3_1 hold656 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][1] ),
    .X(net3253));
 sg13g2_dlygate4sd3_1 hold657 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[30] ),
    .X(net3254));
 sg13g2_dlygate4sd3_1 hold658 (.A(_05571_),
    .X(net3255));
 sg13g2_dlygate4sd3_1 hold659 (.A(_01295_),
    .X(net3256));
 sg13g2_dlygate4sd3_1 hold660 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][26] ),
    .X(net3257));
 sg13g2_dlygate4sd3_1 hold661 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][15] ),
    .X(net3258));
 sg13g2_dlygate4sd3_1 hold662 (.A(\soc_I.rx_uart_i.fifo_i.ram[14][3] ),
    .X(net3259));
 sg13g2_dlygate4sd3_1 hold663 (.A(_00673_),
    .X(net3260));
 sg13g2_dlygate4sd3_1 hold664 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][26] ),
    .X(net3261));
 sg13g2_dlygate4sd3_1 hold665 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][11] ),
    .X(net3262));
 sg13g2_dlygate4sd3_1 hold666 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][8] ),
    .X(net3263));
 sg13g2_dlygate4sd3_1 hold667 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][8] ),
    .X(net3264));
 sg13g2_dlygate4sd3_1 hold668 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][20] ),
    .X(net3265));
 sg13g2_dlygate4sd3_1 hold669 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][4] ),
    .X(net3266));
 sg13g2_dlygate4sd3_1 hold670 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][30] ),
    .X(net3267));
 sg13g2_dlygate4sd3_1 hold671 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][22] ),
    .X(net3268));
 sg13g2_dlygate4sd3_1 hold672 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][26] ),
    .X(net3269));
 sg13g2_dlygate4sd3_1 hold673 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][15] ),
    .X(net3270));
 sg13g2_dlygate4sd3_1 hold674 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][3] ),
    .X(net3271));
 sg13g2_dlygate4sd3_1 hold675 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][8] ),
    .X(net3272));
 sg13g2_dlygate4sd3_1 hold676 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][15] ),
    .X(net3273));
 sg13g2_dlygate4sd3_1 hold677 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][6] ),
    .X(net3274));
 sg13g2_dlygate4sd3_1 hold678 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][24] ),
    .X(net3275));
 sg13g2_dlygate4sd3_1 hold679 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][13] ),
    .X(net3276));
 sg13g2_dlygate4sd3_1 hold680 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][3] ),
    .X(net3277));
 sg13g2_dlygate4sd3_1 hold681 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][20] ),
    .X(net3278));
 sg13g2_dlygate4sd3_1 hold682 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][3] ),
    .X(net3279));
 sg13g2_dlygate4sd3_1 hold683 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][6] ),
    .X(net3280));
 sg13g2_dlygate4sd3_1 hold684 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][26] ),
    .X(net3281));
 sg13g2_dlygate4sd3_1 hold685 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][9] ),
    .X(net3282));
 sg13g2_dlygate4sd3_1 hold686 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][6] ),
    .X(net3283));
 sg13g2_dlygate4sd3_1 hold687 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][15] ),
    .X(net3284));
 sg13g2_dlygate4sd3_1 hold688 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][10] ),
    .X(net3285));
 sg13g2_dlygate4sd3_1 hold689 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][17] ),
    .X(net3286));
 sg13g2_dlygate4sd3_1 hold690 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][8] ),
    .X(net3287));
 sg13g2_dlygate4sd3_1 hold691 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][25] ),
    .X(net3288));
 sg13g2_dlygate4sd3_1 hold692 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][22] ),
    .X(net3289));
 sg13g2_dlygate4sd3_1 hold693 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][17] ),
    .X(net3290));
 sg13g2_dlygate4sd3_1 hold694 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][6] ),
    .X(net3291));
 sg13g2_dlygate4sd3_1 hold695 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][2] ),
    .X(net3292));
 sg13g2_dlygate4sd3_1 hold696 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][26] ),
    .X(net3293));
 sg13g2_dlygate4sd3_1 hold697 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][7] ),
    .X(net3294));
 sg13g2_dlygate4sd3_1 hold698 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][30] ),
    .X(net3295));
 sg13g2_dlygate4sd3_1 hold699 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][20] ),
    .X(net3296));
 sg13g2_dlygate4sd3_1 hold700 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][10] ),
    .X(net3297));
 sg13g2_dlygate4sd3_1 hold701 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][4] ),
    .X(net3298));
 sg13g2_dlygate4sd3_1 hold702 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][2] ),
    .X(net3299));
 sg13g2_dlygate4sd3_1 hold703 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][12] ),
    .X(net3300));
 sg13g2_dlygate4sd3_1 hold704 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][6] ),
    .X(net3301));
 sg13g2_dlygate4sd3_1 hold705 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][19] ),
    .X(net3302));
 sg13g2_dlygate4sd3_1 hold706 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][1] ),
    .X(net3303));
 sg13g2_dlygate4sd3_1 hold707 (.A(\soc_I.rx_uart_i.fifo_i.ram[14][6] ),
    .X(net3304));
 sg13g2_dlygate4sd3_1 hold708 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][6] ),
    .X(net3305));
 sg13g2_dlygate4sd3_1 hold709 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][20] ),
    .X(net3306));
 sg13g2_dlygate4sd3_1 hold710 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][26] ),
    .X(net3307));
 sg13g2_dlygate4sd3_1 hold711 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][9] ),
    .X(net3308));
 sg13g2_dlygate4sd3_1 hold712 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[46] ),
    .X(net3309));
 sg13g2_dlygate4sd3_1 hold713 (.A(_05598_),
    .X(net3310));
 sg13g2_dlygate4sd3_1 hold714 (.A(_01311_),
    .X(net3311));
 sg13g2_dlygate4sd3_1 hold715 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][6] ),
    .X(net3312));
 sg13g2_dlygate4sd3_1 hold716 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[2] ),
    .X(net3313));
 sg13g2_dlygate4sd3_1 hold717 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][5] ),
    .X(net3314));
 sg13g2_dlygate4sd3_1 hold718 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][12] ),
    .X(net3315));
 sg13g2_dlygate4sd3_1 hold719 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][22] ),
    .X(net3316));
 sg13g2_dlygate4sd3_1 hold720 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][4] ),
    .X(net3317));
 sg13g2_dlygate4sd3_1 hold721 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][4] ),
    .X(net3318));
 sg13g2_dlygate4sd3_1 hold722 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][15] ),
    .X(net3319));
 sg13g2_dlygate4sd3_1 hold723 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][14] ),
    .X(net3320));
 sg13g2_dlygate4sd3_1 hold724 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][24] ),
    .X(net3321));
 sg13g2_dlygate4sd3_1 hold725 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][27] ),
    .X(net3322));
 sg13g2_dlygate4sd3_1 hold726 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][27] ),
    .X(net3323));
 sg13g2_dlygate4sd3_1 hold727 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][0] ),
    .X(net3324));
 sg13g2_dlygate4sd3_1 hold728 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][25] ),
    .X(net3325));
 sg13g2_dlygate4sd3_1 hold729 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][16] ),
    .X(net3326));
 sg13g2_dlygate4sd3_1 hold730 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][13] ),
    .X(net3327));
 sg13g2_dlygate4sd3_1 hold731 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][1] ),
    .X(net3328));
 sg13g2_dlygate4sd3_1 hold732 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][0] ),
    .X(net3329));
 sg13g2_dlygate4sd3_1 hold733 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][29] ),
    .X(net3330));
 sg13g2_dlygate4sd3_1 hold734 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][16] ),
    .X(net3331));
 sg13g2_dlygate4sd3_1 hold735 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][14] ),
    .X(net3332));
 sg13g2_dlygate4sd3_1 hold736 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][0] ),
    .X(net3333));
 sg13g2_dlygate4sd3_1 hold737 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][21] ),
    .X(net3334));
 sg13g2_dlygate4sd3_1 hold738 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][2] ),
    .X(net3335));
 sg13g2_dlygate4sd3_1 hold739 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][6] ),
    .X(net3336));
 sg13g2_dlygate4sd3_1 hold740 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][31] ),
    .X(net3337));
 sg13g2_dlygate4sd3_1 hold741 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][31] ),
    .X(net3338));
 sg13g2_dlygate4sd3_1 hold742 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][24] ),
    .X(net3339));
 sg13g2_dlygate4sd3_1 hold743 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][1] ),
    .X(net3340));
 sg13g2_dlygate4sd3_1 hold744 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][24] ),
    .X(net3341));
 sg13g2_dlygate4sd3_1 hold745 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][28] ),
    .X(net3342));
 sg13g2_dlygate4sd3_1 hold746 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][5] ),
    .X(net3343));
 sg13g2_dlygate4sd3_1 hold747 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][27] ),
    .X(net3344));
 sg13g2_dlygate4sd3_1 hold748 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][3] ),
    .X(net3345));
 sg13g2_dlygate4sd3_1 hold749 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][28] ),
    .X(net3346));
 sg13g2_dlygate4sd3_1 hold750 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][15] ),
    .X(net3347));
 sg13g2_dlygate4sd3_1 hold751 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][24] ),
    .X(net3348));
 sg13g2_dlygate4sd3_1 hold752 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][9] ),
    .X(net3349));
 sg13g2_dlygate4sd3_1 hold753 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][3] ),
    .X(net3350));
 sg13g2_dlygate4sd3_1 hold754 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][6] ),
    .X(net3351));
 sg13g2_dlygate4sd3_1 hold755 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][7] ),
    .X(net3352));
 sg13g2_dlygate4sd3_1 hold756 (.A(\soc_I.rx_uart_i.fifo_i.ram[13][1] ),
    .X(net3353));
 sg13g2_dlygate4sd3_1 hold757 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][29] ),
    .X(net3354));
 sg13g2_dlygate4sd3_1 hold758 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][5] ),
    .X(net3355));
 sg13g2_dlygate4sd3_1 hold759 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][25] ),
    .X(net3356));
 sg13g2_dlygate4sd3_1 hold760 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[0][7] ),
    .X(net3357));
 sg13g2_dlygate4sd3_1 hold761 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][6] ),
    .X(net3358));
 sg13g2_dlygate4sd3_1 hold762 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][29] ),
    .X(net3359));
 sg13g2_dlygate4sd3_1 hold763 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][28] ),
    .X(net3360));
 sg13g2_dlygate4sd3_1 hold764 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][7] ),
    .X(net3361));
 sg13g2_dlygate4sd3_1 hold765 (.A(\soc_I.rx_uart_i.fifo_i.ram[13][6] ),
    .X(net3362));
 sg13g2_dlygate4sd3_1 hold766 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][20] ),
    .X(net3363));
 sg13g2_dlygate4sd3_1 hold767 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[10] ),
    .X(net3364));
 sg13g2_dlygate4sd3_1 hold768 (.A(_05538_),
    .X(net3365));
 sg13g2_dlygate4sd3_1 hold769 (.A(_01275_),
    .X(net3366));
 sg13g2_dlygate4sd3_1 hold770 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][26] ),
    .X(net3367));
 sg13g2_dlygate4sd3_1 hold771 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][16] ),
    .X(net3368));
 sg13g2_dlygate4sd3_1 hold772 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][0] ),
    .X(net3369));
 sg13g2_dlygate4sd3_1 hold773 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][16] ),
    .X(net3370));
 sg13g2_dlygate4sd3_1 hold774 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][13] ),
    .X(net3371));
 sg13g2_dlygate4sd3_1 hold775 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][23] ),
    .X(net3372));
 sg13g2_dlygate4sd3_1 hold776 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][20] ),
    .X(net3373));
 sg13g2_dlygate4sd3_1 hold777 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[16] ),
    .X(net3374));
 sg13g2_dlygate4sd3_1 hold778 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][8] ),
    .X(net3375));
 sg13g2_dlygate4sd3_1 hold779 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][15] ),
    .X(net3376));
 sg13g2_dlygate4sd3_1 hold780 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][18] ),
    .X(net3377));
 sg13g2_dlygate4sd3_1 hold781 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][7] ),
    .X(net3378));
 sg13g2_dlygate4sd3_1 hold782 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][30] ),
    .X(net3379));
 sg13g2_dlygate4sd3_1 hold783 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][4] ),
    .X(net3380));
 sg13g2_dlygate4sd3_1 hold784 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[3] ),
    .X(net3381));
 sg13g2_dlygate4sd3_1 hold785 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][28] ),
    .X(net3382));
 sg13g2_dlygate4sd3_1 hold786 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][19] ),
    .X(net3383));
 sg13g2_dlygate4sd3_1 hold787 (.A(\soc_I.rx_uart_i.fifo_i.ram[13][0] ),
    .X(net3384));
 sg13g2_dlygate4sd3_1 hold788 (.A(_00662_),
    .X(net3385));
 sg13g2_dlygate4sd3_1 hold789 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][30] ),
    .X(net3386));
 sg13g2_dlygate4sd3_1 hold790 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][13] ),
    .X(net3387));
 sg13g2_dlygate4sd3_1 hold791 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][16] ),
    .X(net3388));
 sg13g2_dlygate4sd3_1 hold792 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][26] ),
    .X(net3389));
 sg13g2_dlygate4sd3_1 hold793 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][20] ),
    .X(net3390));
 sg13g2_dlygate4sd3_1 hold794 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][10] ),
    .X(net3391));
 sg13g2_dlygate4sd3_1 hold795 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][7] ),
    .X(net3392));
 sg13g2_dlygate4sd3_1 hold796 (.A(\soc_I.rx_uart_i.fifo_i.ram[14][4] ),
    .X(net3393));
 sg13g2_dlygate4sd3_1 hold797 (.A(_00674_),
    .X(net3394));
 sg13g2_dlygate4sd3_1 hold798 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][5] ),
    .X(net3395));
 sg13g2_dlygate4sd3_1 hold799 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][22] ),
    .X(net3396));
 sg13g2_dlygate4sd3_1 hold800 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][13] ),
    .X(net3397));
 sg13g2_dlygate4sd3_1 hold801 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][13] ),
    .X(net3398));
 sg13g2_dlygate4sd3_1 hold802 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][20] ),
    .X(net3399));
 sg13g2_dlygate4sd3_1 hold803 (.A(\soc_I.rx_uart_i.state[2] ),
    .X(net3400));
 sg13g2_dlygate4sd3_1 hold804 (.A(_06696_),
    .X(net3401));
 sg13g2_dlygate4sd3_1 hold805 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][20] ),
    .X(net3402));
 sg13g2_dlygate4sd3_1 hold806 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][29] ),
    .X(net3403));
 sg13g2_dlygate4sd3_1 hold807 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][6] ),
    .X(net3404));
 sg13g2_dlygate4sd3_1 hold808 (.A(\gpio_uo_out[1] ),
    .X(net3405));
 sg13g2_dlygate4sd3_1 hold809 (.A(_01788_),
    .X(net3406));
 sg13g2_dlygate4sd3_1 hold810 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][5] ),
    .X(net3407));
 sg13g2_dlygate4sd3_1 hold811 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][20] ),
    .X(net3408));
 sg13g2_dlygate4sd3_1 hold812 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][31] ),
    .X(net3409));
 sg13g2_dlygate4sd3_1 hold813 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][16] ),
    .X(net3410));
 sg13g2_dlygate4sd3_1 hold814 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][12] ),
    .X(net3411));
 sg13g2_dlygate4sd3_1 hold815 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][5] ),
    .X(net3412));
 sg13g2_dlygate4sd3_1 hold816 (.A(\soc_I.clint_I.mtime[7] ),
    .X(net3413));
 sg13g2_dlygate4sd3_1 hold817 (.A(_01639_),
    .X(net3414));
 sg13g2_dlygate4sd3_1 hold818 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][19] ),
    .X(net3415));
 sg13g2_dlygate4sd3_1 hold819 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][30] ),
    .X(net3416));
 sg13g2_dlygate4sd3_1 hold820 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][7] ),
    .X(net3417));
 sg13g2_dlygate4sd3_1 hold821 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][19] ),
    .X(net3418));
 sg13g2_dlygate4sd3_1 hold822 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[16] ),
    .X(net3419));
 sg13g2_dlygate4sd3_1 hold823 (.A(_05548_),
    .X(net3420));
 sg13g2_dlygate4sd3_1 hold824 (.A(_01281_),
    .X(net3421));
 sg13g2_dlygate4sd3_1 hold825 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][19] ),
    .X(net3422));
 sg13g2_dlygate4sd3_1 hold826 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][24] ),
    .X(net3423));
 sg13g2_dlygate4sd3_1 hold827 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][15] ),
    .X(net3424));
 sg13g2_dlygate4sd3_1 hold828 (.A(\soc_I.spi0_I.tick_cnt[6] ),
    .X(net3425));
 sg13g2_dlygate4sd3_1 hold829 (.A(_06621_),
    .X(net3426));
 sg13g2_dlygate4sd3_1 hold830 (.A(_01769_),
    .X(net3427));
 sg13g2_dlygate4sd3_1 hold831 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][21] ),
    .X(net3428));
 sg13g2_dlygate4sd3_1 hold832 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][12] ),
    .X(net3429));
 sg13g2_dlygate4sd3_1 hold833 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][18] ),
    .X(net3430));
 sg13g2_dlygate4sd3_1 hold834 (.A(\soc_I.rx_uart_i.fifo_i.ram[13][3] ),
    .X(net3431));
 sg13g2_dlygate4sd3_1 hold835 (.A(_00665_),
    .X(net3432));
 sg13g2_dlygate4sd3_1 hold836 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][8] ),
    .X(net3433));
 sg13g2_dlygate4sd3_1 hold837 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][2] ),
    .X(net3434));
 sg13g2_dlygate4sd3_1 hold838 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][14] ),
    .X(net3435));
 sg13g2_dlygate4sd3_1 hold839 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][15] ),
    .X(net3436));
 sg13g2_dlygate4sd3_1 hold840 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][9] ),
    .X(net3437));
 sg13g2_dlygate4sd3_1 hold841 (.A(\soc_I.rx_uart_i.fifo_i.ram[13][5] ),
    .X(net3438));
 sg13g2_dlygate4sd3_1 hold842 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][3] ),
    .X(net3439));
 sg13g2_dlygate4sd3_1 hold843 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][16] ),
    .X(net3440));
 sg13g2_dlygate4sd3_1 hold844 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][19] ),
    .X(net3441));
 sg13g2_dlygate4sd3_1 hold845 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][15] ),
    .X(net3442));
 sg13g2_dlygate4sd3_1 hold846 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][14] ),
    .X(net3443));
 sg13g2_dlygate4sd3_1 hold847 (.A(\soc_I.qqspi_I.rdata[3] ),
    .X(net3444));
 sg13g2_dlygate4sd3_1 hold848 (.A(_01799_),
    .X(net3445));
 sg13g2_dlygate4sd3_1 hold849 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][30] ),
    .X(net3446));
 sg13g2_dlygate4sd3_1 hold850 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][27] ),
    .X(net3447));
 sg13g2_dlygate4sd3_1 hold851 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][21] ),
    .X(net3448));
 sg13g2_dlygate4sd3_1 hold852 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][29] ),
    .X(net3449));
 sg13g2_dlygate4sd3_1 hold853 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][27] ),
    .X(net3450));
 sg13g2_dlygate4sd3_1 hold854 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][29] ),
    .X(net3451));
 sg13g2_dlygate4sd3_1 hold855 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][28] ),
    .X(net3452));
 sg13g2_dlygate4sd3_1 hold856 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][8] ),
    .X(net3453));
 sg13g2_dlygate4sd3_1 hold857 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][4] ),
    .X(net3454));
 sg13g2_dlygate4sd3_1 hold858 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][13] ),
    .X(net3455));
 sg13g2_dlygate4sd3_1 hold859 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][14] ),
    .X(net3456));
 sg13g2_dlygate4sd3_1 hold860 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][4] ),
    .X(net3457));
 sg13g2_dlygate4sd3_1 hold861 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][12] ),
    .X(net3458));
 sg13g2_dlygate4sd3_1 hold862 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[2] ),
    .X(net3459));
 sg13g2_dlygate4sd3_1 hold863 (.A(_05522_),
    .X(net3460));
 sg13g2_dlygate4sd3_1 hold864 (.A(_01267_),
    .X(net3461));
 sg13g2_dlygate4sd3_1 hold865 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][11] ),
    .X(net3462));
 sg13g2_dlygate4sd3_1 hold866 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][25] ),
    .X(net3463));
 sg13g2_dlygate4sd3_1 hold867 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][8] ),
    .X(net3464));
 sg13g2_dlygate4sd3_1 hold868 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][19] ),
    .X(net3465));
 sg13g2_dlygate4sd3_1 hold869 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][30] ),
    .X(net3466));
 sg13g2_dlygate4sd3_1 hold870 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][31] ),
    .X(net3467));
 sg13g2_dlygate4sd3_1 hold871 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][13] ),
    .X(net3468));
 sg13g2_dlygate4sd3_1 hold872 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[6][15] ),
    .X(net3469));
 sg13g2_dlygate4sd3_1 hold873 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][3] ),
    .X(net3470));
 sg13g2_dlygate4sd3_1 hold874 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[60] ),
    .X(net3471));
 sg13g2_dlygate4sd3_1 hold875 (.A(_05621_),
    .X(net3472));
 sg13g2_dlygate4sd3_1 hold876 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][0] ),
    .X(net3473));
 sg13g2_dlygate4sd3_1 hold877 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][29] ),
    .X(net3474));
 sg13g2_dlygate4sd3_1 hold878 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][29] ),
    .X(net3475));
 sg13g2_dlygate4sd3_1 hold879 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][2] ),
    .X(net3476));
 sg13g2_dlygate4sd3_1 hold880 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][15] ),
    .X(net3477));
 sg13g2_dlygate4sd3_1 hold881 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][13] ),
    .X(net3478));
 sg13g2_dlygate4sd3_1 hold882 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][10] ),
    .X(net3479));
 sg13g2_dlygate4sd3_1 hold883 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][29] ),
    .X(net3480));
 sg13g2_dlygate4sd3_1 hold884 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][27] ),
    .X(net3481));
 sg13g2_dlygate4sd3_1 hold885 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][27] ),
    .X(net3482));
 sg13g2_dlygate4sd3_1 hold886 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][25] ),
    .X(net3483));
 sg13g2_dlygate4sd3_1 hold887 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[52] ),
    .X(net3484));
 sg13g2_dlygate4sd3_1 hold888 (.A(_05608_),
    .X(net3485));
 sg13g2_dlygate4sd3_1 hold889 (.A(_01317_),
    .X(net3486));
 sg13g2_dlygate4sd3_1 hold890 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][31] ),
    .X(net3487));
 sg13g2_dlygate4sd3_1 hold891 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][25] ),
    .X(net3488));
 sg13g2_dlygate4sd3_1 hold892 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][23] ),
    .X(net3489));
 sg13g2_dlygate4sd3_1 hold893 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][7] ),
    .X(net3490));
 sg13g2_dlygate4sd3_1 hold894 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][8] ),
    .X(net3491));
 sg13g2_dlygate4sd3_1 hold895 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][11] ),
    .X(net3492));
 sg13g2_dlygate4sd3_1 hold896 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][23] ),
    .X(net3493));
 sg13g2_dlygate4sd3_1 hold897 (.A(\soc_I.qqspi_I.rdata[17] ),
    .X(net3494));
 sg13g2_dlygate4sd3_1 hold898 (.A(_01813_),
    .X(net3495));
 sg13g2_dlygate4sd3_1 hold899 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][16] ),
    .X(net3496));
 sg13g2_dlygate4sd3_1 hold900 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][14] ),
    .X(net3497));
 sg13g2_dlygate4sd3_1 hold901 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][6] ),
    .X(net3498));
 sg13g2_dlygate4sd3_1 hold902 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][29] ),
    .X(net3499));
 sg13g2_dlygate4sd3_1 hold903 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][1] ),
    .X(net3500));
 sg13g2_dlygate4sd3_1 hold904 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][9] ),
    .X(net3501));
 sg13g2_dlygate4sd3_1 hold905 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][22] ),
    .X(net3502));
 sg13g2_dlygate4sd3_1 hold906 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][11] ),
    .X(net3503));
 sg13g2_dlygate4sd3_1 hold907 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][8] ),
    .X(net3504));
 sg13g2_dlygate4sd3_1 hold908 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][27] ),
    .X(net3505));
 sg13g2_dlygate4sd3_1 hold909 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][24] ),
    .X(net3506));
 sg13g2_dlygate4sd3_1 hold910 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][15] ),
    .X(net3507));
 sg13g2_dlygate4sd3_1 hold911 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][24] ),
    .X(net3508));
 sg13g2_dlygate4sd3_1 hold912 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][1] ),
    .X(net3509));
 sg13g2_dlygate4sd3_1 hold913 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][3] ),
    .X(net3510));
 sg13g2_dlygate4sd3_1 hold914 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][27] ),
    .X(net3511));
 sg13g2_dlygate4sd3_1 hold915 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][11] ),
    .X(net3512));
 sg13g2_dlygate4sd3_1 hold916 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][17] ),
    .X(net3513));
 sg13g2_dlygate4sd3_1 hold917 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[9] ),
    .X(net3514));
 sg13g2_dlygate4sd3_1 hold918 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][27] ),
    .X(net3515));
 sg13g2_dlygate4sd3_1 hold919 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][24] ),
    .X(net3516));
 sg13g2_dlygate4sd3_1 hold920 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][17] ),
    .X(net3517));
 sg13g2_dlygate4sd3_1 hold921 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][17] ),
    .X(net3518));
 sg13g2_dlygate4sd3_1 hold922 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][14] ),
    .X(net3519));
 sg13g2_dlygate4sd3_1 hold923 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][16] ),
    .X(net3520));
 sg13g2_dlygate4sd3_1 hold924 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][11] ),
    .X(net3521));
 sg13g2_dlygate4sd3_1 hold925 (.A(\soc_I.tx_uart_i.wait_states[11] ),
    .X(net3522));
 sg13g2_dlygate4sd3_1 hold926 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][3] ),
    .X(net3523));
 sg13g2_dlygate4sd3_1 hold927 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][18] ),
    .X(net3524));
 sg13g2_dlygate4sd3_1 hold928 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][26] ),
    .X(net3525));
 sg13g2_dlygate4sd3_1 hold929 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][27] ),
    .X(net3526));
 sg13g2_dlygate4sd3_1 hold930 (.A(\soc_I.tx_uart_i.wait_states[10] ),
    .X(net3527));
 sg13g2_dlygate4sd3_1 hold931 (.A(_01933_),
    .X(net3528));
 sg13g2_dlygate4sd3_1 hold932 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][28] ),
    .X(net3529));
 sg13g2_dlygate4sd3_1 hold933 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][3] ),
    .X(net3530));
 sg13g2_dlygate4sd3_1 hold934 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][3] ),
    .X(net3531));
 sg13g2_dlygate4sd3_1 hold935 (.A(\soc_I.rx_uart_i.fifo_i.ram[8][7] ),
    .X(net3532));
 sg13g2_dlygate4sd3_1 hold936 (.A(_02107_),
    .X(net3533));
 sg13g2_dlygate4sd3_1 hold937 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][30] ),
    .X(net3534));
 sg13g2_dlygate4sd3_1 hold938 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][5] ),
    .X(net3535));
 sg13g2_dlygate4sd3_1 hold939 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][24] ),
    .X(net3536));
 sg13g2_dlygate4sd3_1 hold940 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][21] ),
    .X(net3537));
 sg13g2_dlygate4sd3_1 hold941 (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[24] ),
    .X(net3538));
 sg13g2_dlygate4sd3_1 hold942 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][12] ),
    .X(net3539));
 sg13g2_dlygate4sd3_1 hold943 (.A(\soc_I.rx_uart_i.fifo_i.ram[10][2] ),
    .X(net3540));
 sg13g2_dlygate4sd3_1 hold944 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][25] ),
    .X(net3541));
 sg13g2_dlygate4sd3_1 hold945 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][10] ),
    .X(net3542));
 sg13g2_dlygate4sd3_1 hold946 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][8] ),
    .X(net3543));
 sg13g2_dlygate4sd3_1 hold947 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][13] ),
    .X(net3544));
 sg13g2_dlygate4sd3_1 hold948 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][15] ),
    .X(net3545));
 sg13g2_dlygate4sd3_1 hold949 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][31] ),
    .X(net3546));
 sg13g2_dlygate4sd3_1 hold950 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][21] ),
    .X(net3547));
 sg13g2_dlygate4sd3_1 hold951 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][31] ),
    .X(net3548));
 sg13g2_dlygate4sd3_1 hold952 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][18] ),
    .X(net3549));
 sg13g2_dlygate4sd3_1 hold953 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][3] ),
    .X(net3550));
 sg13g2_dlygate4sd3_1 hold954 (.A(\soc_I.rx_uart_i.fifo_i.ram[14][7] ),
    .X(net3551));
 sg13g2_dlygate4sd3_1 hold955 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][7] ),
    .X(net3552));
 sg13g2_dlygate4sd3_1 hold956 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][21] ),
    .X(net3553));
 sg13g2_dlygate4sd3_1 hold957 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][4] ),
    .X(net3554));
 sg13g2_dlygate4sd3_1 hold958 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][7] ),
    .X(net3555));
 sg13g2_dlygate4sd3_1 hold959 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][22] ),
    .X(net3556));
 sg13g2_dlygate4sd3_1 hold960 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][24] ),
    .X(net3557));
 sg13g2_dlygate4sd3_1 hold961 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[0] ),
    .X(net3558));
 sg13g2_dlygate4sd3_1 hold962 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][20] ),
    .X(net3559));
 sg13g2_dlygate4sd3_1 hold963 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][25] ),
    .X(net3560));
 sg13g2_dlygate4sd3_1 hold964 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][18] ),
    .X(net3561));
 sg13g2_dlygate4sd3_1 hold965 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][4] ),
    .X(net3562));
 sg13g2_dlygate4sd3_1 hold966 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][0] ),
    .X(net3563));
 sg13g2_dlygate4sd3_1 hold967 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][11] ),
    .X(net3564));
 sg13g2_dlygate4sd3_1 hold968 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][0] ),
    .X(net3565));
 sg13g2_dlygate4sd3_1 hold969 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][18] ),
    .X(net3566));
 sg13g2_dlygate4sd3_1 hold970 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][2] ),
    .X(net3567));
 sg13g2_dlygate4sd3_1 hold971 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][26] ),
    .X(net3568));
 sg13g2_dlygate4sd3_1 hold972 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][20] ),
    .X(net3569));
 sg13g2_dlygate4sd3_1 hold973 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][23] ),
    .X(net3570));
 sg13g2_dlygate4sd3_1 hold974 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][19] ),
    .X(net3571));
 sg13g2_dlygate4sd3_1 hold975 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][26] ),
    .X(net3572));
 sg13g2_dlygate4sd3_1 hold976 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][6] ),
    .X(net3573));
 sg13g2_dlygate4sd3_1 hold977 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][28] ),
    .X(net3574));
 sg13g2_dlygate4sd3_1 hold978 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][25] ),
    .X(net3575));
 sg13g2_dlygate4sd3_1 hold979 (.A(\soc_I.rx_uart_i.fifo_i.rd_ptr[2] ),
    .X(net3576));
 sg13g2_dlygate4sd3_1 hold980 (.A(_06958_),
    .X(net3577));
 sg13g2_dlygate4sd3_1 hold981 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][18] ),
    .X(net3578));
 sg13g2_dlygate4sd3_1 hold982 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][17] ),
    .X(net3579));
 sg13g2_dlygate4sd3_1 hold983 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][28] ),
    .X(net3580));
 sg13g2_dlygate4sd3_1 hold984 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][14] ),
    .X(net3581));
 sg13g2_dlygate4sd3_1 hold985 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][24] ),
    .X(net3582));
 sg13g2_dlygate4sd3_1 hold986 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][16] ),
    .X(net3583));
 sg13g2_dlygate4sd3_1 hold987 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][7] ),
    .X(net3584));
 sg13g2_dlygate4sd3_1 hold988 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[15] ),
    .X(net3585));
 sg13g2_dlygate4sd3_1 hold989 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][27] ),
    .X(net3586));
 sg13g2_dlygate4sd3_1 hold990 (.A(sio1_so_miso_o),
    .X(net3587));
 sg13g2_dlygate4sd3_1 hold991 (.A(_07298_),
    .X(net3588));
 sg13g2_dlygate4sd3_1 hold992 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][16] ),
    .X(net3589));
 sg13g2_dlygate4sd3_1 hold993 (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[10] ),
    .X(net3590));
 sg13g2_dlygate4sd3_1 hold994 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][26] ),
    .X(net3591));
 sg13g2_dlygate4sd3_1 hold995 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][21] ),
    .X(net3592));
 sg13g2_dlygate4sd3_1 hold996 (.A(\soc_I.clint_I.mtime[5] ),
    .X(net3593));
 sg13g2_dlygate4sd3_1 hold997 (.A(_01637_),
    .X(net3594));
 sg13g2_dlygate4sd3_1 hold998 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][3] ),
    .X(net3595));
 sg13g2_dlygate4sd3_1 hold999 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][23] ),
    .X(net3596));
 sg13g2_dlygate4sd3_1 hold1000 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][26] ),
    .X(net3597));
 sg13g2_dlygate4sd3_1 hold1001 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][31] ),
    .X(net3598));
 sg13g2_dlygate4sd3_1 hold1002 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][6] ),
    .X(net3599));
 sg13g2_dlygate4sd3_1 hold1003 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][31] ),
    .X(net3600));
 sg13g2_dlygate4sd3_1 hold1004 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][16] ),
    .X(net3601));
 sg13g2_dlygate4sd3_1 hold1005 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][19] ),
    .X(net3602));
 sg13g2_dlygate4sd3_1 hold1006 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][12] ),
    .X(net3603));
 sg13g2_dlygate4sd3_1 hold1007 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[13] ),
    .X(net3604));
 sg13g2_dlygate4sd3_1 hold1008 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][11] ),
    .X(net3605));
 sg13g2_dlygate4sd3_1 hold1009 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][11] ),
    .X(net3606));
 sg13g2_dlygate4sd3_1 hold1010 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[10] ),
    .X(net3607));
 sg13g2_dlygate4sd3_1 hold1011 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][12] ),
    .X(net3608));
 sg13g2_dlygate4sd3_1 hold1012 (.A(\soc_I.rx_uart_i.fifo_i.ram[10][5] ),
    .X(net3609));
 sg13g2_dlygate4sd3_1 hold1013 (.A(_00643_),
    .X(net3610));
 sg13g2_dlygate4sd3_1 hold1014 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][16] ),
    .X(net3611));
 sg13g2_dlygate4sd3_1 hold1015 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][3] ),
    .X(net3612));
 sg13g2_dlygate4sd3_1 hold1016 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][2] ),
    .X(net3613));
 sg13g2_dlygate4sd3_1 hold1017 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][2] ),
    .X(net3614));
 sg13g2_dlygate4sd3_1 hold1018 (.A(\soc_I.tx_uart_i.wait_states[5] ),
    .X(net3615));
 sg13g2_dlygate4sd3_1 hold1019 (.A(_01928_),
    .X(net3616));
 sg13g2_dlygate4sd3_1 hold1020 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][12] ),
    .X(net3617));
 sg13g2_dlygate4sd3_1 hold1021 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][30] ),
    .X(net3618));
 sg13g2_dlygate4sd3_1 hold1022 (.A(\soc_I.rx_uart_i.fifo_i.ram[14][1] ),
    .X(net3619));
 sg13g2_dlygate4sd3_1 hold1023 (.A(\soc_I.rx_uart_i.fifo_i.ram[8][6] ),
    .X(net3620));
 sg13g2_dlygate4sd3_1 hold1024 (.A(_02106_),
    .X(net3621));
 sg13g2_dlygate4sd3_1 hold1025 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[1] ),
    .X(net3622));
 sg13g2_dlygate4sd3_1 hold1026 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][23] ),
    .X(net3623));
 sg13g2_dlygate4sd3_1 hold1027 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][10] ),
    .X(net3624));
 sg13g2_dlygate4sd3_1 hold1028 (.A(\soc_I.clint_I.tick_cnt[2] ),
    .X(net3625));
 sg13g2_dlygate4sd3_1 hold1029 (.A(_06225_),
    .X(net3626));
 sg13g2_dlygate4sd3_1 hold1030 (.A(_01603_),
    .X(net3627));
 sg13g2_dlygate4sd3_1 hold1031 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][7] ),
    .X(net3628));
 sg13g2_dlygate4sd3_1 hold1032 (.A(\soc_I.qqspi_I.rdata[20] ),
    .X(net3629));
 sg13g2_dlygate4sd3_1 hold1033 (.A(_01816_),
    .X(net3630));
 sg13g2_dlygate4sd3_1 hold1034 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][8] ),
    .X(net3631));
 sg13g2_dlygate4sd3_1 hold1035 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][21] ),
    .X(net3632));
 sg13g2_dlygate4sd3_1 hold1036 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][4] ),
    .X(net3633));
 sg13g2_dlygate4sd3_1 hold1037 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][1] ),
    .X(net3634));
 sg13g2_dlygate4sd3_1 hold1038 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][15] ),
    .X(net3635));
 sg13g2_dlygate4sd3_1 hold1039 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][17] ),
    .X(net3636));
 sg13g2_dlygate4sd3_1 hold1040 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][7] ),
    .X(net3637));
 sg13g2_dlygate4sd3_1 hold1041 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][12] ),
    .X(net3638));
 sg13g2_dlygate4sd3_1 hold1042 (.A(\soc_I.rx_uart_i.fifo_i.ram[10][1] ),
    .X(net3639));
 sg13g2_dlygate4sd3_1 hold1043 (.A(_00639_),
    .X(net3640));
 sg13g2_dlygate4sd3_1 hold1044 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][8] ),
    .X(net3641));
 sg13g2_dlygate4sd3_1 hold1045 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][25] ),
    .X(net3642));
 sg13g2_dlygate4sd3_1 hold1046 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[20] ),
    .X(net3643));
 sg13g2_dlygate4sd3_1 hold1047 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][7] ),
    .X(net3644));
 sg13g2_dlygate4sd3_1 hold1048 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][20] ),
    .X(net3645));
 sg13g2_dlygate4sd3_1 hold1049 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[21] ),
    .X(net3646));
 sg13g2_dlygate4sd3_1 hold1050 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][26] ),
    .X(net3647));
 sg13g2_dlygate4sd3_1 hold1051 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][17] ),
    .X(net3648));
 sg13g2_dlygate4sd3_1 hold1052 (.A(_02232_),
    .X(net3649));
 sg13g2_dlygate4sd3_1 hold1053 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][11] ),
    .X(net3650));
 sg13g2_dlygate4sd3_1 hold1054 (.A(\soc_I.qqspi_I.rdata[12] ),
    .X(net3651));
 sg13g2_dlygate4sd3_1 hold1055 (.A(_01808_),
    .X(net3652));
 sg13g2_dlygate4sd3_1 hold1056 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][29] ),
    .X(net3653));
 sg13g2_dlygate4sd3_1 hold1057 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][1] ),
    .X(net3654));
 sg13g2_dlygate4sd3_1 hold1058 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][22] ),
    .X(net3655));
 sg13g2_dlygate4sd3_1 hold1059 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][28] ),
    .X(net3656));
 sg13g2_dlygate4sd3_1 hold1060 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][27] ),
    .X(net3657));
 sg13g2_dlygate4sd3_1 hold1061 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][12] ),
    .X(net3658));
 sg13g2_dlygate4sd3_1 hold1062 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][18] ),
    .X(net3659));
 sg13g2_dlygate4sd3_1 hold1063 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][28] ),
    .X(net3660));
 sg13g2_dlygate4sd3_1 hold1064 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][15] ),
    .X(net3661));
 sg13g2_dlygate4sd3_1 hold1065 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][31] ),
    .X(net3662));
 sg13g2_dlygate4sd3_1 hold1066 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][30] ),
    .X(net3663));
 sg13g2_dlygate4sd3_1 hold1067 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][4] ),
    .X(net3664));
 sg13g2_dlygate4sd3_1 hold1068 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][22] ),
    .X(net3665));
 sg13g2_dlygate4sd3_1 hold1069 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][17] ),
    .X(net3666));
 sg13g2_dlygate4sd3_1 hold1070 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][2] ),
    .X(net3667));
 sg13g2_dlygate4sd3_1 hold1071 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][23] ),
    .X(net3668));
 sg13g2_dlygate4sd3_1 hold1072 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][11] ),
    .X(net3669));
 sg13g2_dlygate4sd3_1 hold1073 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[63] ),
    .X(net3670));
 sg13g2_dlygate4sd3_1 hold1074 (.A(_01328_),
    .X(net3671));
 sg13g2_dlygate4sd3_1 hold1075 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][1] ),
    .X(net3672));
 sg13g2_dlygate4sd3_1 hold1076 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[25] ),
    .X(net3673));
 sg13g2_dlygate4sd3_1 hold1077 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[15] ),
    .X(net3674));
 sg13g2_dlygate4sd3_1 hold1078 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][7] ),
    .X(net3675));
 sg13g2_dlygate4sd3_1 hold1079 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][15] ),
    .X(net3676));
 sg13g2_dlygate4sd3_1 hold1080 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][29] ),
    .X(net3677));
 sg13g2_dlygate4sd3_1 hold1081 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][26] ),
    .X(net3678));
 sg13g2_dlygate4sd3_1 hold1082 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][23] ),
    .X(net3679));
 sg13g2_dlygate4sd3_1 hold1083 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][19] ),
    .X(net3680));
 sg13g2_dlygate4sd3_1 hold1084 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][21] ),
    .X(net3681));
 sg13g2_dlygate4sd3_1 hold1085 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][4] ),
    .X(net3682));
 sg13g2_dlygate4sd3_1 hold1086 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][0] ),
    .X(net3683));
 sg13g2_dlygate4sd3_1 hold1087 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][23] ),
    .X(net3684));
 sg13g2_dlygate4sd3_1 hold1088 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][28] ),
    .X(net3685));
 sg13g2_dlygate4sd3_1 hold1089 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][31] ),
    .X(net3686));
 sg13g2_dlygate4sd3_1 hold1090 (.A(\soc_I.tx_uart_i.wait_states[12] ),
    .X(net3687));
 sg13g2_dlygate4sd3_1 hold1091 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[34] ),
    .X(net3688));
 sg13g2_dlygate4sd3_1 hold1092 (.A(_05578_),
    .X(net3689));
 sg13g2_dlygate4sd3_1 hold1093 (.A(_01299_),
    .X(net3690));
 sg13g2_dlygate4sd3_1 hold1094 (.A(\soc_I.rx_uart_i.fifo_i.ram[8][3] ),
    .X(net3691));
 sg13g2_dlygate4sd3_1 hold1095 (.A(_02103_),
    .X(net3692));
 sg13g2_dlygate4sd3_1 hold1096 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][28] ),
    .X(net3693));
 sg13g2_dlygate4sd3_1 hold1097 (.A(\soc_I.clint_I.mtime[3] ),
    .X(net3694));
 sg13g2_dlygate4sd3_1 hold1098 (.A(_01635_),
    .X(net3695));
 sg13g2_dlygate4sd3_1 hold1099 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][29] ),
    .X(net3696));
 sg13g2_dlygate4sd3_1 hold1100 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][22] ),
    .X(net3697));
 sg13g2_dlygate4sd3_1 hold1101 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][10] ),
    .X(net3698));
 sg13g2_dlygate4sd3_1 hold1102 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][20] ),
    .X(net3699));
 sg13g2_dlygate4sd3_1 hold1103 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][6] ),
    .X(net3700));
 sg13g2_dlygate4sd3_1 hold1104 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[26] ),
    .X(net3701));
 sg13g2_dlygate4sd3_1 hold1105 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][22] ),
    .X(net3702));
 sg13g2_dlygate4sd3_1 hold1106 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][5] ),
    .X(net3703));
 sg13g2_dlygate4sd3_1 hold1107 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][12] ),
    .X(net3704));
 sg13g2_dlygate4sd3_1 hold1108 (.A(\soc_I.spi0_I.spi_buf[7] ),
    .X(net3705));
 sg13g2_dlygate4sd3_1 hold1109 (.A(_01978_),
    .X(net3706));
 sg13g2_dlygate4sd3_1 hold1110 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][12] ),
    .X(net3707));
 sg13g2_dlygate4sd3_1 hold1111 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][0] ),
    .X(net3708));
 sg13g2_dlygate4sd3_1 hold1112 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][23] ),
    .X(net3709));
 sg13g2_dlygate4sd3_1 hold1113 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[42] ),
    .X(net3710));
 sg13g2_dlygate4sd3_1 hold1114 (.A(_05591_),
    .X(net3711));
 sg13g2_dlygate4sd3_1 hold1115 (.A(_01307_),
    .X(net3712));
 sg13g2_dlygate4sd3_1 hold1116 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][25] ),
    .X(net3713));
 sg13g2_dlygate4sd3_1 hold1117 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][14] ),
    .X(net3714));
 sg13g2_dlygate4sd3_1 hold1118 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][29] ),
    .X(net3715));
 sg13g2_dlygate4sd3_1 hold1119 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][3] ),
    .X(net3716));
 sg13g2_dlygate4sd3_1 hold1120 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][19] ),
    .X(net3717));
 sg13g2_dlygate4sd3_1 hold1121 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][12] ),
    .X(net3718));
 sg13g2_dlygate4sd3_1 hold1122 (.A(\soc_I.spi0_I.spi_buf[1] ),
    .X(net3719));
 sg13g2_dlygate4sd3_1 hold1123 (.A(_01972_),
    .X(net3720));
 sg13g2_dlygate4sd3_1 hold1124 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][14] ),
    .X(net3721));
 sg13g2_dlygate4sd3_1 hold1125 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][30] ),
    .X(net3722));
 sg13g2_dlygate4sd3_1 hold1126 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][21] ),
    .X(net3723));
 sg13g2_dlygate4sd3_1 hold1127 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][17] ),
    .X(net3724));
 sg13g2_dlygate4sd3_1 hold1128 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][2] ),
    .X(net3725));
 sg13g2_dlygate4sd3_1 hold1129 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][27] ),
    .X(net3726));
 sg13g2_dlygate4sd3_1 hold1130 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][27] ),
    .X(net3727));
 sg13g2_dlygate4sd3_1 hold1131 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][20] ),
    .X(net3728));
 sg13g2_dlygate4sd3_1 hold1132 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][1] ),
    .X(net3729));
 sg13g2_dlygate4sd3_1 hold1133 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][14] ),
    .X(net3730));
 sg13g2_dlygate4sd3_1 hold1134 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][2] ),
    .X(net3731));
 sg13g2_dlygate4sd3_1 hold1135 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][8] ),
    .X(net3732));
 sg13g2_dlygate4sd3_1 hold1136 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][13] ),
    .X(net3733));
 sg13g2_dlygate4sd3_1 hold1137 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][23] ),
    .X(net3734));
 sg13g2_dlygate4sd3_1 hold1138 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][24] ),
    .X(net3735));
 sg13g2_dlygate4sd3_1 hold1139 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][18] ),
    .X(net3736));
 sg13g2_dlygate4sd3_1 hold1140 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[40] ),
    .X(net3737));
 sg13g2_dlygate4sd3_1 hold1141 (.A(_05588_),
    .X(net3738));
 sg13g2_dlygate4sd3_1 hold1142 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][23] ),
    .X(net3739));
 sg13g2_dlygate4sd3_1 hold1143 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][22] ),
    .X(net3740));
 sg13g2_dlygate4sd3_1 hold1144 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][14] ),
    .X(net3741));
 sg13g2_dlygate4sd3_1 hold1145 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][20] ),
    .X(net3742));
 sg13g2_dlygate4sd3_1 hold1146 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[22][25] ),
    .X(net3743));
 sg13g2_dlygate4sd3_1 hold1147 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][4] ),
    .X(net3744));
 sg13g2_dlygate4sd3_1 hold1148 (.A(\soc_I.qqspi_I.rdata[8] ),
    .X(net3745));
 sg13g2_dlygate4sd3_1 hold1149 (.A(_01804_),
    .X(net3746));
 sg13g2_dlygate4sd3_1 hold1150 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[18][26] ),
    .X(net3747));
 sg13g2_dlygate4sd3_1 hold1151 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][1] ),
    .X(net3748));
 sg13g2_dlygate4sd3_1 hold1152 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][2] ),
    .X(net3749));
 sg13g2_dlygate4sd3_1 hold1153 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][4] ),
    .X(net3750));
 sg13g2_dlygate4sd3_1 hold1154 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][19] ),
    .X(net3751));
 sg13g2_dlygate4sd3_1 hold1155 (.A(\soc_I.rx_uart_i.fifo_i.ram[10][4] ),
    .X(net3752));
 sg13g2_dlygate4sd3_1 hold1156 (.A(_00642_),
    .X(net3753));
 sg13g2_dlygate4sd3_1 hold1157 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][23] ),
    .X(net3754));
 sg13g2_dlygate4sd3_1 hold1158 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][8] ),
    .X(net3755));
 sg13g2_dlygate4sd3_1 hold1159 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][5] ),
    .X(net3756));
 sg13g2_dlygate4sd3_1 hold1160 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.bit_idx[0] ),
    .X(net3757));
 sg13g2_dlygate4sd3_1 hold1161 (.A(_05628_),
    .X(net3758));
 sg13g2_dlygate4sd3_1 hold1162 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][23] ),
    .X(net3759));
 sg13g2_dlygate4sd3_1 hold1163 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[24] ),
    .X(net3760));
 sg13g2_dlygate4sd3_1 hold1164 (.A(_05561_),
    .X(net3761));
 sg13g2_dlygate4sd3_1 hold1165 (.A(_01289_),
    .X(net3762));
 sg13g2_dlygate4sd3_1 hold1166 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][17] ),
    .X(net3763));
 sg13g2_dlygate4sd3_1 hold1167 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][16] ),
    .X(net3764));
 sg13g2_dlygate4sd3_1 hold1168 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][7] ),
    .X(net3765));
 sg13g2_dlygate4sd3_1 hold1169 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][18] ),
    .X(net3766));
 sg13g2_dlygate4sd3_1 hold1170 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][5] ),
    .X(net3767));
 sg13g2_dlygate4sd3_1 hold1171 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][2] ),
    .X(net3768));
 sg13g2_dlygate4sd3_1 hold1172 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][23] ),
    .X(net3769));
 sg13g2_dlygate4sd3_1 hold1173 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][22] ),
    .X(net3770));
 sg13g2_dlygate4sd3_1 hold1174 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][13] ),
    .X(net3771));
 sg13g2_dlygate4sd3_1 hold1175 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[5] ),
    .X(net3772));
 sg13g2_dlygate4sd3_1 hold1176 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][21] ),
    .X(net3773));
 sg13g2_dlygate4sd3_1 hold1177 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[48] ),
    .X(net3774));
 sg13g2_dlygate4sd3_1 hold1178 (.A(_05601_),
    .X(net3775));
 sg13g2_dlygate4sd3_1 hold1179 (.A(_01313_),
    .X(net3776));
 sg13g2_dlygate4sd3_1 hold1180 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][17] ),
    .X(net3777));
 sg13g2_dlygate4sd3_1 hold1181 (.A(_02352_),
    .X(net3778));
 sg13g2_dlygate4sd3_1 hold1182 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][25] ),
    .X(net3779));
 sg13g2_dlygate4sd3_1 hold1183 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[22] ),
    .X(net3780));
 sg13g2_dlygate4sd3_1 hold1184 (.A(_05558_),
    .X(net3781));
 sg13g2_dlygate4sd3_1 hold1185 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][24] ),
    .X(net3782));
 sg13g2_dlygate4sd3_1 hold1186 (.A(\soc_I.clint_I.mtime[1] ),
    .X(net3783));
 sg13g2_dlygate4sd3_1 hold1187 (.A(_06283_),
    .X(net3784));
 sg13g2_dlygate4sd3_1 hold1188 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][24] ),
    .X(net3785));
 sg13g2_dlygate4sd3_1 hold1189 (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[28] ),
    .X(net3786));
 sg13g2_dlygate4sd3_1 hold1190 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][16] ),
    .X(net3787));
 sg13g2_dlygate4sd3_1 hold1191 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][19] ),
    .X(net3788));
 sg13g2_dlygate4sd3_1 hold1192 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][26] ),
    .X(net3789));
 sg13g2_dlygate4sd3_1 hold1193 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][4] ),
    .X(net3790));
 sg13g2_dlygate4sd3_1 hold1194 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[48] ),
    .X(net3791));
 sg13g2_dlygate4sd3_1 hold1195 (.A(_01185_),
    .X(net3792));
 sg13g2_dlygate4sd3_1 hold1196 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][26] ),
    .X(net3793));
 sg13g2_dlygate4sd3_1 hold1197 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][24] ),
    .X(net3794));
 sg13g2_dlygate4sd3_1 hold1198 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[12] ),
    .X(net3795));
 sg13g2_dlygate4sd3_1 hold1199 (.A(_05541_),
    .X(net3796));
 sg13g2_dlygate4sd3_1 hold1200 (.A(_01277_),
    .X(net3797));
 sg13g2_dlygate4sd3_1 hold1201 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][4] ),
    .X(net3798));
 sg13g2_dlygate4sd3_1 hold1202 (.A(\soc_I.clint_I.mtime[6] ),
    .X(net3799));
 sg13g2_dlygate4sd3_1 hold1203 (.A(_06298_),
    .X(net3800));
 sg13g2_dlygate4sd3_1 hold1204 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][4] ),
    .X(net3801));
 sg13g2_dlygate4sd3_1 hold1205 (.A(\gpio_uo_out[5] ),
    .X(net3802));
 sg13g2_dlygate4sd3_1 hold1206 (.A(_01792_),
    .X(net3803));
 sg13g2_dlygate4sd3_1 hold1207 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][9] ),
    .X(net3804));
 sg13g2_dlygate4sd3_1 hold1208 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][24] ),
    .X(net3805));
 sg13g2_dlygate4sd3_1 hold1209 (.A(\soc_I.rx_uart_i.fifo_i.ram[8][5] ),
    .X(net3806));
 sg13g2_dlygate4sd3_1 hold1210 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][12] ),
    .X(net3807));
 sg13g2_dlygate4sd3_1 hold1211 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][6] ),
    .X(net3808));
 sg13g2_dlygate4sd3_1 hold1212 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][30] ),
    .X(net3809));
 sg13g2_dlygate4sd3_1 hold1213 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][14] ),
    .X(net3810));
 sg13g2_dlygate4sd3_1 hold1214 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][31] ),
    .X(net3811));
 sg13g2_dlygate4sd3_1 hold1215 (.A(\soc_I.rx_uart_i.fifo_i.ram[12][5] ),
    .X(net3812));
 sg13g2_dlygate4sd3_1 hold1216 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][3] ),
    .X(net3813));
 sg13g2_dlygate4sd3_1 hold1217 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][19] ),
    .X(net3814));
 sg13g2_dlygate4sd3_1 hold1218 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][27] ),
    .X(net3815));
 sg13g2_dlygate4sd3_1 hold1219 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][27] ),
    .X(net3816));
 sg13g2_dlygate4sd3_1 hold1220 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[6] ),
    .X(net3817));
 sg13g2_dlygate4sd3_1 hold1221 (.A(_05530_),
    .X(net3818));
 sg13g2_dlygate4sd3_1 hold1222 (.A(\soc_I.spi0_I.tick_cnt[2] ),
    .X(net3819));
 sg13g2_dlygate4sd3_1 hold1223 (.A(_06614_),
    .X(net3820));
 sg13g2_dlygate4sd3_1 hold1224 (.A(_01765_),
    .X(net3821));
 sg13g2_dlygate4sd3_1 hold1225 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][14] ),
    .X(net3822));
 sg13g2_dlygate4sd3_1 hold1226 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][13] ),
    .X(net3823));
 sg13g2_dlygate4sd3_1 hold1227 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][25] ),
    .X(net3824));
 sg13g2_dlygate4sd3_1 hold1228 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][15] ),
    .X(net3825));
 sg13g2_dlygate4sd3_1 hold1229 (.A(_01728_),
    .X(net3826));
 sg13g2_dlygate4sd3_1 hold1230 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][1] ),
    .X(net3827));
 sg13g2_dlygate4sd3_1 hold1231 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][28] ),
    .X(net3828));
 sg13g2_dlygate4sd3_1 hold1232 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][4] ),
    .X(net3829));
 sg13g2_dlygate4sd3_1 hold1233 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][25] ),
    .X(net3830));
 sg13g2_dlygate4sd3_1 hold1234 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][29] ),
    .X(net3831));
 sg13g2_dlygate4sd3_1 hold1235 (.A(\soc_I.rx_uart_i.fifo_i.ram[12][2] ),
    .X(net3832));
 sg13g2_dlygate4sd3_1 hold1236 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][3] ),
    .X(net3833));
 sg13g2_dlygate4sd3_1 hold1237 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][17] ),
    .X(net3834));
 sg13g2_dlygate4sd3_1 hold1238 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][0] ),
    .X(net3835));
 sg13g2_dlygate4sd3_1 hold1239 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][31] ),
    .X(net3836));
 sg13g2_dlygate4sd3_1 hold1240 (.A(\soc_I.rx_uart_i.fifo_i.cnt[3] ),
    .X(net3837));
 sg13g2_dlygate4sd3_1 hold1241 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][27] ),
    .X(net3838));
 sg13g2_dlygate4sd3_1 hold1242 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][12] ),
    .X(net3839));
 sg13g2_dlygate4sd3_1 hold1243 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][18] ),
    .X(net3840));
 sg13g2_dlygate4sd3_1 hold1244 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][12] ),
    .X(net3841));
 sg13g2_dlygate4sd3_1 hold1245 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][20] ),
    .X(net3842));
 sg13g2_dlygate4sd3_1 hold1246 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][31] ),
    .X(net3843));
 sg13g2_dlygate4sd3_1 hold1247 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][5] ),
    .X(net3844));
 sg13g2_dlygate4sd3_1 hold1248 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][21] ),
    .X(net3845));
 sg13g2_dlygate4sd3_1 hold1249 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][24] ),
    .X(net3846));
 sg13g2_dlygate4sd3_1 hold1250 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][0] ),
    .X(net3847));
 sg13g2_dlygate4sd3_1 hold1251 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][12] ),
    .X(net3848));
 sg13g2_dlygate4sd3_1 hold1252 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][27] ),
    .X(net3849));
 sg13g2_dlygate4sd3_1 hold1253 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][10] ),
    .X(net3850));
 sg13g2_dlygate4sd3_1 hold1254 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][20] ),
    .X(net3851));
 sg13g2_dlygate4sd3_1 hold1255 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[12] ),
    .X(net3852));
 sg13g2_dlygate4sd3_1 hold1256 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][27] ),
    .X(net3853));
 sg13g2_dlygate4sd3_1 hold1257 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[24] ),
    .X(net3854));
 sg13g2_dlygate4sd3_1 hold1258 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][16] ),
    .X(net3855));
 sg13g2_dlygate4sd3_1 hold1259 (.A(\soc_I.spi0_I.state ),
    .X(net3856));
 sg13g2_dlygate4sd3_1 hold1260 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[27] ),
    .X(net3857));
 sg13g2_dlygate4sd3_1 hold1261 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][11] ),
    .X(net3858));
 sg13g2_dlygate4sd3_1 hold1262 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[30] ),
    .X(net3859));
 sg13g2_dlygate4sd3_1 hold1263 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[53] ),
    .X(net3860));
 sg13g2_dlygate4sd3_1 hold1264 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][30] ),
    .X(net3861));
 sg13g2_dlygate4sd3_1 hold1265 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][18] ),
    .X(net3862));
 sg13g2_dlygate4sd3_1 hold1266 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][21] ),
    .X(net3863));
 sg13g2_dlygate4sd3_1 hold1267 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][23] ),
    .X(net3864));
 sg13g2_dlygate4sd3_1 hold1268 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][23] ),
    .X(net3865));
 sg13g2_dlygate4sd3_1 hold1269 (.A(\soc_I.spi0_I.rx_data[0] ),
    .X(net3866));
 sg13g2_dlygate4sd3_1 hold1270 (.A(_07177_),
    .X(net3867));
 sg13g2_dlygate4sd3_1 hold1271 (.A(_01971_),
    .X(net3868));
 sg13g2_dlygate4sd3_1 hold1272 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[26] ),
    .X(net3869));
 sg13g2_dlygate4sd3_1 hold1273 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][31] ),
    .X(net3870));
 sg13g2_dlygate4sd3_1 hold1274 (.A(\soc_I.spi0_I.tick_cnt[3] ),
    .X(net3871));
 sg13g2_dlygate4sd3_1 hold1275 (.A(_06616_),
    .X(net3872));
 sg13g2_dlygate4sd3_1 hold1276 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][11] ),
    .X(net3873));
 sg13g2_dlygate4sd3_1 hold1277 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][1] ),
    .X(net3874));
 sg13g2_dlygate4sd3_1 hold1278 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][29] ),
    .X(net3875));
 sg13g2_dlygate4sd3_1 hold1279 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[25][26] ),
    .X(net3876));
 sg13g2_dlygate4sd3_1 hold1280 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][8] ),
    .X(net3877));
 sg13g2_dlygate4sd3_1 hold1281 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][21] ),
    .X(net3878));
 sg13g2_dlygate4sd3_1 hold1282 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][29] ),
    .X(net3879));
 sg13g2_dlygate4sd3_1 hold1283 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][11] ),
    .X(net3880));
 sg13g2_dlygate4sd3_1 hold1284 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][14] ),
    .X(net3881));
 sg13g2_dlygate4sd3_1 hold1285 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][3] ),
    .X(net3882));
 sg13g2_dlygate4sd3_1 hold1286 (.A(\soc_I.qqspi_I.rdata[9] ),
    .X(net3883));
 sg13g2_dlygate4sd3_1 hold1287 (.A(_01805_),
    .X(net3884));
 sg13g2_dlygate4sd3_1 hold1288 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[30] ),
    .X(net3885));
 sg13g2_dlygate4sd3_1 hold1289 (.A(_04556_),
    .X(net3886));
 sg13g2_dlygate4sd3_1 hold1290 (.A(_01033_),
    .X(net3887));
 sg13g2_dlygate4sd3_1 hold1291 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][30] ),
    .X(net3888));
 sg13g2_dlygate4sd3_1 hold1292 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][15] ),
    .X(net3889));
 sg13g2_dlygate4sd3_1 hold1293 (.A(_00251_),
    .X(net3890));
 sg13g2_dlygate4sd3_1 hold1294 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[2][19] ),
    .X(net3891));
 sg13g2_dlygate4sd3_1 hold1295 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][18] ),
    .X(net3892));
 sg13g2_dlygate4sd3_1 hold1296 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][5] ),
    .X(net3893));
 sg13g2_dlygate4sd3_1 hold1297 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[16][27] ),
    .X(net3894));
 sg13g2_dlygate4sd3_1 hold1298 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[17][26] ),
    .X(net3895));
 sg13g2_dlygate4sd3_1 hold1299 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][19] ),
    .X(net3896));
 sg13g2_dlygate4sd3_1 hold1300 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][14] ),
    .X(net3897));
 sg13g2_dlygate4sd3_1 hold1301 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][15] ),
    .X(net3898));
 sg13g2_dlygate4sd3_1 hold1302 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][7] ),
    .X(net3899));
 sg13g2_dlygate4sd3_1 hold1303 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][10] ),
    .X(net3900));
 sg13g2_dlygate4sd3_1 hold1304 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][22] ),
    .X(net3901));
 sg13g2_dlygate4sd3_1 hold1305 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][7] ),
    .X(net3902));
 sg13g2_dlygate4sd3_1 hold1306 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][15] ),
    .X(net3903));
 sg13g2_dlygate4sd3_1 hold1307 (.A(_00725_),
    .X(net3904));
 sg13g2_dlygate4sd3_1 hold1308 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[14][4] ),
    .X(net3905));
 sg13g2_dlygate4sd3_1 hold1309 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][21] ),
    .X(net3906));
 sg13g2_dlygate4sd3_1 hold1310 (.A(\soc_I.rx_uart_i.fifo_i.rd_ptr[1] ),
    .X(net3907));
 sg13g2_dlygate4sd3_1 hold1311 (.A(_06954_),
    .X(net3908));
 sg13g2_dlygate4sd3_1 hold1312 (.A(_01864_),
    .X(net3909));
 sg13g2_dlygate4sd3_1 hold1313 (.A(_00302_),
    .X(net3910));
 sg13g2_dlygate4sd3_1 hold1314 (.A(_01632_),
    .X(net3911));
 sg13g2_dlygate4sd3_1 hold1315 (.A(\soc_I.rx_uart_i.fifo_i.ram[11][3] ),
    .X(net3912));
 sg13g2_dlygate4sd3_1 hold1316 (.A(_00649_),
    .X(net3913));
 sg13g2_dlygate4sd3_1 hold1317 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][13] ),
    .X(net3914));
 sg13g2_dlygate4sd3_1 hold1318 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][25] ),
    .X(net3915));
 sg13g2_dlygate4sd3_1 hold1319 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][31] ),
    .X(net3916));
 sg13g2_dlygate4sd3_1 hold1320 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][30] ),
    .X(net3917));
 sg13g2_dlygate4sd3_1 hold1321 (.A(\gpio_uo_out[4] ),
    .X(net3918));
 sg13g2_dlygate4sd3_1 hold1322 (.A(_01791_),
    .X(net3919));
 sg13g2_dlygate4sd3_1 hold1323 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[1][16] ),
    .X(net3920));
 sg13g2_dlygate4sd3_1 hold1324 (.A(\soc_I.rx_uart_i.fifo_i.ram[4][5] ),
    .X(net3921));
 sg13g2_dlygate4sd3_1 hold1325 (.A(_00335_),
    .X(net3922));
 sg13g2_dlygate4sd3_1 hold1326 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[6] ),
    .X(net3923));
 sg13g2_dlygate4sd3_1 hold1327 (.A(_04459_),
    .X(net3924));
 sg13g2_dlygate4sd3_1 hold1328 (.A(_01009_),
    .X(net3925));
 sg13g2_dlygate4sd3_1 hold1329 (.A(\soc_I.rx_uart_i.fifo_i.rd_ptr[0] ),
    .X(net3926));
 sg13g2_dlygate4sd3_1 hold1330 (.A(\soc_I.tx_uart_i.return_state[0] ),
    .X(net3927));
 sg13g2_dlygate4sd3_1 hold1331 (.A(_02138_),
    .X(net3928));
 sg13g2_dlygate4sd3_1 hold1332 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][28] ),
    .X(net3929));
 sg13g2_dlygate4sd3_1 hold1333 (.A(\soc_I.tx_uart_i.wait_states[9] ),
    .X(net3930));
 sg13g2_dlygate4sd3_1 hold1334 (.A(_01932_),
    .X(net3931));
 sg13g2_dlygate4sd3_1 hold1335 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][25] ),
    .X(net3932));
 sg13g2_dlygate4sd3_1 hold1336 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[18] ),
    .X(net3933));
 sg13g2_dlygate4sd3_1 hold1337 (.A(_05551_),
    .X(net3934));
 sg13g2_dlygate4sd3_1 hold1338 (.A(_01283_),
    .X(net3935));
 sg13g2_dlygate4sd3_1 hold1339 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][30] ),
    .X(net3936));
 sg13g2_dlygate4sd3_1 hold1340 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[21][26] ),
    .X(net3937));
 sg13g2_dlygate4sd3_1 hold1341 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[31] ),
    .X(net3938));
 sg13g2_dlygate4sd3_1 hold1342 (.A(\soc_I.rx_uart_i.fifo_i.ram[9][4] ),
    .X(net3939));
 sg13g2_dlygate4sd3_1 hold1343 (.A(_01888_),
    .X(net3940));
 sg13g2_dlygate4sd3_1 hold1344 (.A(\soc_I.rx_uart_i.fifo_i.ram[4][2] ),
    .X(net3941));
 sg13g2_dlygate4sd3_1 hold1345 (.A(_00332_),
    .X(net3942));
 sg13g2_dlygate4sd3_1 hold1346 (.A(\soc_I.clint_I.mtime[19] ),
    .X(net3943));
 sg13g2_dlygate4sd3_1 hold1347 (.A(_01651_),
    .X(net3944));
 sg13g2_dlygate4sd3_1 hold1348 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][23] ),
    .X(net3945));
 sg13g2_dlygate4sd3_1 hold1349 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][13] ),
    .X(net3946));
 sg13g2_dlygate4sd3_1 hold1350 (.A(\soc_I.spi0_I.spi_buf[2] ),
    .X(net3947));
 sg13g2_dlygate4sd3_1 hold1351 (.A(_01973_),
    .X(net3948));
 sg13g2_dlygate4sd3_1 hold1352 (.A(\soc_I.rx_uart_i.fifo_i.ram[5][5] ),
    .X(net3949));
 sg13g2_dlygate4sd3_1 hold1353 (.A(_02300_),
    .X(net3950));
 sg13g2_dlygate4sd3_1 hold1354 (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[11] ),
    .X(net3951));
 sg13g2_dlygate4sd3_1 hold1355 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][18] ),
    .X(net3952));
 sg13g2_dlygate4sd3_1 hold1356 (.A(\soc_I.rx_uart_i.fifo_i.wr_ptr[1] ),
    .X(net3953));
 sg13g2_dlygate4sd3_1 hold1357 (.A(_06948_),
    .X(net3954));
 sg13g2_dlygate4sd3_1 hold1358 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][14] ),
    .X(net3955));
 sg13g2_dlygate4sd3_1 hold1359 (.A(\soc_I.rx_uart_i.fifo_i.ram[6][2] ),
    .X(net3956));
 sg13g2_dlygate4sd3_1 hold1360 (.A(_02289_),
    .X(net3957));
 sg13g2_dlygate4sd3_1 hold1361 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][16] ),
    .X(net3958));
 sg13g2_dlygate4sd3_1 hold1362 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][11] ),
    .X(net3959));
 sg13g2_dlygate4sd3_1 hold1363 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][27] ),
    .X(net3960));
 sg13g2_dlygate4sd3_1 hold1364 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][21] ),
    .X(net3961));
 sg13g2_dlygate4sd3_1 hold1365 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[23] ),
    .X(net3962));
 sg13g2_dlygate4sd3_1 hold1366 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[24][18] ),
    .X(net3963));
 sg13g2_dlygate4sd3_1 hold1367 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[7] ),
    .X(net3964));
 sg13g2_dlygate4sd3_1 hold1368 (.A(\soc_I.rx_uart_i.fifo_i.ram[11][7] ),
    .X(net3965));
 sg13g2_dlygate4sd3_1 hold1369 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[8] ),
    .X(net3966));
 sg13g2_dlygate4sd3_1 hold1370 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[11] ),
    .X(net3967));
 sg13g2_dlygate4sd3_1 hold1371 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[21] ),
    .X(net3968));
 sg13g2_dlygate4sd3_1 hold1372 (.A(_04518_),
    .X(net3969));
 sg13g2_dlygate4sd3_1 hold1373 (.A(_01024_),
    .X(net3970));
 sg13g2_dlygate4sd3_1 hold1374 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[7] ),
    .X(net3971));
 sg13g2_dlygate4sd3_1 hold1375 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][1] ),
    .X(net3972));
 sg13g2_dlygate4sd3_1 hold1376 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][12] ),
    .X(net3973));
 sg13g2_dlygate4sd3_1 hold1377 (.A(\soc_I.rx_uart_i.fifo_i.ram[15][7] ),
    .X(net3974));
 sg13g2_dlygate4sd3_1 hold1378 (.A(_01104_),
    .X(net3975));
 sg13g2_dlygate4sd3_1 hold1379 (.A(\soc_I.qqspi_I.rdata[10] ),
    .X(net3976));
 sg13g2_dlygate4sd3_1 hold1380 (.A(_01806_),
    .X(net3977));
 sg13g2_dlygate4sd3_1 hold1381 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.bit_idx[2] ),
    .X(net3978));
 sg13g2_dlygate4sd3_1 hold1382 (.A(_01331_),
    .X(net3979));
 sg13g2_dlygate4sd3_1 hold1383 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][2] ),
    .X(net3980));
 sg13g2_dlygate4sd3_1 hold1384 (.A(\soc_I.rx_uart_i.fifo_i.din[2] ),
    .X(net3981));
 sg13g2_dlygate4sd3_1 hold1385 (.A(_00632_),
    .X(net3982));
 sg13g2_dlygate4sd3_1 hold1386 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][9] ),
    .X(net3983));
 sg13g2_dlygate4sd3_1 hold1387 (.A(\soc_I.rx_uart_i.fifo_i.ram[14][0] ),
    .X(net3984));
 sg13g2_dlygate4sd3_1 hold1388 (.A(_02814_),
    .X(net3985));
 sg13g2_dlygate4sd3_1 hold1389 (.A(_00670_),
    .X(net3986));
 sg13g2_dlygate4sd3_1 hold1390 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][18] ),
    .X(net3987));
 sg13g2_dlygate4sd3_1 hold1391 (.A(\soc_I.rx_uart_i.fifo_i.ram[2][4] ),
    .X(net3988));
 sg13g2_dlygate4sd3_1 hold1392 (.A(_01085_),
    .X(net3989));
 sg13g2_dlygate4sd3_1 hold1393 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][27] ),
    .X(net3990));
 sg13g2_dlygate4sd3_1 hold1394 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][0] ),
    .X(net3991));
 sg13g2_dlygate4sd3_1 hold1395 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][24] ),
    .X(net3992));
 sg13g2_dlygate4sd3_1 hold1396 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[7] ),
    .X(net3993));
 sg13g2_dlygate4sd3_1 hold1397 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][30] ),
    .X(net3994));
 sg13g2_dlygate4sd3_1 hold1398 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][24] ),
    .X(net3995));
 sg13g2_dlygate4sd3_1 hold1399 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[19] ),
    .X(net3996));
 sg13g2_dlygate4sd3_1 hold1400 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][19] ),
    .X(net3997));
 sg13g2_dlygate4sd3_1 hold1401 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][10] ),
    .X(net3998));
 sg13g2_dlygate4sd3_1 hold1402 (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[0] ),
    .X(net3999));
 sg13g2_dlygate4sd3_1 hold1403 (.A(_04122_),
    .X(net4000));
 sg13g2_dlygate4sd3_1 hold1404 (.A(\soc_I.clint_I.mtime[47] ),
    .X(net4001));
 sg13g2_dlygate4sd3_1 hold1405 (.A(_06410_),
    .X(net4002));
 sg13g2_dlygate4sd3_1 hold1406 (.A(\soc_I.rx_uart_i.fifo_i.ram[3][4] ),
    .X(net4003));
 sg13g2_dlygate4sd3_1 hold1407 (.A(_01077_),
    .X(net4004));
 sg13g2_dlygate4sd3_1 hold1408 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][4] ),
    .X(net4005));
 sg13g2_dlygate4sd3_1 hold1409 (.A(\soc_I.rx_uart_i.fifo_i.ram[8][2] ),
    .X(net4006));
 sg13g2_dlygate4sd3_1 hold1410 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[23][28] ),
    .X(net4007));
 sg13g2_dlygate4sd3_1 hold1411 (.A(\soc_I.spi0_I.spi_buf[4] ),
    .X(net4008));
 sg13g2_dlygate4sd3_1 hold1412 (.A(_01975_),
    .X(net4009));
 sg13g2_dlygate4sd3_1 hold1413 (.A(\soc_I.rx_uart_i.fifo_i.ram[6][4] ),
    .X(net4010));
 sg13g2_dlygate4sd3_1 hold1414 (.A(_02291_),
    .X(net4011));
 sg13g2_dlygate4sd3_1 hold1415 (.A(_00292_),
    .X(net4012));
 sg13g2_dlygate4sd3_1 hold1416 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][11] ),
    .X(net4013));
 sg13g2_dlygate4sd3_1 hold1417 (.A(\soc_I.rx_uart_i.fifo_i.ram[6][5] ),
    .X(net4014));
 sg13g2_dlygate4sd3_1 hold1418 (.A(_02292_),
    .X(net4015));
 sg13g2_dlygate4sd3_1 hold1419 (.A(\soc_I.rx_uart_i.fifo_i.ram[7][4] ),
    .X(net4016));
 sg13g2_dlygate4sd3_1 hold1420 (.A(_02283_),
    .X(net4017));
 sg13g2_dlygate4sd3_1 hold1421 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][5] ),
    .X(net4018));
 sg13g2_dlygate4sd3_1 hold1422 (.A(\soc_I.rx_uart_i.fifo_i.ram[1][2] ),
    .X(net4019));
 sg13g2_dlygate4sd3_1 hold1423 (.A(\soc_I.tx_uart_i.wait_states[1] ),
    .X(net4020));
 sg13g2_dlygate4sd3_1 hold1424 (.A(_01924_),
    .X(net4021));
 sg13g2_dlygate4sd3_1 hold1425 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][12] ),
    .X(net4022));
 sg13g2_dlygate4sd3_1 hold1426 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[20][11] ),
    .X(net4023));
 sg13g2_dlygate4sd3_1 hold1427 (.A(\soc_I.rx_uart_i.fifo_i.ram[0][5] ),
    .X(net4024));
 sg13g2_dlygate4sd3_1 hold1428 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][3] ),
    .X(net4025));
 sg13g2_dlygate4sd3_1 hold1429 (.A(\soc_I.rx_uart_i.fifo_i.ram[1][3] ),
    .X(net4026));
 sg13g2_dlygate4sd3_1 hold1430 (.A(_01092_),
    .X(net4027));
 sg13g2_dlygate4sd3_1 hold1431 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[63] ),
    .X(net4028));
 sg13g2_dlygate4sd3_1 hold1432 (.A(_01200_),
    .X(net4029));
 sg13g2_dlygate4sd3_1 hold1433 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][1] ),
    .X(net4030));
 sg13g2_dlygate4sd3_1 hold1434 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][30] ),
    .X(net4031));
 sg13g2_dlygate4sd3_1 hold1435 (.A(_00152_),
    .X(net4032));
 sg13g2_dlygate4sd3_1 hold1436 (.A(_07469_),
    .X(net4033));
 sg13g2_dlygate4sd3_1 hold1437 (.A(\soc_I.rx_uart_i.fifo_i.ram[1][1] ),
    .X(net4034));
 sg13g2_dlygate4sd3_1 hold1438 (.A(_01090_),
    .X(net4035));
 sg13g2_dlygate4sd3_1 hold1439 (.A(\soc_I.rx_uart_i.fifo_i.ram[5][7] ),
    .X(net4036));
 sg13g2_dlygate4sd3_1 hold1440 (.A(\soc_I.rx_uart_i.fifo_i.ram[7][5] ),
    .X(net4037));
 sg13g2_dlygate4sd3_1 hold1441 (.A(_02284_),
    .X(net4038));
 sg13g2_dlygate4sd3_1 hold1442 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[6] ),
    .X(net4039));
 sg13g2_dlygate4sd3_1 hold1443 (.A(\soc_I.rx_uart_i.fifo_i.ram[5][4] ),
    .X(net4040));
 sg13g2_dlygate4sd3_1 hold1444 (.A(_02299_),
    .X(net4041));
 sg13g2_dlygate4sd3_1 hold1445 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][1] ),
    .X(net4042));
 sg13g2_dlygate4sd3_1 hold1446 (.A(\soc_I.rx_uart_i.fifo_i.ram[15][6] ),
    .X(net4043));
 sg13g2_dlygate4sd3_1 hold1447 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[7][11] ),
    .X(net4044));
 sg13g2_dlygate4sd3_1 hold1448 (.A(\soc_I.tx_uart_i.tx_data_reg[4] ),
    .X(net4045));
 sg13g2_dlygate4sd3_1 hold1449 (.A(_01880_),
    .X(net4046));
 sg13g2_dlygate4sd3_1 hold1450 (.A(\soc_I.rx_uart_i.fifo_i.ram[0][7] ),
    .X(net4047));
 sg13g2_dlygate4sd3_1 hold1451 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][14] ),
    .X(net4048));
 sg13g2_dlygate4sd3_1 hold1452 (.A(\soc_I.rx_uart_i.fifo_i.ram[12][1] ),
    .X(net4049));
 sg13g2_dlygate4sd3_1 hold1453 (.A(\soc_I.rx_uart_i.fifo_i.ram[11][2] ),
    .X(net4050));
 sg13g2_dlygate4sd3_1 hold1454 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[11][18] ),
    .X(net4051));
 sg13g2_dlygate4sd3_1 hold1455 (.A(\soc_I.rx_uart_i.fifo_i.ram[3][7] ),
    .X(net4052));
 sg13g2_dlygate4sd3_1 hold1456 (.A(\soc_I.rx_uart_i.fifo_i.ram[6][3] ),
    .X(net4053));
 sg13g2_dlygate4sd3_1 hold1457 (.A(_02290_),
    .X(net4054));
 sg13g2_dlygate4sd3_1 hold1458 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[10] ),
    .X(net4055));
 sg13g2_dlygate4sd3_1 hold1459 (.A(_04474_),
    .X(net4056));
 sg13g2_dlygate4sd3_1 hold1460 (.A(_01013_),
    .X(net4057));
 sg13g2_dlygate4sd3_1 hold1461 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[43] ),
    .X(net4058));
 sg13g2_dlygate4sd3_1 hold1462 (.A(_04759_),
    .X(net4059));
 sg13g2_dlygate4sd3_1 hold1463 (.A(_01180_),
    .X(net4060));
 sg13g2_dlygate4sd3_1 hold1464 (.A(\gpio_uo_out[7] ),
    .X(net4061));
 sg13g2_dlygate4sd3_1 hold1465 (.A(_01794_),
    .X(net4062));
 sg13g2_dlygate4sd3_1 hold1466 (.A(\soc_I.rx_uart_i.fifo_i.ram[2][5] ),
    .X(net4063));
 sg13g2_dlygate4sd3_1 hold1467 (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[14] ),
    .X(net4064));
 sg13g2_dlygate4sd3_1 hold1468 (.A(\soc_I.rx_uart_i.fifo_i.ram[1][7] ),
    .X(net4065));
 sg13g2_dlygate4sd3_1 hold1469 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][4] ),
    .X(net4066));
 sg13g2_dlygate4sd3_1 hold1470 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][23] ),
    .X(net4067));
 sg13g2_dlygate4sd3_1 hold1471 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[30] ),
    .X(net4068));
 sg13g2_dlygate4sd3_1 hold1472 (.A(\soc_I.qqspi_I.state[2] ),
    .X(net4069));
 sg13g2_dlygate4sd3_1 hold1473 (.A(_12567_),
    .X(net4070));
 sg13g2_dlygate4sd3_1 hold1474 (.A(\soc_I.rx_uart_i.fifo_i.ram[3][2] ),
    .X(net4071));
 sg13g2_dlygate4sd3_1 hold1475 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][4] ),
    .X(net4072));
 sg13g2_dlygate4sd3_1 hold1476 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[12][16] ),
    .X(net4073));
 sg13g2_dlygate4sd3_1 hold1477 (.A(\soc_I.rx_uart_i.fifo_i.ram[4][3] ),
    .X(net4074));
 sg13g2_dlygate4sd3_1 hold1478 (.A(_00333_),
    .X(net4075));
 sg13g2_dlygate4sd3_1 hold1479 (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[30] ),
    .X(net4076));
 sg13g2_dlygate4sd3_1 hold1480 (.A(\soc_I.rx_uart_i.fifo_i.ram[10][7] ),
    .X(net4077));
 sg13g2_dlygate4sd3_1 hold1481 (.A(_00645_),
    .X(net4078));
 sg13g2_dlygate4sd3_1 hold1482 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[29] ),
    .X(net4079));
 sg13g2_dlygate4sd3_1 hold1483 (.A(_00178_),
    .X(net4080));
 sg13g2_dlygate4sd3_1 hold1484 (.A(_05373_),
    .X(net4081));
 sg13g2_dlygate4sd3_1 hold1485 (.A(\soc_I.rx_uart_i.fifo_i.ram[4][4] ),
    .X(net4082));
 sg13g2_dlygate4sd3_1 hold1486 (.A(_00334_),
    .X(net4083));
 sg13g2_dlygate4sd3_1 hold1487 (.A(\soc_I.rx_uart_i.fifo_i.ram[2][6] ),
    .X(net4084));
 sg13g2_dlygate4sd3_1 hold1488 (.A(_01087_),
    .X(net4085));
 sg13g2_dlygate4sd3_1 hold1489 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[25] ),
    .X(net4086));
 sg13g2_dlygate4sd3_1 hold1490 (.A(_04534_),
    .X(net4087));
 sg13g2_dlygate4sd3_1 hold1491 (.A(_01028_),
    .X(net4088));
 sg13g2_dlygate4sd3_1 hold1492 (.A(\soc_I.rx_uart_i.fifo_i.ram[15][4] ),
    .X(net4089));
 sg13g2_dlygate4sd3_1 hold1493 (.A(_01101_),
    .X(net4090));
 sg13g2_dlygate4sd3_1 hold1494 (.A(\soc_I.rx_uart_i.fifo_i.ram[6][1] ),
    .X(net4091));
 sg13g2_dlygate4sd3_1 hold1495 (.A(\soc_I.rx_uart_i.fifo_i.ram[15][3] ),
    .X(net4092));
 sg13g2_dlygate4sd3_1 hold1496 (.A(_01100_),
    .X(net4093));
 sg13g2_dlygate4sd3_1 hold1497 (.A(\soc_I.rx_uart_i.fifo_i.ram[1][4] ),
    .X(net4094));
 sg13g2_dlygate4sd3_1 hold1498 (.A(_01093_),
    .X(net4095));
 sg13g2_dlygate4sd3_1 hold1499 (.A(\soc_I.rx_uart_i.fifo_i.ram[2][1] ),
    .X(net4096));
 sg13g2_dlygate4sd3_1 hold1500 (.A(_01082_),
    .X(net4097));
 sg13g2_dlygate4sd3_1 hold1501 (.A(\soc_I.rx_uart_i.fifo_i.ram[15][1] ),
    .X(net4098));
 sg13g2_dlygate4sd3_1 hold1502 (.A(\soc_I.rx_uart_i.fifo_i.ram[11][5] ),
    .X(net4099));
 sg13g2_dlygate4sd3_1 hold1503 (.A(_00651_),
    .X(net4100));
 sg13g2_dlygate4sd3_1 hold1504 (.A(\soc_I.rx_uart_i.fifo_i.ram[5][6] ),
    .X(net4101));
 sg13g2_dlygate4sd3_1 hold1505 (.A(\soc_I.spi0_I.spi_buf[5] ),
    .X(net4102));
 sg13g2_dlygate4sd3_1 hold1506 (.A(_01976_),
    .X(net4103));
 sg13g2_dlygate4sd3_1 hold1507 (.A(\soc_I.rx_uart_i.fifo_i.ram[10][6] ),
    .X(net4104));
 sg13g2_dlygate4sd3_1 hold1508 (.A(_00644_),
    .X(net4105));
 sg13g2_dlygate4sd3_1 hold1509 (.A(\soc_I.rx_uart_i.fifo_i.ram[7][6] ),
    .X(net4106));
 sg13g2_dlygate4sd3_1 hold1510 (.A(\soc_I.rx_uart_i.fifo_i.ram[7][2] ),
    .X(net4107));
 sg13g2_dlygate4sd3_1 hold1511 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][3] ),
    .X(net4108));
 sg13g2_dlygate4sd3_1 hold1512 (.A(\soc_I.rx_uart_i.fifo_i.ram[12][4] ),
    .X(net4109));
 sg13g2_dlygate4sd3_1 hold1513 (.A(_00658_),
    .X(net4110));
 sg13g2_dlygate4sd3_1 hold1514 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[10][7] ),
    .X(net4111));
 sg13g2_dlygate4sd3_1 hold1515 (.A(\soc_I.rx_uart_i.fifo_i.ram[7][7] ),
    .X(net4112));
 sg13g2_dlygate4sd3_1 hold1516 (.A(_02286_),
    .X(net4113));
 sg13g2_dlygate4sd3_1 hold1517 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[9] ),
    .X(net4114));
 sg13g2_dlygate4sd3_1 hold1518 (.A(_04677_),
    .X(net4115));
 sg13g2_dlygate4sd3_1 hold1519 (.A(_01146_),
    .X(net4116));
 sg13g2_dlygate4sd3_1 hold1520 (.A(\soc_I.tx_uart_i.wait_states[0] ),
    .X(net4117));
 sg13g2_dlygate4sd3_1 hold1521 (.A(\soc_I.kianv_I.Instr[1] ),
    .X(net4118));
 sg13g2_dlygate4sd3_1 hold1522 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[24] ),
    .X(net4119));
 sg13g2_dlygate4sd3_1 hold1523 (.A(_04530_),
    .X(net4120));
 sg13g2_dlygate4sd3_1 hold1524 (.A(_01027_),
    .X(net4121));
 sg13g2_dlygate4sd3_1 hold1525 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][21] ),
    .X(net4122));
 sg13g2_dlygate4sd3_1 hold1526 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[13] ),
    .X(net4123));
 sg13g2_dlygate4sd3_1 hold1527 (.A(_04486_),
    .X(net4124));
 sg13g2_dlygate4sd3_1 hold1528 (.A(_01016_),
    .X(net4125));
 sg13g2_dlygate4sd3_1 hold1529 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[29] ),
    .X(net4126));
 sg13g2_dlygate4sd3_1 hold1530 (.A(\soc_I.rx_uart_i.fifo_i.ram[0][6] ),
    .X(net4127));
 sg13g2_dlygate4sd3_1 hold1531 (.A(_00636_),
    .X(net4128));
 sg13g2_dlygate4sd3_1 hold1532 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[2] ),
    .X(net4129));
 sg13g2_dlygate4sd3_1 hold1533 (.A(_01139_),
    .X(net4130));
 sg13g2_dlygate4sd3_1 hold1534 (.A(\soc_I.rx_uart_i.fifo_i.ram[1][6] ),
    .X(net4131));
 sg13g2_dlygate4sd3_1 hold1535 (.A(_01095_),
    .X(net4132));
 sg13g2_dlygate4sd3_1 hold1536 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[12] ),
    .X(net4133));
 sg13g2_dlygate4sd3_1 hold1537 (.A(_04482_),
    .X(net4134));
 sg13g2_dlygate4sd3_1 hold1538 (.A(_01015_),
    .X(net4135));
 sg13g2_dlygate4sd3_1 hold1539 (.A(\soc_I.rx_uart_i.fifo_i.ram[4][1] ),
    .X(net4136));
 sg13g2_dlygate4sd3_1 hold1540 (.A(_00331_),
    .X(net4137));
 sg13g2_dlygate4sd3_1 hold1541 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[20] ),
    .X(net4138));
 sg13g2_dlygate4sd3_1 hold1542 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[15] ),
    .X(net4139));
 sg13g2_dlygate4sd3_1 hold1543 (.A(_04494_),
    .X(net4140));
 sg13g2_dlygate4sd3_1 hold1544 (.A(_01018_),
    .X(net4141));
 sg13g2_dlygate4sd3_1 hold1545 (.A(\soc_I.rx_uart_i.fifo_i.ram[0][3] ),
    .X(net4142));
 sg13g2_dlygate4sd3_1 hold1546 (.A(_00633_),
    .X(net4143));
 sg13g2_dlygate4sd3_1 hold1547 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[3] ),
    .X(net4144));
 sg13g2_dlygate4sd3_1 hold1548 (.A(_01006_),
    .X(net4145));
 sg13g2_dlygate4sd3_1 hold1549 (.A(\soc_I.rx_uart_i.fifo_i.ram[8][1] ),
    .X(net4146));
 sg13g2_dlygate4sd3_1 hold1550 (.A(_02101_),
    .X(net4147));
 sg13g2_dlygate4sd3_1 hold1551 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[55] ),
    .X(net4148));
 sg13g2_dlygate4sd3_1 hold1552 (.A(_05613_),
    .X(net4149));
 sg13g2_dlygate4sd3_1 hold1553 (.A(\soc_I.rx_uart_i.fifo_i.ram[9][6] ),
    .X(net4150));
 sg13g2_dlygate4sd3_1 hold1554 (.A(_01890_),
    .X(net4151));
 sg13g2_dlygate4sd3_1 hold1555 (.A(\soc_I.rx_uart_i.fifo_i.ram[2][3] ),
    .X(net4152));
 sg13g2_dlygate4sd3_1 hold1556 (.A(_01084_),
    .X(net4153));
 sg13g2_dlygate4sd3_1 hold1557 (.A(\soc_I.rx_uart_i.fifo_i.ram[12][7] ),
    .X(net4154));
 sg13g2_dlygate4sd3_1 hold1558 (.A(\soc_I.clint_I.tick_cnt[12] ),
    .X(net4155));
 sg13g2_dlygate4sd3_1 hold1559 (.A(_06244_),
    .X(net4156));
 sg13g2_dlygate4sd3_1 hold1560 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[4][24] ),
    .X(net4157));
 sg13g2_dlygate4sd3_1 hold1561 (.A(\soc_I.rx_uart_i.fifo_i.ram[3][3] ),
    .X(net4158));
 sg13g2_dlygate4sd3_1 hold1562 (.A(_01076_),
    .X(net4159));
 sg13g2_dlygate4sd3_1 hold1563 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[10] ),
    .X(net4160));
 sg13g2_dlygate4sd3_1 hold1564 (.A(\soc_I.rx_uart_i.fifo_i.ram[10][3] ),
    .X(net4161));
 sg13g2_dlygate4sd3_1 hold1565 (.A(_00641_),
    .X(net4162));
 sg13g2_dlygate4sd3_1 hold1566 (.A(\soc_I.rx_uart_i.fifo_i.ram[2][7] ),
    .X(net4163));
 sg13g2_dlygate4sd3_1 hold1567 (.A(_00149_),
    .X(net4164));
 sg13g2_dlygate4sd3_1 hold1568 (.A(_01782_),
    .X(net4165));
 sg13g2_dlygate4sd3_1 hold1569 (.A(\soc_I.qqspi_I.rdata[14] ),
    .X(net4166));
 sg13g2_dlygate4sd3_1 hold1570 (.A(_01810_),
    .X(net4167));
 sg13g2_dlygate4sd3_1 hold1571 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[43] ),
    .X(net4168));
 sg13g2_dlygate4sd3_1 hold1572 (.A(_05593_),
    .X(net4169));
 sg13g2_dlygate4sd3_1 hold1573 (.A(\soc_I.rx_uart_i.fifo_i.ram[1][5] ),
    .X(net4170));
 sg13g2_dlygate4sd3_1 hold1574 (.A(_00018_),
    .X(net4171));
 sg13g2_dlygate4sd3_1 hold1575 (.A(_06356_),
    .X(net4172));
 sg13g2_dlygate4sd3_1 hold1576 (.A(_01657_),
    .X(net4173));
 sg13g2_dlygate4sd3_1 hold1577 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[3][8] ),
    .X(net4174));
 sg13g2_dlygate4sd3_1 hold1578 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[28][30] ),
    .X(net4175));
 sg13g2_dlygate4sd3_1 hold1579 (.A(\soc_I.rx_uart_i.fifo_i.ram[9][7] ),
    .X(net4176));
 sg13g2_dlygate4sd3_1 hold1580 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[11] ),
    .X(net4177));
 sg13g2_dlygate4sd3_1 hold1581 (.A(_04478_),
    .X(net4178));
 sg13g2_dlygate4sd3_1 hold1582 (.A(_01014_),
    .X(net4179));
 sg13g2_dlygate4sd3_1 hold1583 (.A(\soc_I.rx_uart_i.fifo_i.ram[3][1] ),
    .X(net4180));
 sg13g2_dlygate4sd3_1 hold1584 (.A(_01074_),
    .X(net4181));
 sg13g2_dlygate4sd3_1 hold1585 (.A(\soc_I.rx_uart_i.fifo_i.ram[4][7] ),
    .X(net4182));
 sg13g2_dlygate4sd3_1 hold1586 (.A(_00337_),
    .X(net4183));
 sg13g2_dlygate4sd3_1 hold1587 (.A(\soc_I.rx_uart_i.fifo_i.ram[9][1] ),
    .X(net4184));
 sg13g2_dlygate4sd3_1 hold1588 (.A(_01885_),
    .X(net4185));
 sg13g2_dlygate4sd3_1 hold1589 (.A(\soc_I.rx_uart_i.fifo_i.ram[15][5] ),
    .X(net4186));
 sg13g2_dlygate4sd3_1 hold1590 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][4] ),
    .X(net4187));
 sg13g2_dlygate4sd3_1 hold1591 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[27] ),
    .X(net4188));
 sg13g2_dlygate4sd3_1 hold1592 (.A(\soc_I.spi0_I.tick_cnt[10] ),
    .X(net4189));
 sg13g2_dlygate4sd3_1 hold1593 (.A(_06629_),
    .X(net4190));
 sg13g2_dlygate4sd3_1 hold1594 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[27][7] ),
    .X(net4191));
 sg13g2_dlygate4sd3_1 hold1595 (.A(\soc_I.rx_uart_i.fifo_i.ram[12][3] ),
    .X(net4192));
 sg13g2_dlygate4sd3_1 hold1596 (.A(_00657_),
    .X(net4193));
 sg13g2_dlygate4sd3_1 hold1597 (.A(\soc_I.rx_uart_i.fifo_i.ram[2][2] ),
    .X(net4194));
 sg13g2_dlygate4sd3_1 hold1598 (.A(\soc_I.tx_uart_i.wait_states[13] ),
    .X(net4195));
 sg13g2_dlygate4sd3_1 hold1599 (.A(_01936_),
    .X(net4196));
 sg13g2_dlygate4sd3_1 hold1600 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[7] ),
    .X(net4197));
 sg13g2_dlygate4sd3_1 hold1601 (.A(\soc_I.rx_uart_i.fifo_i.ram[5][1] ),
    .X(net4198));
 sg13g2_dlygate4sd3_1 hold1602 (.A(\soc_I.rx_uart_i.fifo_i.ram[9][2] ),
    .X(net4199));
 sg13g2_dlygate4sd3_1 hold1603 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[19][16] ),
    .X(net4200));
 sg13g2_dlygate4sd3_1 hold1604 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[31] ),
    .X(net4201));
 sg13g2_dlygate4sd3_1 hold1605 (.A(_05573_),
    .X(net4202));
 sg13g2_dlygate4sd3_1 hold1606 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[16] ),
    .X(net4203));
 sg13g2_dlygate4sd3_1 hold1607 (.A(_04498_),
    .X(net4204));
 sg13g2_dlygate4sd3_1 hold1608 (.A(_01019_),
    .X(net4205));
 sg13g2_dlygate4sd3_1 hold1609 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][8] ),
    .X(net4206));
 sg13g2_dlygate4sd3_1 hold1610 (.A(\soc_I.rx_uart_i.fifo_i.ram[3][6] ),
    .X(net4207));
 sg13g2_dlygate4sd3_1 hold1611 (.A(_01079_),
    .X(net4208));
 sg13g2_dlygate4sd3_1 hold1612 (.A(\soc_I.rx_uart_i.fifo_i.ram[8][4] ),
    .X(net4209));
 sg13g2_dlygate4sd3_1 hold1613 (.A(_02104_),
    .X(net4210));
 sg13g2_dlygate4sd3_1 hold1614 (.A(\soc_I.rx_uart_i.fifo_i.ram[7][1] ),
    .X(net4211));
 sg13g2_dlygate4sd3_1 hold1615 (.A(\soc_I.rx_uart_i.fifo_i.ram[11][1] ),
    .X(net4212));
 sg13g2_dlygate4sd3_1 hold1616 (.A(_00647_),
    .X(net4213));
 sg13g2_dlygate4sd3_1 hold1617 (.A(\soc_I.rx_uart_i.fifo_i.ram[0][4] ),
    .X(net4214));
 sg13g2_dlygate4sd3_1 hold1618 (.A(_00634_),
    .X(net4215));
 sg13g2_dlygate4sd3_1 hold1619 (.A(\soc_I.gpio0_I.rdata[0] ),
    .X(net4216));
 sg13g2_dlygate4sd3_1 hold1620 (.A(_01787_),
    .X(net4217));
 sg13g2_dlygate4sd3_1 hold1621 (.A(\soc_I.rx_uart_i.fifo_i.ram[6][6] ),
    .X(net4218));
 sg13g2_dlygate4sd3_1 hold1622 (.A(\soc_I.rx_uart_i.fifo_i.ram[11][4] ),
    .X(net4219));
 sg13g2_dlygate4sd3_1 hold1623 (.A(_00650_),
    .X(net4220));
 sg13g2_dlygate4sd3_1 hold1624 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[7] ),
    .X(net4221));
 sg13g2_dlygate4sd3_1 hold1625 (.A(_01068_),
    .X(net4222));
 sg13g2_dlygate4sd3_1 hold1626 (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[12] ),
    .X(net4223));
 sg13g2_dlygate4sd3_1 hold1627 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][11] ),
    .X(net4224));
 sg13g2_dlygate4sd3_1 hold1628 (.A(\soc_I.clint_I.mtimecmp[19] ),
    .X(net4225));
 sg13g2_dlygate4sd3_1 hold1629 (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[15] ),
    .X(net4226));
 sg13g2_dlygate4sd3_1 hold1630 (.A(_01454_),
    .X(net4227));
 sg13g2_dlygate4sd3_1 hold1631 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[7] ),
    .X(net4228));
 sg13g2_dlygate4sd3_1 hold1632 (.A(_04462_),
    .X(net4229));
 sg13g2_dlygate4sd3_1 hold1633 (.A(_01010_),
    .X(net4230));
 sg13g2_dlygate4sd3_1 hold1634 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[1] ),
    .X(net4231));
 sg13g2_dlygate4sd3_1 hold1635 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[20] ),
    .X(net4232));
 sg13g2_dlygate4sd3_1 hold1636 (.A(_04514_),
    .X(net4233));
 sg13g2_dlygate4sd3_1 hold1637 (.A(_01023_),
    .X(net4234));
 sg13g2_dlygate4sd3_1 hold1638 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[19] ),
    .X(net4235));
 sg13g2_dlygate4sd3_1 hold1639 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[15][27] ),
    .X(net4236));
 sg13g2_dlygate4sd3_1 hold1640 (.A(\soc_I.rx_uart_i.fifo_i.ram[11][6] ),
    .X(net4237));
 sg13g2_dlygate4sd3_1 hold1641 (.A(_00652_),
    .X(net4238));
 sg13g2_dlygate4sd3_1 hold1642 (.A(\soc_I.tx_uart_i.wait_states[4] ),
    .X(net4239));
 sg13g2_dlygate4sd3_1 hold1643 (.A(\soc_I.rx_uart_i.fifo_i.ram[12][6] ),
    .X(net4240));
 sg13g2_dlygate4sd3_1 hold1644 (.A(\soc_I.PC[3] ),
    .X(net4241));
 sg13g2_dlygate4sd3_1 hold1645 (.A(\soc_I.PC[30] ),
    .X(net4242));
 sg13g2_dlygate4sd3_1 hold1646 (.A(_01469_),
    .X(net4243));
 sg13g2_dlygate4sd3_1 hold1647 (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[6] ),
    .X(net4244));
 sg13g2_dlygate4sd3_1 hold1648 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[17] ),
    .X(net4245));
 sg13g2_dlygate4sd3_1 hold1649 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[17] ),
    .X(net4246));
 sg13g2_dlygate4sd3_1 hold1650 (.A(_04502_),
    .X(net4247));
 sg13g2_dlygate4sd3_1 hold1651 (.A(_01020_),
    .X(net4248));
 sg13g2_dlygate4sd3_1 hold1652 (.A(\soc_I.rx_uart_i.fifo_i.cnt[2] ),
    .X(net4249));
 sg13g2_dlygate4sd3_1 hold1653 (.A(\soc_I.rx_uart_i.fifo_i.ram[9][3] ),
    .X(net4250));
 sg13g2_dlygate4sd3_1 hold1654 (.A(\soc_I.spi0_I.tick_cnt[14] ),
    .X(net4251));
 sg13g2_dlygate4sd3_1 hold1655 (.A(_06637_),
    .X(net4252));
 sg13g2_dlygate4sd3_1 hold1656 (.A(\soc_I.rx_uart_i.fifo_i.ram[4][6] ),
    .X(net4253));
 sg13g2_dlygate4sd3_1 hold1657 (.A(\soc_I.rx_uart_i.fifo_i.ram[7][3] ),
    .X(net4254));
 sg13g2_dlygate4sd3_1 hold1658 (.A(_02282_),
    .X(net4255));
 sg13g2_dlygate4sd3_1 hold1659 (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[20] ),
    .X(net4256));
 sg13g2_dlygate4sd3_1 hold1660 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[10] ),
    .X(net4257));
 sg13g2_dlygate4sd3_1 hold1661 (.A(_00850_),
    .X(net4258));
 sg13g2_dlygate4sd3_1 hold1662 (.A(\soc_I.tx_uart_i.wait_states[14] ),
    .X(net4259));
 sg13g2_dlygate4sd3_1 hold1663 (.A(\soc_I.rx_uart_i.fifo_i.ram[5][2] ),
    .X(net4260));
 sg13g2_dlygate4sd3_1 hold1664 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[22] ),
    .X(net4261));
 sg13g2_dlygate4sd3_1 hold1665 (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[5] ),
    .X(net4262));
 sg13g2_dlygate4sd3_1 hold1666 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[26] ),
    .X(net4263));
 sg13g2_dlygate4sd3_1 hold1667 (.A(_04538_),
    .X(net4264));
 sg13g2_dlygate4sd3_1 hold1668 (.A(_01029_),
    .X(net4265));
 sg13g2_dlygate4sd3_1 hold1669 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[20] ),
    .X(net4266));
 sg13g2_dlygate4sd3_1 hold1670 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[5][14] ),
    .X(net4267));
 sg13g2_dlygate4sd3_1 hold1671 (.A(\soc_I.clint_I.mtime[57] ),
    .X(net4268));
 sg13g2_dlygate4sd3_1 hold1672 (.A(_06430_),
    .X(net4269));
 sg13g2_dlygate4sd3_1 hold1673 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[8][2] ),
    .X(net4270));
 sg13g2_dlygate4sd3_1 hold1674 (.A(\soc_I.rx_uart_i.fifo_i.ram[9][5] ),
    .X(net4271));
 sg13g2_dlygate4sd3_1 hold1675 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[14] ),
    .X(net4272));
 sg13g2_dlygate4sd3_1 hold1676 (.A(\soc_I.clint_I.mtimecmp[12] ),
    .X(net4273));
 sg13g2_dlygate4sd3_1 hold1677 (.A(\soc_I.clint_I.mtime[54] ),
    .X(net4274));
 sg13g2_dlygate4sd3_1 hold1678 (.A(_06424_),
    .X(net4275));
 sg13g2_dlygate4sd3_1 hold1679 (.A(_01686_),
    .X(net4276));
 sg13g2_dlygate4sd3_1 hold1680 (.A(\soc_I.gpio0_I.rdata[6] ),
    .X(net4277));
 sg13g2_dlygate4sd3_1 hold1681 (.A(_01793_),
    .X(net4278));
 sg13g2_dlygate4sd3_1 hold1682 (.A(\soc_I.spi0_I.tick_cnt[7] ),
    .X(net4279));
 sg13g2_dlygate4sd3_1 hold1683 (.A(_06623_),
    .X(net4280));
 sg13g2_dlygate4sd3_1 hold1684 (.A(\soc_I.tx_uart_i.ready ),
    .X(net4281));
 sg13g2_dlygate4sd3_1 hold1685 (.A(_06968_),
    .X(net4282));
 sg13g2_dlygate4sd3_1 hold1686 (.A(_01870_),
    .X(net4283));
 sg13g2_dlygate4sd3_1 hold1687 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[1] ),
    .X(net4284));
 sg13g2_dlygate4sd3_1 hold1688 (.A(_01266_),
    .X(net4285));
 sg13g2_dlygate4sd3_1 hold1689 (.A(\soc_I.rx_uart_i.fifo_i.ram[15][2] ),
    .X(net4286));
 sg13g2_dlygate4sd3_1 hold1690 (.A(\soc_I.spi0_I.tick_cnt[9] ),
    .X(net4287));
 sg13g2_dlygate4sd3_1 hold1691 (.A(_06627_),
    .X(net4288));
 sg13g2_dlygate4sd3_1 hold1692 (.A(\soc_I.tx_uart_i.tx_data_reg[1] ),
    .X(net4289));
 sg13g2_dlygate4sd3_1 hold1693 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[23] ),
    .X(net4290));
 sg13g2_dlygate4sd3_1 hold1694 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[1] ),
    .X(net4291));
 sg13g2_dlygate4sd3_1 hold1695 (.A(\soc_I.spi0_I.xfer_cycles[4] ),
    .X(net4292));
 sg13g2_dlygate4sd3_1 hold1696 (.A(_01750_),
    .X(net4293));
 sg13g2_dlygate4sd3_1 hold1697 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[15] ),
    .X(net4294));
 sg13g2_dlygate4sd3_1 hold1698 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[12] ),
    .X(net4295));
 sg13g2_dlygate4sd3_1 hold1699 (.A(_04146_),
    .X(net4296));
 sg13g2_dlygate4sd3_1 hold1700 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[13] ),
    .X(net4297));
 sg13g2_dlygate4sd3_1 hold1701 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.bit_idx[4] ),
    .X(net4298));
 sg13g2_dlygate4sd3_1 hold1702 (.A(_01333_),
    .X(net4299));
 sg13g2_dlygate4sd3_1 hold1703 (.A(\soc_I.kianv_I.Instr[0] ),
    .X(net4300));
 sg13g2_dlygate4sd3_1 hold1704 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[61] ),
    .X(net4301));
 sg13g2_dlygate4sd3_1 hold1705 (.A(_05623_),
    .X(net4302));
 sg13g2_dlygate4sd3_1 hold1706 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[16] ),
    .X(net4303));
 sg13g2_dlygate4sd3_1 hold1707 (.A(\soc_I.clint_I.mtime[60] ),
    .X(net4304));
 sg13g2_dlygate4sd3_1 hold1708 (.A(_06436_),
    .X(net4305));
 sg13g2_dlygate4sd3_1 hold1709 (.A(_01692_),
    .X(net4306));
 sg13g2_dlygate4sd3_1 hold1710 (.A(\soc_I.spi0_I.sclk ),
    .X(net4307));
 sg13g2_dlygate4sd3_1 hold1711 (.A(_06565_),
    .X(net4308));
 sg13g2_dlygate4sd3_1 hold1712 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[29] ),
    .X(net4309));
 sg13g2_dlygate4sd3_1 hold1713 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[1] ),
    .X(net4310));
 sg13g2_dlygate4sd3_1 hold1714 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[28] ),
    .X(net4311));
 sg13g2_dlygate4sd3_1 hold1715 (.A(\soc_I.spi_div_reg[29] ),
    .X(net4312));
 sg13g2_dlygate4sd3_1 hold1716 (.A(_00289_),
    .X(net4313));
 sg13g2_dlygate4sd3_1 hold1717 (.A(_06823_),
    .X(net4314));
 sg13g2_dlygate4sd3_1 hold1718 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[15] ),
    .X(net4315));
 sg13g2_dlygate4sd3_1 hold1719 (.A(\soc_I.spi0_I.spi_buf[3] ),
    .X(net4316));
 sg13g2_dlygate4sd3_1 hold1720 (.A(_01974_),
    .X(net4317));
 sg13g2_dlygate4sd3_1 hold1721 (.A(\soc_I.rx_uart_i.fifo_i.ram[6][7] ),
    .X(net4318));
 sg13g2_dlygate4sd3_1 hold1722 (.A(_02294_),
    .X(net4319));
 sg13g2_dlygate4sd3_1 hold1723 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[5] ),
    .X(net4320));
 sg13g2_dlygate4sd3_1 hold1724 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[2] ),
    .X(net4321));
 sg13g2_dlygate4sd3_1 hold1725 (.A(_04432_),
    .X(net4322));
 sg13g2_dlygate4sd3_1 hold1726 (.A(_01005_),
    .X(net4323));
 sg13g2_dlygate4sd3_1 hold1727 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[8] ),
    .X(net4324));
 sg13g2_dlygate4sd3_1 hold1728 (.A(_08485_),
    .X(net4325));
 sg13g2_dlygate4sd3_1 hold1729 (.A(\soc_I.clint_I.tick_cnt[8] ),
    .X(net4326));
 sg13g2_dlygate4sd3_1 hold1730 (.A(_06237_),
    .X(net4327));
 sg13g2_dlygate4sd3_1 hold1731 (.A(\soc_I.rx_uart_i.fifo_i.ram[0][1] ),
    .X(net4328));
 sg13g2_dlygate4sd3_1 hold1732 (.A(_00631_),
    .X(net4329));
 sg13g2_dlygate4sd3_1 hold1733 (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[11] ),
    .X(net4330));
 sg13g2_dlygate4sd3_1 hold1734 (.A(_01450_),
    .X(net4331));
 sg13g2_dlygate4sd3_1 hold1735 (.A(\soc_I.clint_I.mtime[9] ),
    .X(net4332));
 sg13g2_dlygate4sd3_1 hold1736 (.A(_01641_),
    .X(net4333));
 sg13g2_dlygate4sd3_1 hold1737 (.A(\soc_I.clint_I.tick_cnt[17] ),
    .X(net4334));
 sg13g2_dlygate4sd3_1 hold1738 (.A(_06253_),
    .X(net4335));
 sg13g2_dlygate4sd3_1 hold1739 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[4] ),
    .X(net4336));
 sg13g2_dlygate4sd3_1 hold1740 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[20] ),
    .X(net4337));
 sg13g2_dlygate4sd3_1 hold1741 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[14] ),
    .X(net4338));
 sg13g2_dlygate4sd3_1 hold1742 (.A(_04490_),
    .X(net4339));
 sg13g2_dlygate4sd3_1 hold1743 (.A(_01017_),
    .X(net4340));
 sg13g2_dlygate4sd3_1 hold1744 (.A(\soc_I.spi_div_reg[17] ),
    .X(net4341));
 sg13g2_dlygate4sd3_1 hold1745 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[26][18] ),
    .X(net4342));
 sg13g2_dlygate4sd3_1 hold1746 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[36] ),
    .X(net4343));
 sg13g2_dlygate4sd3_1 hold1747 (.A(_05581_),
    .X(net4344));
 sg13g2_dlygate4sd3_1 hold1748 (.A(_01301_),
    .X(net4345));
 sg13g2_dlygate4sd3_1 hold1749 (.A(\soc_I.spi0_I.tick_cnt[13] ),
    .X(net4346));
 sg13g2_dlygate4sd3_1 hold1750 (.A(_06635_),
    .X(net4347));
 sg13g2_dlygate4sd3_1 hold1751 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[21] ),
    .X(net4348));
 sg13g2_dlygate4sd3_1 hold1752 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[15] ),
    .X(net4349));
 sg13g2_dlygate4sd3_1 hold1753 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[0] ),
    .X(net4350));
 sg13g2_dlygate4sd3_1 hold1754 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[14] ),
    .X(net4351));
 sg13g2_dlygate4sd3_1 hold1755 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[31][19] ),
    .X(net4352));
 sg13g2_dlygate4sd3_1 hold1756 (.A(\soc_I.PC[29] ),
    .X(net4353));
 sg13g2_dlygate4sd3_1 hold1757 (.A(_01468_),
    .X(net4354));
 sg13g2_dlygate4sd3_1 hold1758 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[29] ),
    .X(net4355));
 sg13g2_dlygate4sd3_1 hold1759 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[13] ),
    .X(net4356));
 sg13g2_dlygate4sd3_1 hold1760 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[17] ),
    .X(net4357));
 sg13g2_dlygate4sd3_1 hold1761 (.A(_00857_),
    .X(net4358));
 sg13g2_dlygate4sd3_1 hold1762 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[4] ),
    .X(net4359));
 sg13g2_dlygate4sd3_1 hold1763 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[19] ),
    .X(net4360));
 sg13g2_dlygate4sd3_1 hold1764 (.A(\soc_I.spi_div_reg[31] ),
    .X(net4361));
 sg13g2_dlygate4sd3_1 hold1765 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[1] ),
    .X(net4362));
 sg13g2_dlygate4sd3_1 hold1766 (.A(_05316_),
    .X(net4363));
 sg13g2_dlygate4sd3_1 hold1767 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[19] ),
    .X(net4364));
 sg13g2_dlygate4sd3_1 hold1768 (.A(_05553_),
    .X(net4365));
 sg13g2_dlygate4sd3_1 hold1769 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[18] ),
    .X(net4366));
 sg13g2_dlygate4sd3_1 hold1770 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[49] ),
    .X(net4367));
 sg13g2_dlygate4sd3_1 hold1771 (.A(_02159_),
    .X(net4368));
 sg13g2_dlygate4sd3_1 hold1772 (.A(\soc_I.spi_div_reg[21] ),
    .X(net4369));
 sg13g2_dlygate4sd3_1 hold1773 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[19] ),
    .X(net4370));
 sg13g2_dlygate4sd3_1 hold1774 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[31] ),
    .X(net4371));
 sg13g2_dlygate4sd3_1 hold1775 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[19] ),
    .X(net4372));
 sg13g2_dlygate4sd3_1 hold1776 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[21] ),
    .X(net4373));
 sg13g2_dlygate4sd3_1 hold1777 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[25] ),
    .X(net4374));
 sg13g2_dlygate4sd3_1 hold1778 (.A(_05563_),
    .X(net4375));
 sg13g2_dlygate4sd3_1 hold1779 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[7] ),
    .X(net4376));
 sg13g2_dlygate4sd3_1 hold1780 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[31] ),
    .X(net4377));
 sg13g2_dlygate4sd3_1 hold1781 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[23] ),
    .X(net4378));
 sg13g2_dlygate4sd3_1 hold1782 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[23] ),
    .X(net4379));
 sg13g2_dlygate4sd3_1 hold1783 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[17] ),
    .X(net4380));
 sg13g2_dlygate4sd3_1 hold1784 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[29] ),
    .X(net4381));
 sg13g2_dlygate4sd3_1 hold1785 (.A(\soc_I.qqspi_I.rdata[23] ),
    .X(net4382));
 sg13g2_dlygate4sd3_1 hold1786 (.A(_01819_),
    .X(net4383));
 sg13g2_dlygate4sd3_1 hold1787 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[5] ),
    .X(net4384));
 sg13g2_dlygate4sd3_1 hold1788 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[22] ),
    .X(net4385));
 sg13g2_dlygate4sd3_1 hold1789 (.A(\soc_I.clint_I.mtimecmp[41] ),
    .X(net4386));
 sg13g2_dlygate4sd3_1 hold1790 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[15] ),
    .X(net4387));
 sg13g2_dlygate4sd3_1 hold1791 (.A(_04688_),
    .X(net4388));
 sg13g2_dlygate4sd3_1 hold1792 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[49] ),
    .X(net4389));
 sg13g2_dlygate4sd3_1 hold1793 (.A(_05603_),
    .X(net4390));
 sg13g2_dlygate4sd3_1 hold1794 (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[4] ),
    .X(net4391));
 sg13g2_dlygate4sd3_1 hold1795 (.A(\soc_I.spi_div_reg[28] ),
    .X(net4392));
 sg13g2_dlygate4sd3_1 hold1796 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[7] ),
    .X(net4393));
 sg13g2_dlygate4sd3_1 hold1797 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[9] ),
    .X(net4394));
 sg13g2_dlygate4sd3_1 hold1798 (.A(\soc_I.rx_uart_i.fifo_i.ram[3][5] ),
    .X(net4395));
 sg13g2_dlygate4sd3_1 hold1799 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[8] ),
    .X(net4396));
 sg13g2_dlygate4sd3_1 hold1800 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[28] ),
    .X(net4397));
 sg13g2_dlygate4sd3_1 hold1801 (.A(_04178_),
    .X(net4398));
 sg13g2_dlygate4sd3_1 hold1802 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[18] ),
    .X(net4399));
 sg13g2_dlygate4sd3_1 hold1803 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[27] ),
    .X(net4400));
 sg13g2_dlygate4sd3_1 hold1804 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[30] ),
    .X(net4401));
 sg13g2_dlygate4sd3_1 hold1805 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[10] ),
    .X(net4402));
 sg13g2_dlygate4sd3_1 hold1806 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[22] ),
    .X(net4403));
 sg13g2_dlygate4sd3_1 hold1807 (.A(_04522_),
    .X(net4404));
 sg13g2_dlygate4sd3_1 hold1808 (.A(_01025_),
    .X(net4405));
 sg13g2_dlygate4sd3_1 hold1809 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[31] ),
    .X(net4406));
 sg13g2_dlygate4sd3_1 hold1810 (.A(_04184_),
    .X(net4407));
 sg13g2_dlygate4sd3_1 hold1811 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[23] ),
    .X(net4408));
 sg13g2_dlygate4sd3_1 hold1812 (.A(_05465_),
    .X(net4409));
 sg13g2_dlygate4sd3_1 hold1813 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[17] ),
    .X(net4410));
 sg13g2_dlygate4sd3_1 hold1814 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[2] ),
    .X(net4411));
 sg13g2_dlygate4sd3_1 hold1815 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[27] ),
    .X(net4412));
 sg13g2_dlygate4sd3_1 hold1816 (.A(\soc_I.spi0_I.tick_cnt[4] ),
    .X(net4413));
 sg13g2_dlygate4sd3_1 hold1817 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[2] ),
    .X(net4414));
 sg13g2_dlygate4sd3_1 hold1818 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[18] ),
    .X(net4415));
 sg13g2_dlygate4sd3_1 hold1819 (.A(_04506_),
    .X(net4416));
 sg13g2_dlygate4sd3_1 hold1820 (.A(_01021_),
    .X(net4417));
 sg13g2_dlygate4sd3_1 hold1821 (.A(\soc_I.clint_I.div[12] ),
    .X(net4418));
 sg13g2_dlygate4sd3_1 hold1822 (.A(\soc_I.tx_uart_i.tx_data_reg[6] ),
    .X(net4419));
 sg13g2_dlygate4sd3_1 hold1823 (.A(\soc_I.clint_I.div[4] ),
    .X(net4420));
 sg13g2_dlygate4sd3_1 hold1824 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[16] ),
    .X(net4421));
 sg13g2_dlygate4sd3_1 hold1825 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[23] ),
    .X(net4422));
 sg13g2_dlygate4sd3_1 hold1826 (.A(_04526_),
    .X(net4423));
 sg13g2_dlygate4sd3_1 hold1827 (.A(_01026_),
    .X(net4424));
 sg13g2_dlygate4sd3_1 hold1828 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[30][11] ),
    .X(net4425));
 sg13g2_dlygate4sd3_1 hold1829 (.A(\soc_I.tx_uart_i.wait_states[15] ),
    .X(net4426));
 sg13g2_dlygate4sd3_1 hold1830 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[5] ),
    .X(net4427));
 sg13g2_dlygate4sd3_1 hold1831 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[30] ),
    .X(net4428));
 sg13g2_dlygate4sd3_1 hold1832 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[14] ),
    .X(net4429));
 sg13g2_dlygate4sd3_1 hold1833 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[9] ),
    .X(net4430));
 sg13g2_dlygate4sd3_1 hold1834 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[25] ),
    .X(net4431));
 sg13g2_dlygate4sd3_1 hold1835 (.A(\soc_I.clint_I.tick_cnt[3] ),
    .X(net4432));
 sg13g2_dlygate4sd3_1 hold1836 (.A(_06227_),
    .X(net4433));
 sg13g2_dlygate4sd3_1 hold1837 (.A(\soc_I.spi0_I.tick_cnt[11] ),
    .X(net4434));
 sg13g2_dlygate4sd3_1 hold1838 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[10] ),
    .X(net4435));
 sg13g2_dlygate4sd3_1 hold1839 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[0] ),
    .X(net4436));
 sg13g2_dlygate4sd3_1 hold1840 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[30] ),
    .X(net4437));
 sg13g2_dlygate4sd3_1 hold1841 (.A(\soc_I.spi_div_reg[16] ),
    .X(net4438));
 sg13g2_dlygate4sd3_1 hold1842 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[40] ),
    .X(net4439));
 sg13g2_dlygate4sd3_1 hold1843 (.A(_04751_),
    .X(net4440));
 sg13g2_dlygate4sd3_1 hold1844 (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[9] ),
    .X(net4441));
 sg13g2_dlygate4sd3_1 hold1845 (.A(\soc_I.rx_uart_i.rx_in_sync[1] ),
    .X(net4442));
 sg13g2_dlygate4sd3_1 hold1846 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[2] ),
    .X(net4443));
 sg13g2_dlygate4sd3_1 hold1847 (.A(\soc_I.spi_div_reg[25] ),
    .X(net4444));
 sg13g2_dlygate4sd3_1 hold1848 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[17] ),
    .X(net4445));
 sg13g2_dlygate4sd3_1 hold1849 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[24] ),
    .X(net4446));
 sg13g2_dlygate4sd3_1 hold1850 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[11] ),
    .X(net4447));
 sg13g2_dlygate4sd3_1 hold1851 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[0] ),
    .X(net4448));
 sg13g2_dlygate4sd3_1 hold1852 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[15] ),
    .X(net4449));
 sg13g2_dlygate4sd3_1 hold1853 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[12] ),
    .X(net4450));
 sg13g2_dlygate4sd3_1 hold1854 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[0] ),
    .X(net4451));
 sg13g2_dlygate4sd3_1 hold1855 (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[3] ),
    .X(net4452));
 sg13g2_dlygate4sd3_1 hold1856 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[15] ),
    .X(net4453));
 sg13g2_dlygate4sd3_1 hold1857 (.A(\soc_I.clint_I.div[8] ),
    .X(net4454));
 sg13g2_dlygate4sd3_1 hold1858 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[9] ),
    .X(net4455));
 sg13g2_dlygate4sd3_1 hold1859 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[27] ),
    .X(net4456));
 sg13g2_dlygate4sd3_1 hold1860 (.A(_00867_),
    .X(net4457));
 sg13g2_dlygate4sd3_1 hold1861 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[13] ),
    .X(net4458));
 sg13g2_dlygate4sd3_1 hold1862 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[16] ),
    .X(net4459));
 sg13g2_dlygate4sd3_1 hold1863 (.A(_00856_),
    .X(net4460));
 sg13g2_dlygate4sd3_1 hold1864 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[29] ),
    .X(net4461));
 sg13g2_dlygate4sd3_1 hold1865 (.A(_00869_),
    .X(net4462));
 sg13g2_dlygate4sd3_1 hold1866 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[28] ),
    .X(net4463));
 sg13g2_dlygate4sd3_1 hold1867 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[8] ),
    .X(net4464));
 sg13g2_dlygate4sd3_1 hold1868 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[22] ),
    .X(net4465));
 sg13g2_dlygate4sd3_1 hold1869 (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[13] ),
    .X(net4466));
 sg13g2_dlygate4sd3_1 hold1870 (.A(\soc_I.spi0_I.tick_cnt[12] ),
    .X(net4467));
 sg13g2_dlygate4sd3_1 hold1871 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[31] ),
    .X(net4468));
 sg13g2_dlygate4sd3_1 hold1872 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[5] ),
    .X(net4469));
 sg13g2_dlygate4sd3_1 hold1873 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[22] ),
    .X(net4470));
 sg13g2_dlygate4sd3_1 hold1874 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[24] ),
    .X(net4471));
 sg13g2_dlygate4sd3_1 hold1875 (.A(\soc_I.rx_uart_i.bit_idx[2] ),
    .X(net4472));
 sg13g2_dlygate4sd3_1 hold1876 (.A(_06831_),
    .X(net4473));
 sg13g2_dlygate4sd3_1 hold1877 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[29] ),
    .X(net4474));
 sg13g2_dlygate4sd3_1 hold1878 (.A(_04723_),
    .X(net4475));
 sg13g2_dlygate4sd3_1 hold1879 (.A(_01166_),
    .X(net4476));
 sg13g2_dlygate4sd3_1 hold1880 (.A(\soc_I.qqspi_I.xfer_cycles[1] ),
    .X(net4477));
 sg13g2_dlygate4sd3_1 hold1881 (.A(_00775_),
    .X(net4478));
 sg13g2_dlygate4sd3_1 hold1882 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[20] ),
    .X(net4479));
 sg13g2_dlygate4sd3_1 hold1883 (.A(\soc_I.rst_cnt[1] ),
    .X(net4480));
 sg13g2_dlygate4sd3_1 hold1884 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[31] ),
    .X(net4481));
 sg13g2_dlygate4sd3_1 hold1885 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[13] ),
    .X(net4482));
 sg13g2_dlygate4sd3_1 hold1886 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[13] ),
    .X(net4483));
 sg13g2_dlygate4sd3_1 hold1887 (.A(_04685_),
    .X(net4484));
 sg13g2_dlygate4sd3_1 hold1888 (.A(_01150_),
    .X(net4485));
 sg13g2_dlygate4sd3_1 hold1889 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[16] ),
    .X(net4486));
 sg13g2_dlygate4sd3_1 hold1890 (.A(\soc_I.spi0_I.tick_cnt[17] ),
    .X(net4487));
 sg13g2_dlygate4sd3_1 hold1891 (.A(_06642_),
    .X(net4488));
 sg13g2_dlygate4sd3_1 hold1892 (.A(\soc_I.clint_I.mtime[4] ),
    .X(net4489));
 sg13g2_dlygate4sd3_1 hold1893 (.A(_01636_),
    .X(net4490));
 sg13g2_dlygate4sd3_1 hold1894 (.A(_00253_),
    .X(net4491));
 sg13g2_dlygate4sd3_1 hold1895 (.A(_02208_),
    .X(net4492));
 sg13g2_dlygate4sd3_1 hold1896 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[18] ),
    .X(net4493));
 sg13g2_dlygate4sd3_1 hold1897 (.A(_00112_),
    .X(net4494));
 sg13g2_dlygate4sd3_1 hold1898 (.A(_06379_),
    .X(net4495));
 sg13g2_dlygate4sd3_1 hold1899 (.A(_01665_),
    .X(net4496));
 sg13g2_dlygate4sd3_1 hold1900 (.A(\soc_I.clint_I.mtime[17] ),
    .X(net4497));
 sg13g2_dlygate4sd3_1 hold1901 (.A(_01649_),
    .X(net4498));
 sg13g2_dlygate4sd3_1 hold1902 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[13] ),
    .X(net4499));
 sg13g2_dlygate4sd3_1 hold1903 (.A(_05543_),
    .X(net4500));
 sg13g2_dlygate4sd3_1 hold1904 (.A(_00093_),
    .X(net4501));
 sg13g2_dlygate4sd3_1 hold1905 (.A(_06319_),
    .X(net4502));
 sg13g2_dlygate4sd3_1 hold1906 (.A(_01645_),
    .X(net4503));
 sg13g2_dlygate4sd3_1 hold1907 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[4] ),
    .X(net4504));
 sg13g2_dlygate4sd3_1 hold1908 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[30] ),
    .X(net4505));
 sg13g2_dlygate4sd3_1 hold1909 (.A(_00870_),
    .X(net4506));
 sg13g2_dlygate4sd3_1 hold1910 (.A(\soc_I.spi_div_reg[27] ),
    .X(net4507));
 sg13g2_dlygate4sd3_1 hold1911 (.A(\soc_I.spi0_I.tick_cnt[16] ),
    .X(net4508));
 sg13g2_dlygate4sd3_1 hold1912 (.A(_06641_),
    .X(net4509));
 sg13g2_dlygate4sd3_1 hold1913 (.A(\soc_I.clint_I.mtimecmp[33] ),
    .X(net4510));
 sg13g2_dlygate4sd3_1 hold1914 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[56] ),
    .X(net4511));
 sg13g2_dlygate4sd3_1 hold1915 (.A(_01193_),
    .X(net4512));
 sg13g2_dlygate4sd3_1 hold1916 (.A(\soc_I.tx_uart_i.tx_data_reg[2] ),
    .X(net4513));
 sg13g2_dlygate4sd3_1 hold1917 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[24] ),
    .X(net4514));
 sg13g2_dlygate4sd3_1 hold1918 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[26] ),
    .X(net4515));
 sg13g2_dlygate4sd3_1 hold1919 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[18] ),
    .X(net4516));
 sg13g2_dlygate4sd3_1 hold1920 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[13] ),
    .X(net4517));
 sg13g2_dlygate4sd3_1 hold1921 (.A(\soc_I.clint_I.mtime[11] ),
    .X(net4518));
 sg13g2_dlygate4sd3_1 hold1922 (.A(_01643_),
    .X(net4519));
 sg13g2_dlygate4sd3_1 hold1923 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[5] ),
    .X(net4520));
 sg13g2_dlygate4sd3_1 hold1924 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[15] ),
    .X(net4521));
 sg13g2_dlygate4sd3_1 hold1925 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[1] ),
    .X(net4522));
 sg13g2_dlygate4sd3_1 hold1926 (.A(\soc_I.spi_div_reg[18] ),
    .X(net4523));
 sg13g2_dlygate4sd3_1 hold1927 (.A(_00249_),
    .X(net4524));
 sg13g2_dlygate4sd3_1 hold1928 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[23] ),
    .X(net4525));
 sg13g2_dlygate4sd3_1 hold1929 (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[7] ),
    .X(net4526));
 sg13g2_dlygate4sd3_1 hold1930 (.A(_01446_),
    .X(net4527));
 sg13g2_dlygate4sd3_1 hold1931 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[27] ),
    .X(net4528));
 sg13g2_dlygate4sd3_1 hold1932 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[7] ),
    .X(net4529));
 sg13g2_dlygate4sd3_1 hold1933 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[6] ),
    .X(net4530));
 sg13g2_dlygate4sd3_1 hold1934 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[56] ),
    .X(net4531));
 sg13g2_dlygate4sd3_1 hold1935 (.A(_02152_),
    .X(net4532));
 sg13g2_dlygate4sd3_1 hold1936 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[18] ),
    .X(net4533));
 sg13g2_dlygate4sd3_1 hold1937 (.A(\soc_I.rx_uart_i.wait_states[2] ),
    .X(net4534));
 sg13g2_dlygate4sd3_1 hold1938 (.A(_01844_),
    .X(net4535));
 sg13g2_dlygate4sd3_1 hold1939 (.A(\soc_I.tx_uart_i.tx_data_reg[3] ),
    .X(net4536));
 sg13g2_dlygate4sd3_1 hold1940 (.A(\soc_I.spi0_I.ready_xfer ),
    .X(net4537));
 sg13g2_dlygate4sd3_1 hold1941 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[20] ),
    .X(net4538));
 sg13g2_dlygate4sd3_1 hold1942 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[11] ),
    .X(net4539));
 sg13g2_dlygate4sd3_1 hold1943 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[2] ),
    .X(net4540));
 sg13g2_dlygate4sd3_1 hold1944 (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[1] ),
    .X(net4541));
 sg13g2_dlygate4sd3_1 hold1945 (.A(_01440_),
    .X(net4542));
 sg13g2_dlygate4sd3_1 hold1946 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[2] ),
    .X(net4543));
 sg13g2_dlygate4sd3_1 hold1947 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[31] ),
    .X(net4544));
 sg13g2_dlygate4sd3_1 hold1948 (.A(\soc_I.rx_uart_i.bit_idx[1] ),
    .X(net4545));
 sg13g2_dlygate4sd3_1 hold1949 (.A(_06811_),
    .X(net4546));
 sg13g2_dlygate4sd3_1 hold1950 (.A(\soc_I.rx_uart_i.fifo_i.ram[5][3] ),
    .X(net4547));
 sg13g2_dlygate4sd3_1 hold1951 (.A(_02298_),
    .X(net4548));
 sg13g2_dlygate4sd3_1 hold1952 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[17] ),
    .X(net4549));
 sg13g2_dlygate4sd3_1 hold1953 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[19] ),
    .X(net4550));
 sg13g2_dlygate4sd3_1 hold1954 (.A(_04510_),
    .X(net4551));
 sg13g2_dlygate4sd3_1 hold1955 (.A(_01022_),
    .X(net4552));
 sg13g2_dlygate4sd3_1 hold1956 (.A(\soc_I.clint_I.mtimecmp[40] ),
    .X(net4553));
 sg13g2_dlygate4sd3_1 hold1957 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[6] ),
    .X(net4554));
 sg13g2_dlygate4sd3_1 hold1958 (.A(\soc_I.clint_I.mtime[29] ),
    .X(net4555));
 sg13g2_dlygate4sd3_1 hold1959 (.A(_01661_),
    .X(net4556));
 sg13g2_dlygate4sd3_1 hold1960 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[29] ),
    .X(net4557));
 sg13g2_dlygate4sd3_1 hold1961 (.A(\soc_I.tx_uart_i.tx_data_reg[5] ),
    .X(net4558));
 sg13g2_dlygate4sd3_1 hold1962 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.privilege_mode[0] ),
    .X(net4559));
 sg13g2_dlygate4sd3_1 hold1963 (.A(_01071_),
    .X(net4560));
 sg13g2_dlygate4sd3_1 hold1964 (.A(\soc_I.spi0_I.cen ),
    .X(net4561));
 sg13g2_dlygate4sd3_1 hold1965 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[5] ),
    .X(net4562));
 sg13g2_dlygate4sd3_1 hold1966 (.A(\soc_I.spi_div_reg[19] ),
    .X(net4563));
 sg13g2_dlygate4sd3_1 hold1967 (.A(\soc_I.clint_I.mtime[62] ),
    .X(net4564));
 sg13g2_dlygate4sd3_1 hold1968 (.A(_01694_),
    .X(net4565));
 sg13g2_dlygate4sd3_1 hold1969 (.A(\soc_I.PC[1] ),
    .X(net4566));
 sg13g2_dlygate4sd3_1 hold1970 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[3] ),
    .X(net4567));
 sg13g2_dlygate4sd3_1 hold1971 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[6] ),
    .X(net4568));
 sg13g2_dlygate4sd3_1 hold1972 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[21] ),
    .X(net4569));
 sg13g2_dlygate4sd3_1 hold1973 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[18] ),
    .X(net4570));
 sg13g2_dlygate4sd3_1 hold1974 (.A(\soc_I.spi0_I.tick_cnt[8] ),
    .X(net4571));
 sg13g2_dlygate4sd3_1 hold1975 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[28] ),
    .X(net4572));
 sg13g2_dlygate4sd3_1 hold1976 (.A(_00868_),
    .X(net4573));
 sg13g2_dlygate4sd3_1 hold1977 (.A(\soc_I.qqspi_I.state[6] ),
    .X(net4574));
 sg13g2_dlygate4sd3_1 hold1978 (.A(_12572_),
    .X(net4575));
 sg13g2_dlygate4sd3_1 hold1979 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[28] ),
    .X(net4576));
 sg13g2_dlygate4sd3_1 hold1980 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[24] ),
    .X(net4577));
 sg13g2_dlygate4sd3_1 hold1981 (.A(_00864_),
    .X(net4578));
 sg13g2_dlygate4sd3_1 hold1982 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[30] ),
    .X(net4579));
 sg13g2_dlygate4sd3_1 hold1983 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[9] ),
    .X(net4580));
 sg13g2_dlygate4sd3_1 hold1984 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[19] ),
    .X(net4581));
 sg13g2_dlygate4sd3_1 hold1985 (.A(\soc_I.clint_I.mtime[31] ),
    .X(net4582));
 sg13g2_dlygate4sd3_1 hold1986 (.A(_01663_),
    .X(net4583));
 sg13g2_dlygate4sd3_1 hold1987 (.A(sio0_si_mosi_o),
    .X(net4584));
 sg13g2_dlygate4sd3_1 hold1988 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[14] ),
    .X(net4585));
 sg13g2_dlygate4sd3_1 hold1989 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[12] ),
    .X(net4586));
 sg13g2_dlygate4sd3_1 hold1990 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[13][7] ),
    .X(net4587));
 sg13g2_dlygate4sd3_1 hold1991 (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[23] ),
    .X(net4588));
 sg13g2_dlygate4sd3_1 hold1992 (.A(_01462_),
    .X(net4589));
 sg13g2_dlygate4sd3_1 hold1993 (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[2] ),
    .X(net4590));
 sg13g2_dlygate4sd3_1 hold1994 (.A(_01441_),
    .X(net4591));
 sg13g2_dlygate4sd3_1 hold1995 (.A(\soc_I.clint_I.mtimecmp[0] ),
    .X(net4592));
 sg13g2_dlygate4sd3_1 hold1996 (.A(\soc_I.spi_div_reg[24] ),
    .X(net4593));
 sg13g2_dlygate4sd3_1 hold1997 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[57] ),
    .X(net4594));
 sg13g2_dlygate4sd3_1 hold1998 (.A(_05617_),
    .X(net4595));
 sg13g2_dlygate4sd3_1 hold1999 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[28] ),
    .X(net4596));
 sg13g2_dlygate4sd3_1 hold2000 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[0] ),
    .X(net4597));
 sg13g2_dlygate4sd3_1 hold2001 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[11] ),
    .X(net4598));
 sg13g2_dlygate4sd3_1 hold2002 (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[3] ),
    .X(net4599));
 sg13g2_dlygate4sd3_1 hold2003 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[25] ),
    .X(net4600));
 sg13g2_dlygate4sd3_1 hold2004 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[26] ),
    .X(net4601));
 sg13g2_dlygate4sd3_1 hold2005 (.A(\soc_I.clint_I.mtime[15] ),
    .X(net4602));
 sg13g2_dlygate4sd3_1 hold2006 (.A(_01647_),
    .X(net4603));
 sg13g2_dlygate4sd3_1 hold2007 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[23] ),
    .X(net4604));
 sg13g2_dlygate4sd3_1 hold2008 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[13] ),
    .X(net4605));
 sg13g2_dlygate4sd3_1 hold2009 (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[29] ),
    .X(net4606));
 sg13g2_dlygate4sd3_1 hold2010 (.A(\soc_I.clint_I.tick_cnt[6] ),
    .X(net4607));
 sg13g2_dlygate4sd3_1 hold2011 (.A(_06233_),
    .X(net4608));
 sg13g2_dlygate4sd3_1 hold2012 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[10] ),
    .X(net4609));
 sg13g2_dlygate4sd3_1 hold2013 (.A(_00252_),
    .X(net4610));
 sg13g2_dlygate4sd3_1 hold2014 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[16] ),
    .X(net4611));
 sg13g2_dlygate4sd3_1 hold2015 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[9] ),
    .X(net4612));
 sg13g2_dlygate4sd3_1 hold2016 (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[27] ),
    .X(net4613));
 sg13g2_dlygate4sd3_1 hold2017 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[24] ),
    .X(net4614));
 sg13g2_dlygate4sd3_1 hold2018 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[62] ),
    .X(net4615));
 sg13g2_dlygate4sd3_1 hold2019 (.A(_02146_),
    .X(net4616));
 sg13g2_dlygate4sd3_1 hold2020 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[4] ),
    .X(net4617));
 sg13g2_dlygate4sd3_1 hold2021 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[27] ),
    .X(net4618));
 sg13g2_dlygate4sd3_1 hold2022 (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[2] ),
    .X(net4619));
 sg13g2_dlygate4sd3_1 hold2023 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[7] ),
    .X(net4620));
 sg13g2_dlygate4sd3_1 hold2024 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[9] ),
    .X(net4621));
 sg13g2_dlygate4sd3_1 hold2025 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[12] ),
    .X(net4622));
 sg13g2_dlygate4sd3_1 hold2026 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[14] ),
    .X(net4623));
 sg13g2_dlygate4sd3_1 hold2027 (.A(_00854_),
    .X(net4624));
 sg13g2_dlygate4sd3_1 hold2028 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[14] ),
    .X(net4625));
 sg13g2_dlygate4sd3_1 hold2029 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[20] ),
    .X(net4626));
 sg13g2_dlygate4sd3_1 hold2030 (.A(\soc_I.spi0_I.rx_data[6] ),
    .X(net4627));
 sg13g2_dlygate4sd3_1 hold2031 (.A(_01977_),
    .X(net4628));
 sg13g2_dlygate4sd3_1 hold2032 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[25] ),
    .X(net4629));
 sg13g2_dlygate4sd3_1 hold2033 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[8] ),
    .X(net4630));
 sg13g2_dlygate4sd3_1 hold2034 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[22] ),
    .X(net4631));
 sg13g2_dlygate4sd3_1 hold2035 (.A(\soc_I.spi_div_reg[23] ),
    .X(net4632));
 sg13g2_dlygate4sd3_1 hold2036 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[16] ),
    .X(net4633));
 sg13g2_dlygate4sd3_1 hold2037 (.A(\soc_I.gpio0_I.rdata[3] ),
    .X(net4634));
 sg13g2_dlygate4sd3_1 hold2038 (.A(_01790_),
    .X(net4635));
 sg13g2_dlygate4sd3_1 hold2039 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[53] ),
    .X(net4636));
 sg13g2_dlygate4sd3_1 hold2040 (.A(_05610_),
    .X(net4637));
 sg13g2_dlygate4sd3_1 hold2041 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[6] ),
    .X(net4638));
 sg13g2_dlygate4sd3_1 hold2042 (.A(\soc_I.spi_div_reg[22] ),
    .X(net4639));
 sg13g2_dlygate4sd3_1 hold2043 (.A(\soc_I.gpio0_I.rdata[2] ),
    .X(net4640));
 sg13g2_dlygate4sd3_1 hold2044 (.A(_01789_),
    .X(net4641));
 sg13g2_dlygate4sd3_1 hold2045 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[1] ),
    .X(net4642));
 sg13g2_dlygate4sd3_1 hold2046 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[20] ),
    .X(net4643));
 sg13g2_dlygate4sd3_1 hold2047 (.A(_04162_),
    .X(net4644));
 sg13g2_dlygate4sd3_1 hold2048 (.A(\soc_I.spi0_I.spi_buf[6] ),
    .X(net4645));
 sg13g2_dlygate4sd3_1 hold2049 (.A(\soc_I.tx_uart_i.tx_data_reg[0] ),
    .X(net4646));
 sg13g2_dlygate4sd3_1 hold2050 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[54] ),
    .X(net4647));
 sg13g2_dlygate4sd3_1 hold2051 (.A(_04785_),
    .X(net4648));
 sg13g2_dlygate4sd3_1 hold2052 (.A(_01191_),
    .X(net4649));
 sg13g2_dlygate4sd3_1 hold2053 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[31] ),
    .X(net4650));
 sg13g2_dlygate4sd3_1 hold2054 (.A(_00871_),
    .X(net4651));
 sg13g2_dlygate4sd3_1 hold2055 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[25] ),
    .X(net4652));
 sg13g2_dlygate4sd3_1 hold2056 (.A(_00865_),
    .X(net4653));
 sg13g2_dlygate4sd3_1 hold2057 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[26] ),
    .X(net4654));
 sg13g2_dlygate4sd3_1 hold2058 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[3] ),
    .X(net4655));
 sg13g2_dlygate4sd3_1 hold2059 (.A(\soc_I.spi0_I.tick_cnt[15] ),
    .X(net4656));
 sg13g2_dlygate4sd3_1 hold2060 (.A(\soc_I.tx_uart_i.tx_data_reg[7] ),
    .X(net4657));
 sg13g2_dlygate4sd3_1 hold2061 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[55] ),
    .X(net4658));
 sg13g2_dlygate4sd3_1 hold2062 (.A(_08226_),
    .X(net4659));
 sg13g2_dlygate4sd3_1 hold2063 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[3] ),
    .X(net4660));
 sg13g2_dlygate4sd3_1 hold2064 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[21] ),
    .X(net4661));
 sg13g2_dlygate4sd3_1 hold2065 (.A(\soc_I.clint_I.mtimecmp[3] ),
    .X(net4662));
 sg13g2_dlygate4sd3_1 hold2066 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[23] ),
    .X(net4663));
 sg13g2_dlygate4sd3_1 hold2067 (.A(\soc_I.PC[14] ),
    .X(net4664));
 sg13g2_dlygate4sd3_1 hold2068 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[12] ),
    .X(net4665));
 sg13g2_dlygate4sd3_1 hold2069 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[48] ),
    .X(net4666));
 sg13g2_dlygate4sd3_1 hold2070 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[2] ),
    .X(net4667));
 sg13g2_dlygate4sd3_1 hold2071 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[31] ),
    .X(net4668));
 sg13g2_dlygate4sd3_1 hold2072 (.A(_05520_),
    .X(net4669));
 sg13g2_dlygate4sd3_1 hold2073 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[8] ),
    .X(net4670));
 sg13g2_dlygate4sd3_1 hold2074 (.A(_04138_),
    .X(net4671));
 sg13g2_dlygate4sd3_1 hold2075 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[29] ),
    .X(net4672));
 sg13g2_dlygate4sd3_1 hold2076 (.A(\soc_I.qqspi_I.state[3] ),
    .X(net4673));
 sg13g2_dlygate4sd3_1 hold2077 (.A(_12568_),
    .X(net4674));
 sg13g2_dlygate4sd3_1 hold2078 (.A(\soc_I.spi0_I.xfer_cycles[2] ),
    .X(net4675));
 sg13g2_dlygate4sd3_1 hold2079 (.A(_06571_),
    .X(net4676));
 sg13g2_dlygate4sd3_1 hold2080 (.A(_01748_),
    .X(net4677));
 sg13g2_dlygate4sd3_1 hold2081 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[20] ),
    .X(net4678));
 sg13g2_dlygate4sd3_1 hold2082 (.A(_00860_),
    .X(net4679));
 sg13g2_dlygate4sd3_1 hold2083 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[10] ),
    .X(net4680));
 sg13g2_dlygate4sd3_1 hold2084 (.A(\soc_I.rx_uart_i.fifo_i.din[6] ),
    .X(net4681));
 sg13g2_dlygate4sd3_1 hold2085 (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[31] ),
    .X(net4682));
 sg13g2_dlygate4sd3_1 hold2086 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[21] ),
    .X(net4683));
 sg13g2_dlygate4sd3_1 hold2087 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[0] ),
    .X(net4684));
 sg13g2_dlygate4sd3_1 hold2088 (.A(\soc_I.clint_I.tick_cnt[11] ),
    .X(net4685));
 sg13g2_dlygate4sd3_1 hold2089 (.A(_06242_),
    .X(net4686));
 sg13g2_dlygate4sd3_1 hold2090 (.A(\soc_I.clint_I.mtimecmp[5] ),
    .X(net4687));
 sg13g2_dlygate4sd3_1 hold2091 (.A(\soc_I.spi_div_reg[30] ),
    .X(net4688));
 sg13g2_dlygate4sd3_1 hold2092 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[14] ),
    .X(net4689));
 sg13g2_dlygate4sd3_1 hold2093 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[28] ),
    .X(net4690));
 sg13g2_dlygate4sd3_1 hold2094 (.A(_01031_),
    .X(net4691));
 sg13g2_dlygate4sd3_1 hold2095 (.A(\soc_I.clint_I.mtimecmp[49] ),
    .X(net4692));
 sg13g2_dlygate4sd3_1 hold2096 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[10] ),
    .X(net4693));
 sg13g2_dlygate4sd3_1 hold2097 (.A(\soc_I.clint_I.mtimecmp[56] ),
    .X(net4694));
 sg13g2_dlygate4sd3_1 hold2098 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[5] ),
    .X(net4695));
 sg13g2_dlygate4sd3_1 hold2099 (.A(_00909_),
    .X(net4696));
 sg13g2_dlygate4sd3_1 hold2100 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[12] ),
    .X(net4697));
 sg13g2_dlygate4sd3_1 hold2101 (.A(_04684_),
    .X(net4698));
 sg13g2_dlygate4sd3_1 hold2102 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[6] ),
    .X(net4699));
 sg13g2_dlygate4sd3_1 hold2103 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[8] ),
    .X(net4700));
 sg13g2_dlygate4sd3_1 hold2104 (.A(\soc_I.spi_div_reg[20] ),
    .X(net4701));
 sg13g2_dlygate4sd3_1 hold2105 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[14] ),
    .X(net4702));
 sg13g2_dlygate4sd3_1 hold2106 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[26] ),
    .X(net4703));
 sg13g2_dlygate4sd3_1 hold2107 (.A(\soc_I.qqspi_I.xfer_cycles[0] ),
    .X(net4704));
 sg13g2_dlygate4sd3_1 hold2108 (.A(_00774_),
    .X(net4705));
 sg13g2_dlygate4sd3_1 hold2109 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[11] ),
    .X(net4706));
 sg13g2_dlygate4sd3_1 hold2110 (.A(\soc_I.clint_I.mtimecmp[46] ),
    .X(net4707));
 sg13g2_dlygate4sd3_1 hold2111 (.A(\soc_I.clint_I.mtimecmp[37] ),
    .X(net4708));
 sg13g2_dlygate4sd3_1 hold2112 (.A(\gpio_uo_out[6] ),
    .X(net4709));
 sg13g2_dlygate4sd3_1 hold2113 (.A(\soc_I.clint_I.mtimecmp[48] ),
    .X(net4710));
 sg13g2_dlygate4sd3_1 hold2114 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[30] ),
    .X(net4711));
 sg13g2_dlygate4sd3_1 hold2115 (.A(_04182_),
    .X(net4712));
 sg13g2_dlygate4sd3_1 hold2116 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[4] ),
    .X(net4713));
 sg13g2_dlygate4sd3_1 hold2117 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[27] ),
    .X(net4714));
 sg13g2_dlygate4sd3_1 hold2118 (.A(_05567_),
    .X(net4715));
 sg13g2_dlygate4sd3_1 hold2119 (.A(\soc_I.tx_uart_i.wait_states[6] ),
    .X(net4716));
 sg13g2_dlygate4sd3_1 hold2120 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[8] ),
    .X(net4717));
 sg13g2_dlygate4sd3_1 hold2121 (.A(_05536_),
    .X(net4718));
 sg13g2_dlygate4sd3_1 hold2122 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[0] ),
    .X(net4719));
 sg13g2_dlygate4sd3_1 hold2123 (.A(\soc_I.clint_I.mtimecmp[39] ),
    .X(net4720));
 sg13g2_dlygate4sd3_1 hold2124 (.A(\soc_I.clint_I.mtime[52] ),
    .X(net4721));
 sg13g2_dlygate4sd3_1 hold2125 (.A(_06420_),
    .X(net4722));
 sg13g2_dlygate4sd3_1 hold2126 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[37] ),
    .X(net4723));
 sg13g2_dlygate4sd3_1 hold2127 (.A(_05583_),
    .X(net4724));
 sg13g2_dlygate4sd3_1 hold2128 (.A(_00060_),
    .X(net4725));
 sg13g2_dlygate4sd3_1 hold2129 (.A(_01655_),
    .X(net4726));
 sg13g2_dlygate4sd3_1 hold2130 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[21] ),
    .X(net4727));
 sg13g2_dlygate4sd3_1 hold2131 (.A(_00861_),
    .X(net4728));
 sg13g2_dlygate4sd3_1 hold2132 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[14] ),
    .X(net4729));
 sg13g2_dlygate4sd3_1 hold2133 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[26] ),
    .X(net4730));
 sg13g2_dlygate4sd3_1 hold2134 (.A(_00866_),
    .X(net4731));
 sg13g2_dlygate4sd3_1 hold2135 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[6] ),
    .X(net4732));
 sg13g2_dlygate4sd3_1 hold2136 (.A(_00910_),
    .X(net4733));
 sg13g2_dlygate4sd3_1 hold2137 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[9] ),
    .X(net4734));
 sg13g2_dlygate4sd3_1 hold2138 (.A(\soc_I.tx_uart_i.bit_idx[1] ),
    .X(net4735));
 sg13g2_dlygate4sd3_1 hold2139 (.A(_06987_),
    .X(net4736));
 sg13g2_dlygate4sd3_1 hold2140 (.A(\soc_I.clint_I.mtimecmp[27] ),
    .X(net4737));
 sg13g2_dlygate4sd3_1 hold2141 (.A(\soc_I.spi0_I.xfer_cycles[5] ),
    .X(net4738));
 sg13g2_dlygate4sd3_1 hold2142 (.A(_06580_),
    .X(net4739));
 sg13g2_dlygate4sd3_1 hold2143 (.A(_01751_),
    .X(net4740));
 sg13g2_dlygate4sd3_1 hold2144 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[22] ),
    .X(net4741));
 sg13g2_dlygate4sd3_1 hold2145 (.A(_00862_),
    .X(net4742));
 sg13g2_dlygate4sd3_1 hold2146 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[0] ),
    .X(net4743));
 sg13g2_dlygate4sd3_1 hold2147 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[12] ),
    .X(net4744));
 sg13g2_dlygate4sd3_1 hold2148 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[12] ),
    .X(net4745));
 sg13g2_dlygate4sd3_1 hold2149 (.A(_04604_),
    .X(net4746));
 sg13g2_dlygate4sd3_1 hold2150 (.A(\gpio_uo_out[2] ),
    .X(net4747));
 sg13g2_dlygate4sd3_1 hold2151 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[29] ),
    .X(net4748));
 sg13g2_dlygate4sd3_1 hold2152 (.A(\soc_I.clint_I.mtimecmp[51] ),
    .X(net4749));
 sg13g2_dlygate4sd3_1 hold2153 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[16] ),
    .X(net4750));
 sg13g2_dlygate4sd3_1 hold2154 (.A(\soc_I.clint_I.mtimecmp[4] ),
    .X(net4751));
 sg13g2_dlygate4sd3_1 hold2155 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[19] ),
    .X(net4752));
 sg13g2_dlygate4sd3_1 hold2156 (.A(\soc_I.tx_uart_i.bit_idx[2] ),
    .X(net4753));
 sg13g2_dlygate4sd3_1 hold2157 (.A(\soc_I.clint_I.mtimecmp[7] ),
    .X(net4754));
 sg13g2_dlygate4sd3_1 hold2158 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[39] ),
    .X(net4755));
 sg13g2_dlygate4sd3_1 hold2159 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[21] ),
    .X(net4756));
 sg13g2_dlygate4sd3_1 hold2160 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[11] ),
    .X(net4757));
 sg13g2_dlygate4sd3_1 hold2161 (.A(\soc_I.clint_I.mtimecmp[42] ),
    .X(net4758));
 sg13g2_dlygate4sd3_1 hold2162 (.A(\soc_I.rx_uart_i.wait_states[10] ),
    .X(net4759));
 sg13g2_dlygate4sd3_1 hold2163 (.A(_01852_),
    .X(net4760));
 sg13g2_dlygate4sd3_1 hold2164 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[15] ),
    .X(net4761));
 sg13g2_dlygate4sd3_1 hold2165 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[2] ),
    .X(net4762));
 sg13g2_dlygate4sd3_1 hold2166 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[56] ),
    .X(net4763));
 sg13g2_dlygate4sd3_1 hold2167 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[23] ),
    .X(net4764));
 sg13g2_dlygate4sd3_1 hold2168 (.A(\soc_I.clint_I.mtime[30] ),
    .X(net4765));
 sg13g2_dlygate4sd3_1 hold2169 (.A(_06373_),
    .X(net4766));
 sg13g2_dlygate4sd3_1 hold2170 (.A(\soc_I.spi0_I.div[8] ),
    .X(net4767));
 sg13g2_dlygate4sd3_1 hold2171 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[25] ),
    .X(net4768));
 sg13g2_dlygate4sd3_1 hold2172 (.A(_05479_),
    .X(net4769));
 sg13g2_dlygate4sd3_1 hold2173 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[2] ),
    .X(net4770));
 sg13g2_dlygate4sd3_1 hold2174 (.A(_00286_),
    .X(net4771));
 sg13g2_dlygate4sd3_1 hold2175 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[54] ),
    .X(net4772));
 sg13g2_dlygate4sd3_1 hold2176 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[6] ),
    .X(net4773));
 sg13g2_dlygate4sd3_1 hold2177 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mcause[31] ),
    .X(net4774));
 sg13g2_dlygate4sd3_1 hold2178 (.A(\soc_I.clint_I.mtimecmp[6] ),
    .X(net4775));
 sg13g2_dlygate4sd3_1 hold2179 (.A(\soc_I.clint_I.mtime[63] ),
    .X(net4776));
 sg13g2_dlygate4sd3_1 hold2180 (.A(_01695_),
    .X(net4777));
 sg13g2_dlygate4sd3_1 hold2181 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[24] ),
    .X(net4778));
 sg13g2_dlygate4sd3_1 hold2182 (.A(_04170_),
    .X(net4779));
 sg13g2_dlygate4sd3_1 hold2183 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[9] ),
    .X(net4780));
 sg13g2_dlygate4sd3_1 hold2184 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[1] ),
    .X(net4781));
 sg13g2_dlygate4sd3_1 hold2185 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.privilege_mode[1] ),
    .X(net4782));
 sg13g2_dlygate4sd3_1 hold2186 (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[27] ),
    .X(net4783));
 sg13g2_dlygate4sd3_1 hold2187 (.A(_01466_),
    .X(net4784));
 sg13g2_dlygate4sd3_1 hold2188 (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[21] ),
    .X(net4785));
 sg13g2_dlygate4sd3_1 hold2189 (.A(_01460_),
    .X(net4786));
 sg13g2_dlygate4sd3_1 hold2190 (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[15] ),
    .X(net4787));
 sg13g2_dlygate4sd3_1 hold2191 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[19] ),
    .X(net4788));
 sg13g2_dlygate4sd3_1 hold2192 (.A(_00859_),
    .X(net4789));
 sg13g2_dlygate4sd3_1 hold2193 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[31] ),
    .X(net4790));
 sg13g2_dlygate4sd3_1 hold2194 (.A(_01034_),
    .X(net4791));
 sg13g2_dlygate4sd3_1 hold2195 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[13] ),
    .X(net4792));
 sg13g2_dlygate4sd3_1 hold2196 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[62] ),
    .X(net4793));
 sg13g2_dlygate4sd3_1 hold2197 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[4] ),
    .X(net4794));
 sg13g2_dlygate4sd3_1 hold2198 (.A(\soc_I.kianv_I.amo_reserved_state_load ),
    .X(net4795));
 sg13g2_dlygate4sd3_1 hold2199 (.A(\gpio_uo_out[0] ),
    .X(net4796));
 sg13g2_dlygate4sd3_1 hold2200 (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[10] ),
    .X(net4797));
 sg13g2_dlygate4sd3_1 hold2201 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[13] ),
    .X(net4798));
 sg13g2_dlygate4sd3_1 hold2202 (.A(\soc_I.clint_I.mtimecmp[32] ),
    .X(net4799));
 sg13g2_dlygate4sd3_1 hold2203 (.A(\soc_I.PC[0] ),
    .X(net4800));
 sg13g2_dlygate4sd3_1 hold2204 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[27] ),
    .X(net4801));
 sg13g2_dlygate4sd3_1 hold2205 (.A(_00175_),
    .X(net4802));
 sg13g2_dlygate4sd3_1 hold2206 (.A(_05393_),
    .X(net4803));
 sg13g2_dlygate4sd3_1 hold2207 (.A(\soc_I.clint_I.mtimecmp[14] ),
    .X(net4804));
 sg13g2_dlygate4sd3_1 hold2208 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[3] ),
    .X(net4805));
 sg13g2_dlygate4sd3_1 hold2209 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[26] ),
    .X(net4806));
 sg13g2_dlygate4sd3_1 hold2210 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[61] ),
    .X(net4807));
 sg13g2_dlygate4sd3_1 hold2211 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[22] ),
    .X(net4808));
 sg13g2_dlygate4sd3_1 hold2212 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[41] ),
    .X(net4809));
 sg13g2_dlygate4sd3_1 hold2213 (.A(_05590_),
    .X(net4810));
 sg13g2_dlygate4sd3_1 hold2214 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[22] ),
    .X(net4811));
 sg13g2_dlygate4sd3_1 hold2215 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[3] ),
    .X(net4812));
 sg13g2_dlygate4sd3_1 hold2216 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[47] ),
    .X(net4813));
 sg13g2_dlygate4sd3_1 hold2217 (.A(_05600_),
    .X(net4814));
 sg13g2_dlygate4sd3_1 hold2218 (.A(\soc_I.spi_div_reg[26] ),
    .X(net4815));
 sg13g2_dlygate4sd3_1 hold2219 (.A(\soc_I.clint_I.mtimecmp[36] ),
    .X(net4816));
 sg13g2_dlygate4sd3_1 hold2220 (.A(\soc_I.qqspi_I.ready ),
    .X(net4817));
 sg13g2_dlygate4sd3_1 hold2221 (.A(_07293_),
    .X(net4818));
 sg13g2_dlygate4sd3_1 hold2222 (.A(\soc_I.clint_I.mtime[51] ),
    .X(net4819));
 sg13g2_dlygate4sd3_1 hold2223 (.A(_06418_),
    .X(net4820));
 sg13g2_dlygate4sd3_1 hold2224 (.A(_00162_),
    .X(net4821));
 sg13g2_dlygate4sd3_1 hold2225 (.A(_05486_),
    .X(net4822));
 sg13g2_dlygate4sd3_1 hold2226 (.A(\soc_I.spi0_I.xfer_cycles[5] ),
    .X(net4823));
 sg13g2_dlygate4sd3_1 hold2227 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[24] ),
    .X(net4824));
 sg13g2_dlygate4sd3_1 hold2228 (.A(\soc_I.clint_I.mtime[58] ),
    .X(net4825));
 sg13g2_dlygate4sd3_1 hold2229 (.A(_06433_),
    .X(net4826));
 sg13g2_dlygate4sd3_1 hold2230 (.A(_01691_),
    .X(net4827));
 sg13g2_dlygate4sd3_1 hold2231 (.A(\soc_I.spi0_I.spi_buf[0] ),
    .X(net4828));
 sg13g2_dlygate4sd3_1 hold2232 (.A(\soc_I.clint_I.mtimecmp[60] ),
    .X(net4829));
 sg13g2_dlygate4sd3_1 hold2233 (.A(\soc_I.clint_I.mtimecmp[29] ),
    .X(net4830));
 sg13g2_dlygate4sd3_1 hold2234 (.A(\soc_I.clint_I.mtimecmp[59] ),
    .X(net4831));
 sg13g2_dlygate4sd3_1 hold2235 (.A(\soc_I.clint_I.mtimecmp[28] ),
    .X(net4832));
 sg13g2_dlygate4sd3_1 hold2236 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[11] ),
    .X(net4833));
 sg13g2_dlygate4sd3_1 hold2237 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[50] ),
    .X(net4834));
 sg13g2_dlygate4sd3_1 hold2238 (.A(_02158_),
    .X(net4835));
 sg13g2_dlygate4sd3_1 hold2239 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[5] ),
    .X(net4836));
 sg13g2_dlygate4sd3_1 hold2240 (.A(\soc_I.clint_I.mtimecmp[17] ),
    .X(net4837));
 sg13g2_dlygate4sd3_1 hold2241 (.A(\soc_I.clint_I.tick_cnt[15] ),
    .X(net4838));
 sg13g2_dlygate4sd3_1 hold2242 (.A(_06249_),
    .X(net4839));
 sg13g2_dlygate4sd3_1 hold2243 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[22] ),
    .X(net4840));
 sg13g2_dlygate4sd3_1 hold2244 (.A(_04166_),
    .X(net4841));
 sg13g2_dlygate4sd3_1 hold2245 (.A(\soc_I.clint_I.mtimecmp[21] ),
    .X(net4842));
 sg13g2_dlygate4sd3_1 hold2246 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[32] ),
    .X(net4843));
 sg13g2_dlygate4sd3_1 hold2247 (.A(\soc_I.clint_I.tick_cnt[10] ),
    .X(net4844));
 sg13g2_dlygate4sd3_1 hold2248 (.A(_06240_),
    .X(net4845));
 sg13g2_dlygate4sd3_1 hold2249 (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[25] ),
    .X(net4846));
 sg13g2_dlygate4sd3_1 hold2250 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[4] ),
    .X(net4847));
 sg13g2_dlygate4sd3_1 hold2251 (.A(_04447_),
    .X(net4848));
 sg13g2_dlygate4sd3_1 hold2252 (.A(\soc_I.clint_I.mtimecmp[55] ),
    .X(net4849));
 sg13g2_dlygate4sd3_1 hold2253 (.A(\soc_I.rx_uart_i.wait_states[8] ),
    .X(net4850));
 sg13g2_dlygate4sd3_1 hold2254 (.A(_01850_),
    .X(net4851));
 sg13g2_dlygate4sd3_1 hold2255 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[29][18] ),
    .X(net4852));
 sg13g2_dlygate4sd3_1 hold2256 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[4] ),
    .X(net4853));
 sg13g2_dlygate4sd3_1 hold2257 (.A(_00908_),
    .X(net4854));
 sg13g2_dlygate4sd3_1 hold2258 (.A(\soc_I.clint_I.mtimecmp[8] ),
    .X(net4855));
 sg13g2_dlygate4sd3_1 hold2259 (.A(\soc_I.qqspi_I.xfer_cycles[2] ),
    .X(net4856));
 sg13g2_dlygate4sd3_1 hold2260 (.A(_00466_),
    .X(net4857));
 sg13g2_dlygate4sd3_1 hold2261 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[17] ),
    .X(net4858));
 sg13g2_dlygate4sd3_1 hold2262 (.A(\soc_I.clint_I.mtimecmp[52] ),
    .X(net4859));
 sg13g2_dlygate4sd3_1 hold2263 (.A(\soc_I.clint_I.mtimecmp[10] ),
    .X(net4860));
 sg13g2_dlygate4sd3_1 hold2264 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[25] ),
    .X(net4861));
 sg13g2_dlygate4sd3_1 hold2265 (.A(_04172_),
    .X(net4862));
 sg13g2_dlygate4sd3_1 hold2266 (.A(\gpio_uo_en[0] ),
    .X(net4863));
 sg13g2_dlygate4sd3_1 hold2267 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[25] ),
    .X(net4864));
 sg13g2_dlygate4sd3_1 hold2268 (.A(\soc_I.clint_I.mtimecmp[18] ),
    .X(net4865));
 sg13g2_dlygate4sd3_1 hold2269 (.A(\soc_I.rx_uart_i.wait_states[14] ),
    .X(net4866));
 sg13g2_dlygate4sd3_1 hold2270 (.A(_01856_),
    .X(net4867));
 sg13g2_dlygate4sd3_1 hold2271 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[18] ),
    .X(net4868));
 sg13g2_dlygate4sd3_1 hold2272 (.A(_00858_),
    .X(net4869));
 sg13g2_dlygate4sd3_1 hold2273 (.A(\soc_I.clint_I.mtimecmp[11] ),
    .X(net4870));
 sg13g2_dlygate4sd3_1 hold2274 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[13] ),
    .X(net4871));
 sg13g2_dlygate4sd3_1 hold2275 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[28] ),
    .X(net4872));
 sg13g2_dlygate4sd3_1 hold2276 (.A(_05500_),
    .X(net4873));
 sg13g2_dlygate4sd3_1 hold2277 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[29] ),
    .X(net4874));
 sg13g2_dlygate4sd3_1 hold2278 (.A(_01032_),
    .X(net4875));
 sg13g2_dlygate4sd3_1 hold2279 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[26] ),
    .X(net4876));
 sg13g2_dlygate4sd3_1 hold2280 (.A(_00930_),
    .X(net4877));
 sg13g2_dlygate4sd3_1 hold2281 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[1] ),
    .X(net4878));
 sg13g2_dlygate4sd3_1 hold2282 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[33] ),
    .X(net4879));
 sg13g2_dlygate4sd3_1 hold2283 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[0] ),
    .X(net4880));
 sg13g2_dlygate4sd3_1 hold2284 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[14] ),
    .X(net4881));
 sg13g2_dlygate4sd3_1 hold2285 (.A(_00918_),
    .X(net4882));
 sg13g2_dlygate4sd3_1 hold2286 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[17] ),
    .X(net4883));
 sg13g2_dlygate4sd3_1 hold2287 (.A(_00921_),
    .X(net4884));
 sg13g2_dlygate4sd3_1 hold2288 (.A(\soc_I.clint_I.tick_cnt[1] ),
    .X(net4885));
 sg13g2_dlygate4sd3_1 hold2289 (.A(_06223_),
    .X(net4886));
 sg13g2_dlygate4sd3_1 hold2290 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[58] ),
    .X(net4887));
 sg13g2_dlygate4sd3_1 hold2291 (.A(\soc_I.rx_uart_i.wait_states[6] ),
    .X(net4888));
 sg13g2_dlygate4sd3_1 hold2292 (.A(_01848_),
    .X(net4889));
 sg13g2_dlygate4sd3_1 hold2293 (.A(\soc_I.spi0_I.div[5] ),
    .X(net4890));
 sg13g2_dlygate4sd3_1 hold2294 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[3] ),
    .X(net4891));
 sg13g2_dlygate4sd3_1 hold2295 (.A(\gpio_uo_en[3] ),
    .X(net4892));
 sg13g2_dlygate4sd3_1 hold2296 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[45] ),
    .X(net4893));
 sg13g2_dlygate4sd3_1 hold2297 (.A(_05597_),
    .X(net4894));
 sg13g2_dlygate4sd3_1 hold2298 (.A(\soc_I.clint_I.mtimecmp[30] ),
    .X(net4895));
 sg13g2_dlygate4sd3_1 hold2299 (.A(_00167_),
    .X(net4896));
 sg13g2_dlygate4sd3_1 hold2300 (.A(_05450_),
    .X(net4897));
 sg13g2_dlygate4sd3_1 hold2301 (.A(\soc_I.kianv_I.datapath_unit_I.Result_I.d5[8] ),
    .X(net4898));
 sg13g2_dlygate4sd3_1 hold2302 (.A(\soc_I.clint_I.mtimecmp[34] ),
    .X(net4899));
 sg13g2_dlygate4sd3_1 hold2303 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[15] ),
    .X(net4900));
 sg13g2_dlygate4sd3_1 hold2304 (.A(\soc_I.clint_I.mtime[27] ),
    .X(net4901));
 sg13g2_dlygate4sd3_1 hold2305 (.A(_01659_),
    .X(net4902));
 sg13g2_dlygate4sd3_1 hold2306 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[4] ),
    .X(net4903));
 sg13g2_dlygate4sd3_1 hold2307 (.A(_04669_),
    .X(net4904));
 sg13g2_dlygate4sd3_1 hold2308 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[19] ),
    .X(net4905));
 sg13g2_dlygate4sd3_1 hold2309 (.A(_00923_),
    .X(net4906));
 sg13g2_dlygate4sd3_1 hold2310 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[11] ),
    .X(net4907));
 sg13g2_dlygate4sd3_1 hold2311 (.A(\soc_I.clint_I.mtimecmp[15] ),
    .X(net4908));
 sg13g2_dlygate4sd3_1 hold2312 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[27] ),
    .X(net4909));
 sg13g2_dlygate4sd3_1 hold2313 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[15] ),
    .X(net4910));
 sg13g2_dlygate4sd3_1 hold2314 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[16] ),
    .X(net4911));
 sg13g2_dlygate4sd3_1 hold2315 (.A(_05419_),
    .X(net4912));
 sg13g2_dlygate4sd3_1 hold2316 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[28] ),
    .X(net4913));
 sg13g2_dlygate4sd3_1 hold2317 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[13] ),
    .X(net4914));
 sg13g2_dlygate4sd3_1 hold2318 (.A(_05399_),
    .X(net4915));
 sg13g2_dlygate4sd3_1 hold2319 (.A(\soc_I.clint_I.mtimecmp[61] ),
    .X(net4916));
 sg13g2_dlygate4sd3_1 hold2320 (.A(_00158_),
    .X(net4917));
 sg13g2_dlygate4sd3_1 hold2321 (.A(_05514_),
    .X(net4918));
 sg13g2_dlygate4sd3_1 hold2322 (.A(\soc_I.clint_I.mtimecmp[58] ),
    .X(net4919));
 sg13g2_dlygate4sd3_1 hold2323 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[7] ),
    .X(net4920));
 sg13g2_dlygate4sd3_1 hold2324 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[11] ),
    .X(net4921));
 sg13g2_dlygate4sd3_1 hold2325 (.A(\soc_I.clint_I.mtimecmp[50] ),
    .X(net4922));
 sg13g2_dlygate4sd3_1 hold2326 (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[22] ),
    .X(net4923));
 sg13g2_dlygate4sd3_1 hold2327 (.A(\soc_I.clint_I.mtimecmp[9] ),
    .X(net4924));
 sg13g2_dlygate4sd3_1 hold2328 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[0] ),
    .X(net4925));
 sg13g2_dlygate4sd3_1 hold2329 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[50] ),
    .X(net4926));
 sg13g2_dlygate4sd3_1 hold2330 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[21] ),
    .X(net4927));
 sg13g2_dlygate4sd3_1 hold2331 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[52] ),
    .X(net4928));
 sg13g2_dlygate4sd3_1 hold2332 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[6] ),
    .X(net4929));
 sg13g2_dlygate4sd3_1 hold2333 (.A(\soc_I.clint_I.mtimecmp[47] ),
    .X(net4930));
 sg13g2_dlygate4sd3_1 hold2334 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.bit_idx[3] ),
    .X(net4931));
 sg13g2_dlygate4sd3_1 hold2335 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[18] ),
    .X(net4932));
 sg13g2_dlygate4sd3_1 hold2336 (.A(_04158_),
    .X(net4933));
 sg13g2_dlygate4sd3_1 hold2337 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[12] ),
    .X(net4934));
 sg13g2_dlygate4sd3_1 hold2338 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[17] ),
    .X(net4935));
 sg13g2_dlygate4sd3_1 hold2339 (.A(_04691_),
    .X(net4936));
 sg13g2_dlygate4sd3_1 hold2340 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[15] ),
    .X(net4937));
 sg13g2_dlygate4sd3_1 hold2341 (.A(\soc_I.clint_I.mtimecmp[16] ),
    .X(net4938));
 sg13g2_dlygate4sd3_1 hold2342 (.A(\soc_I.spi0_I.div[4] ),
    .X(net4939));
 sg13g2_dlygate4sd3_1 hold2343 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[39] ),
    .X(net4940));
 sg13g2_dlygate4sd3_1 hold2344 (.A(_05587_),
    .X(net4941));
 sg13g2_dlygate4sd3_1 hold2345 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[54] ),
    .X(net4942));
 sg13g2_dlygate4sd3_1 hold2346 (.A(_05611_),
    .X(net4943));
 sg13g2_dlygate4sd3_1 hold2347 (.A(\soc_I.clint_I.mtimecmp[44] ),
    .X(net4944));
 sg13g2_dlygate4sd3_1 hold2348 (.A(\soc_I.clint_I.mtimecmp[1] ),
    .X(net4945));
 sg13g2_dlygate4sd3_1 hold2349 (.A(\soc_I.clint_I.mtime[53] ),
    .X(net4946));
 sg13g2_dlygate4sd3_1 hold2350 (.A(\soc_I.clint_I.tick_cnt[14] ),
    .X(net4947));
 sg13g2_dlygate4sd3_1 hold2351 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor2_abs[23] ),
    .X(net4948));
 sg13g2_dlygate4sd3_1 hold2352 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[60] ),
    .X(net4949));
 sg13g2_dlygate4sd3_1 hold2353 (.A(_02148_),
    .X(net4950));
 sg13g2_dlygate4sd3_1 hold2354 (.A(\gpio_uo_en[6] ),
    .X(net4951));
 sg13g2_dlygate4sd3_1 hold2355 (.A(\soc_I.kianv_I.Instr[3] ),
    .X(net4952));
 sg13g2_dlygate4sd3_1 hold2356 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[35] ),
    .X(net4953));
 sg13g2_dlygate4sd3_1 hold2357 (.A(\soc_I.clint_I.tick_cnt[7] ),
    .X(net4954));
 sg13g2_dlygate4sd3_1 hold2358 (.A(\soc_I.clint_I.mtimecmp[13] ),
    .X(net4955));
 sg13g2_dlygate4sd3_1 hold2359 (.A(\soc_I.clint_I.mtimecmp[20] ),
    .X(net4956));
 sg13g2_dlygate4sd3_1 hold2360 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[8] ),
    .X(net4957));
 sg13g2_dlygate4sd3_1 hold2361 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[59] ),
    .X(net4958));
 sg13g2_dlygate4sd3_1 hold2362 (.A(_04797_),
    .X(net4959));
 sg13g2_dlygate4sd3_1 hold2363 (.A(_01196_),
    .X(net4960));
 sg13g2_dlygate4sd3_1 hold2364 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[23] ),
    .X(net4961));
 sg13g2_dlygate4sd3_1 hold2365 (.A(_05560_),
    .X(net4962));
 sg13g2_dlygate4sd3_1 hold2366 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[27] ),
    .X(net4963));
 sg13g2_dlygate4sd3_1 hold2367 (.A(_01030_),
    .X(net4964));
 sg13g2_dlygate4sd3_1 hold2368 (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[26] ),
    .X(net4965));
 sg13g2_dlygate4sd3_1 hold2369 (.A(\gpio_uo_out[3] ),
    .X(net4966));
 sg13g2_dlygate4sd3_1 hold2370 (.A(\gpio_uo_en[1] ),
    .X(net4967));
 sg13g2_dlygate4sd3_1 hold2371 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[16] ),
    .X(net4968));
 sg13g2_dlygate4sd3_1 hold2372 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[22] ),
    .X(net4969));
 sg13g2_dlygate4sd3_1 hold2373 (.A(\soc_I.gpio0_I.ready ),
    .X(net4970));
 sg13g2_dlygate4sd3_1 hold2374 (.A(\soc_I.clint_I.mtime[55] ),
    .X(net4971));
 sg13g2_dlygate4sd3_1 hold2375 (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[4] ),
    .X(net4972));
 sg13g2_dlygate4sd3_1 hold2376 (.A(_01443_),
    .X(net4973));
 sg13g2_dlygate4sd3_1 hold2377 (.A(\soc_I.clint_I.mtimecmp[43] ),
    .X(net4974));
 sg13g2_dlygate4sd3_1 hold2378 (.A(\soc_I.qqspi_I.spi_buf[24] ),
    .X(net4975));
 sg13g2_dlygate4sd3_1 hold2379 (.A(_07311_),
    .X(net4976));
 sg13g2_dlygate4sd3_1 hold2380 (.A(\soc_I.qqspi_I.state[1] ),
    .X(net4977));
 sg13g2_dlygate4sd3_1 hold2381 (.A(_12571_),
    .X(net4978));
 sg13g2_dlygate4sd3_1 hold2382 (.A(\soc_I.clint_I.mtimecmp[31] ),
    .X(net4979));
 sg13g2_dlygate4sd3_1 hold2383 (.A(\soc_I.PC[2] ),
    .X(net4980));
 sg13g2_dlygate4sd3_1 hold2384 (.A(\soc_I.PC[31] ),
    .X(net4981));
 sg13g2_dlygate4sd3_1 hold2385 (.A(_01470_),
    .X(net4982));
 sg13g2_dlygate4sd3_1 hold2386 (.A(\soc_I.rx_uart_i.wait_states[3] ),
    .X(net4983));
 sg13g2_dlygate4sd3_1 hold2387 (.A(_06877_),
    .X(net4984));
 sg13g2_dlygate4sd3_1 hold2388 (.A(_00245_),
    .X(net4985));
 sg13g2_dlygate4sd3_1 hold2389 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[5] ),
    .X(net4986));
 sg13g2_dlygate4sd3_1 hold2390 (.A(_05529_),
    .X(net4987));
 sg13g2_dlygate4sd3_1 hold2391 (.A(\soc_I.spi0_I.tick_cnt[0] ),
    .X(net4988));
 sg13g2_dlygate4sd3_1 hold2392 (.A(_06612_),
    .X(net4989));
 sg13g2_dlygate4sd3_1 hold2393 (.A(\soc_I.clint_I.tick_cnt[4] ),
    .X(net4990));
 sg13g2_dlygate4sd3_1 hold2394 (.A(\gpio_uo_en[5] ),
    .X(net4991));
 sg13g2_dlygate4sd3_1 hold2395 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[16] ),
    .X(net4992));
 sg13g2_dlygate4sd3_1 hold2396 (.A(_00920_),
    .X(net4993));
 sg13g2_dlygate4sd3_1 hold2397 (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[29] ),
    .X(net4994));
 sg13g2_dlygate4sd3_1 hold2398 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[6] ),
    .X(net4995));
 sg13g2_dlygate4sd3_1 hold2399 (.A(\soc_I.clint_I.mtime[32] ),
    .X(net4996));
 sg13g2_dlygate4sd3_1 hold2400 (.A(_06381_),
    .X(net4997));
 sg13g2_dlygate4sd3_1 hold2401 (.A(_01666_),
    .X(net4998));
 sg13g2_dlygate4sd3_1 hold2402 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[18] ),
    .X(net4999));
 sg13g2_dlygate4sd3_1 hold2403 (.A(_05432_),
    .X(net5000));
 sg13g2_dlygate4sd3_1 hold2404 (.A(\soc_I.div_reg[12] ),
    .X(net5001));
 sg13g2_dlygate4sd3_1 hold2405 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[3] ),
    .X(net5002));
 sg13g2_dlygate4sd3_1 hold2406 (.A(\soc_I.clint_I.mtime[21] ),
    .X(net5003));
 sg13g2_dlygate4sd3_1 hold2407 (.A(_01653_),
    .X(net5004));
 sg13g2_dlygate4sd3_1 hold2408 (.A(\soc_I.clint_I.mtimecmp[2] ),
    .X(net5005));
 sg13g2_dlygate4sd3_1 hold2409 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[8] ),
    .X(net5006));
 sg13g2_dlygate4sd3_1 hold2410 (.A(_04676_),
    .X(net5007));
 sg13g2_dlygate4sd3_1 hold2411 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[8] ),
    .X(net5008));
 sg13g2_dlygate4sd3_1 hold2412 (.A(\soc_I.spi0_I.div[7] ),
    .X(net5009));
 sg13g2_dlygate4sd3_1 hold2413 (.A(\gpio_uo_en[4] ),
    .X(net5010));
 sg13g2_dlygate4sd3_1 hold2414 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[51] ),
    .X(net5011));
 sg13g2_dlygate4sd3_1 hold2415 (.A(\soc_I.spi0_I.tick_cnt[5] ),
    .X(net5012));
 sg13g2_dlygate4sd3_1 hold2416 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[4] ),
    .X(net5013));
 sg13g2_dlygate4sd3_1 hold2417 (.A(_05528_),
    .X(net5014));
 sg13g2_dlygate4sd3_1 hold2418 (.A(\soc_I.rx_uart_i.wait_states[4] ),
    .X(net5015));
 sg13g2_dlygate4sd3_1 hold2419 (.A(_01846_),
    .X(net5016));
 sg13g2_dlygate4sd3_1 hold2420 (.A(\soc_I.clint_I.div[14] ),
    .X(net5017));
 sg13g2_dlygate4sd3_1 hold2421 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[29] ),
    .X(net5018));
 sg13g2_dlygate4sd3_1 hold2422 (.A(\soc_I.clint_I.mtimecmp[45] ),
    .X(net5019));
 sg13g2_dlygate4sd3_1 hold2423 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[10] ),
    .X(net5020));
 sg13g2_dlygate4sd3_1 hold2424 (.A(_05379_),
    .X(net5021));
 sg13g2_dlygate4sd3_1 hold2425 (.A(_00161_),
    .X(net5022));
 sg13g2_dlygate4sd3_1 hold2426 (.A(_05494_),
    .X(net5023));
 sg13g2_dlygate4sd3_1 hold2427 (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[28] ),
    .X(net5024));
 sg13g2_dlygate4sd3_1 hold2428 (.A(_01467_),
    .X(net5025));
 sg13g2_dlygate4sd3_1 hold2429 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[12] ),
    .X(net5026));
 sg13g2_dlygate4sd3_1 hold2430 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[9] ),
    .X(net5027));
 sg13g2_dlygate4sd3_1 hold2431 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[28] ),
    .X(net5028));
 sg13g2_dlygate4sd3_1 hold2432 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[13] ),
    .X(net5029));
 sg13g2_dlygate4sd3_1 hold2433 (.A(\soc_I.clint_I.mtimecmp[53] ),
    .X(net5030));
 sg13g2_dlygate4sd3_1 hold2434 (.A(\soc_I.clint_I.tick_cnt[5] ),
    .X(net5031));
 sg13g2_dlygate4sd3_1 hold2435 (.A(\soc_I.clint_I.mtimecmp[54] ),
    .X(net5032));
 sg13g2_dlygate4sd3_1 hold2436 (.A(\soc_I.clint_I.div[10] ),
    .X(net5033));
 sg13g2_dlygate4sd3_1 hold2437 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[57] ),
    .X(net5034));
 sg13g2_dlygate4sd3_1 hold2438 (.A(_04793_),
    .X(net5035));
 sg13g2_dlygate4sd3_1 hold2439 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[10] ),
    .X(net5036));
 sg13g2_dlygate4sd3_1 hold2440 (.A(\soc_I.spi0_I.div[3] ),
    .X(net5037));
 sg13g2_dlygate4sd3_1 hold2441 (.A(\soc_I.clint_I.mtimecmp[38] ),
    .X(net5038));
 sg13g2_dlygate4sd3_1 hold2442 (.A(\gpio_uo_en[2] ),
    .X(net5039));
 sg13g2_dlygate4sd3_1 hold2443 (.A(\soc_I.clint_I.mtimecmp[35] ),
    .X(net5040));
 sg13g2_dlygate4sd3_1 hold2444 (.A(\soc_I.spi0_I.xfer_cycles[1] ),
    .X(net5041));
 sg13g2_dlygate4sd3_1 hold2445 (.A(_06568_),
    .X(net5042));
 sg13g2_dlygate4sd3_1 hold2446 (.A(_06570_),
    .X(net5043));
 sg13g2_dlygate4sd3_1 hold2447 (.A(\soc_I.spi0_I.xfer_cycles[0] ),
    .X(net5044));
 sg13g2_dlygate4sd3_1 hold2448 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[44] ),
    .X(net5045));
 sg13g2_dlygate4sd3_1 hold2449 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[19] ),
    .X(net5046));
 sg13g2_dlygate4sd3_1 hold2450 (.A(\soc_I.clint_I.div[11] ),
    .X(net5047));
 sg13g2_dlygate4sd3_1 hold2451 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.state[0] ),
    .X(net5048));
 sg13g2_dlygate4sd3_1 hold2452 (.A(_05755_),
    .X(net5049));
 sg13g2_dlygate4sd3_1 hold2453 (.A(\soc_I.qqspi_I.xfer_cycles[4] ),
    .X(net5050));
 sg13g2_dlygate4sd3_1 hold2454 (.A(_00468_),
    .X(net5051));
 sg13g2_dlygate4sd3_1 hold2455 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[4] ),
    .X(net5052));
 sg13g2_dlygate4sd3_1 hold2456 (.A(_05337_),
    .X(net5053));
 sg13g2_dlygate4sd3_1 hold2457 (.A(\soc_I.kianv_I.Instr[10] ),
    .X(net5054));
 sg13g2_dlygate4sd3_1 hold2458 (.A(\soc_I.clint_I.mtimecmp[62] ),
    .X(net5055));
 sg13g2_dlygate4sd3_1 hold2459 (.A(\soc_I.kianv_I.datapath_unit_I.ALUOut[1] ),
    .X(net5056));
 sg13g2_dlygate4sd3_1 hold2460 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[19] ),
    .X(net5057));
 sg13g2_dlygate4sd3_1 hold2461 (.A(_05438_),
    .X(net5058));
 sg13g2_dlygate4sd3_1 hold2462 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[4] ),
    .X(net5059));
 sg13g2_dlygate4sd3_1 hold2463 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[26] ),
    .X(net5060));
 sg13g2_dlygate4sd3_1 hold2464 (.A(\soc_I.clint_I.mtime[39] ),
    .X(net5061));
 sg13g2_dlygate4sd3_1 hold2465 (.A(_06393_),
    .X(net5062));
 sg13g2_dlygate4sd3_1 hold2466 (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[14] ),
    .X(net5063));
 sg13g2_dlygate4sd3_1 hold2467 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[7] ),
    .X(net5064));
 sg13g2_dlygate4sd3_1 hold2468 (.A(\soc_I.rst_cnt[2] ),
    .X(net5065));
 sg13g2_dlygate4sd3_1 hold2469 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[1] ),
    .X(net5066));
 sg13g2_dlygate4sd3_1 hold2470 (.A(\soc_I.qqspi_I.state[0] ),
    .X(net5067));
 sg13g2_dlygate4sd3_1 hold2471 (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[1] ),
    .X(net5068));
 sg13g2_dlygate4sd3_1 hold2472 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[4] ),
    .X(net5069));
 sg13g2_dlygate4sd3_1 hold2473 (.A(_02204_),
    .X(net5070));
 sg13g2_dlygate4sd3_1 hold2474 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[1] ),
    .X(net5071));
 sg13g2_dlygate4sd3_1 hold2475 (.A(_04663_),
    .X(net5072));
 sg13g2_dlygate4sd3_1 hold2476 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[58] ),
    .X(net5073));
 sg13g2_dlygate4sd3_1 hold2477 (.A(\soc_I.clint_I.div[7] ),
    .X(net5074));
 sg13g2_dlygate4sd3_1 hold2478 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[55] ),
    .X(net5075));
 sg13g2_dlygate4sd3_1 hold2479 (.A(_04787_),
    .X(net5076));
 sg13g2_dlygate4sd3_1 hold2480 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[2] ),
    .X(net5077));
 sg13g2_dlygate4sd3_1 hold2481 (.A(\soc_I.clint_I.mtimecmp[24] ),
    .X(net5078));
 sg13g2_dlygate4sd3_1 hold2482 (.A(\soc_I.clint_I.mtime[48] ),
    .X(net5079));
 sg13g2_dlygate4sd3_1 hold2483 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[38] ),
    .X(net5080));
 sg13g2_dlygate4sd3_1 hold2484 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[22] ),
    .X(net5081));
 sg13g2_dlygate4sd3_1 hold2485 (.A(_05458_),
    .X(net5082));
 sg13g2_dlygate4sd3_1 hold2486 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[9] ),
    .X(net5083));
 sg13g2_dlygate4sd3_1 hold2487 (.A(_02199_),
    .X(net5084));
 sg13g2_dlygate4sd3_1 hold2488 (.A(\soc_I.clint_I.mtimecmp[22] ),
    .X(net5085));
 sg13g2_dlygate4sd3_1 hold2489 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[60] ),
    .X(net5086));
 sg13g2_dlygate4sd3_1 hold2490 (.A(\soc_I.clint_I.mtime[8] ),
    .X(net5087));
 sg13g2_dlygate4sd3_1 hold2491 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[7] ),
    .X(net5088));
 sg13g2_dlygate4sd3_1 hold2492 (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[26] ),
    .X(net5089));
 sg13g2_dlygate4sd3_1 hold2493 (.A(_01465_),
    .X(net5090));
 sg13g2_dlygate4sd3_1 hold2494 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[2] ),
    .X(net5091));
 sg13g2_dlygate4sd3_1 hold2495 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[19] ),
    .X(net5092));
 sg13g2_dlygate4sd3_1 hold2496 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[52] ),
    .X(net5093));
 sg13g2_dlygate4sd3_1 hold2497 (.A(_01189_),
    .X(net5094));
 sg13g2_dlygate4sd3_1 hold2498 (.A(\soc_I.clint_I.mtimecmp[25] ),
    .X(net5095));
 sg13g2_dlygate4sd3_1 hold2499 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[1] ),
    .X(net5096));
 sg13g2_dlygate4sd3_1 hold2500 (.A(\soc_I.PC[27] ),
    .X(net5097));
 sg13g2_dlygate4sd3_1 hold2501 (.A(\soc_I.clint_I.tick_cnt[13] ),
    .X(net5098));
 sg13g2_dlygate4sd3_1 hold2502 (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[21] ),
    .X(net5099));
 sg13g2_dlygate4sd3_1 hold2503 (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[19] ),
    .X(net5100));
 sg13g2_dlygate4sd3_1 hold2504 (.A(\soc_I.clint_I.mtimecmp[57] ),
    .X(net5101));
 sg13g2_dlygate4sd3_1 hold2505 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[59] ),
    .X(net5102));
 sg13g2_dlygate4sd3_1 hold2506 (.A(_02149_),
    .X(net5103));
 sg13g2_dlygate4sd3_1 hold2507 (.A(\soc_I.qqspi_I.xfer_cycles[5] ),
    .X(net5104));
 sg13g2_dlygate4sd3_1 hold2508 (.A(_00469_),
    .X(net5105));
 sg13g2_dlygate4sd3_1 hold2509 (.A(\soc_I.rx_uart_i.fifo_i.cnt[4] ),
    .X(net5106));
 sg13g2_dlygate4sd3_1 hold2510 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[20] ),
    .X(net5107));
 sg13g2_dlygate4sd3_1 hold2511 (.A(\soc_I.spi0_I.div[6] ),
    .X(net5108));
 sg13g2_dlygate4sd3_1 hold2512 (.A(\soc_I.rx_uart_i.wait_states[9] ),
    .X(net5109));
 sg13g2_dlygate4sd3_1 hold2513 (.A(_01851_),
    .X(net5110));
 sg13g2_dlygate4sd3_1 hold2514 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[57] ),
    .X(net5111));
 sg13g2_dlygate4sd3_1 hold2515 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[16] ),
    .X(net5112));
 sg13g2_dlygate4sd3_1 hold2516 (.A(\soc_I.clint_I.mtime[56] ),
    .X(net5113));
 sg13g2_dlygate4sd3_1 hold2517 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[38] ),
    .X(net5114));
 sg13g2_dlygate4sd3_1 hold2518 (.A(_02170_),
    .X(net5115));
 sg13g2_dlygate4sd3_1 hold2519 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[28] ),
    .X(net5116));
 sg13g2_dlygate4sd3_1 hold2520 (.A(\soc_I.clint_I.mtime[42] ),
    .X(net5117));
 sg13g2_dlygate4sd3_1 hold2521 (.A(\soc_I.clint_I.tick_cnt[16] ),
    .X(net5118));
 sg13g2_dlygate4sd3_1 hold2522 (.A(\soc_I.clint_I.mtime[20] ),
    .X(net5119));
 sg13g2_dlygate4sd3_1 hold2523 (.A(_01652_),
    .X(net5120));
 sg13g2_dlygate4sd3_1 hold2524 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[18] ),
    .X(net5121));
 sg13g2_dlygate4sd3_1 hold2525 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[30] ),
    .X(net5122));
 sg13g2_dlygate4sd3_1 hold2526 (.A(\soc_I.spi0_I.div[12] ),
    .X(net5123));
 sg13g2_dlygate4sd3_1 hold2527 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[6] ),
    .X(net5124));
 sg13g2_dlygate4sd3_1 hold2528 (.A(\soc_I.clint_I.mtime[10] ),
    .X(net5125));
 sg13g2_dlygate4sd3_1 hold2529 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[26] ),
    .X(net5126));
 sg13g2_dlygate4sd3_1 hold2530 (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[22] ),
    .X(net5127));
 sg13g2_dlygate4sd3_1 hold2531 (.A(_01461_),
    .X(net5128));
 sg13g2_dlygate4sd3_1 hold2532 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.factor1_abs[25] ),
    .X(net5129));
 sg13g2_dlygate4sd3_1 hold2533 (.A(\soc_I.qqspi_I.spi_buf[25] ),
    .X(net5130));
 sg13g2_dlygate4sd3_1 hold2534 (.A(_07317_),
    .X(net5131));
 sg13g2_dlygate4sd3_1 hold2535 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[63] ),
    .X(net5132));
 sg13g2_dlygate4sd3_1 hold2536 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[30] ),
    .X(net5133));
 sg13g2_dlygate4sd3_1 hold2537 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[31] ),
    .X(net5134));
 sg13g2_dlygate4sd3_1 hold2538 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[21] ),
    .X(net5135));
 sg13g2_dlygate4sd3_1 hold2539 (.A(\soc_I.clint_I.mtimecmp[26] ),
    .X(net5136));
 sg13g2_dlygate4sd3_1 hold2540 (.A(\soc_I.clint_I.mtimecmp[63] ),
    .X(net5137));
 sg13g2_dlygate4sd3_1 hold2541 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[17] ),
    .X(net5138));
 sg13g2_dlygate4sd3_1 hold2542 (.A(_05425_),
    .X(net5139));
 sg13g2_dlygate4sd3_1 hold2543 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mie[3] ),
    .X(net5140));
 sg13g2_dlygate4sd3_1 hold2544 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[18] ),
    .X(net5141));
 sg13g2_dlygate4sd3_1 hold2545 (.A(\soc_I.rx_uart_i.rx_in_sync[2] ),
    .X(net5142));
 sg13g2_dlygate4sd3_1 hold2546 (.A(_06810_),
    .X(net5143));
 sg13g2_dlygate4sd3_1 hold2547 (.A(_01828_),
    .X(net5144));
 sg13g2_dlygate4sd3_1 hold2548 (.A(\soc_I.IRQ3 ),
    .X(net5145));
 sg13g2_dlygate4sd3_1 hold2549 (.A(\soc_I.clint_I.div[2] ),
    .X(net5146));
 sg13g2_dlygate4sd3_1 hold2550 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[14] ),
    .X(net5147));
 sg13g2_dlygate4sd3_1 hold2551 (.A(\soc_I.clint_I.div[15] ),
    .X(net5148));
 sg13g2_dlygate4sd3_1 hold2552 (.A(\soc_I.clint_I.mtime[40] ),
    .X(net5149));
 sg13g2_dlygate4sd3_1 hold2553 (.A(_06395_),
    .X(net5150));
 sg13g2_dlygate4sd3_1 hold2554 (.A(\gpio_uo_en[7] ),
    .X(net5151));
 sg13g2_dlygate4sd3_1 hold2555 (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[24] ),
    .X(net5152));
 sg13g2_dlygate4sd3_1 hold2556 (.A(\soc_I.spi0_I.div[2] ),
    .X(net5153));
 sg13g2_dlygate4sd3_1 hold2557 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[3] ),
    .X(net5154));
 sg13g2_dlygate4sd3_1 hold2558 (.A(_05329_),
    .X(net5155));
 sg13g2_dlygate4sd3_1 hold2559 (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[16] ),
    .X(net5156));
 sg13g2_dlygate4sd3_1 hold2560 (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[6] ),
    .X(net5157));
 sg13g2_dlygate4sd3_1 hold2561 (.A(_01445_),
    .X(net5158));
 sg13g2_dlygate4sd3_1 hold2562 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[22] ),
    .X(net5159));
 sg13g2_dlygate4sd3_1 hold2563 (.A(_04704_),
    .X(net5160));
 sg13g2_dlygate4sd3_1 hold2564 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[20] ),
    .X(net5161));
 sg13g2_dlygate4sd3_1 hold2565 (.A(\soc_I.rx_uart_i.wait_states[7] ),
    .X(net5162));
 sg13g2_dlygate4sd3_1 hold2566 (.A(_01849_),
    .X(net5163));
 sg13g2_dlygate4sd3_1 hold2567 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[17] ),
    .X(net5164));
 sg13g2_dlygate4sd3_1 hold2568 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[22] ),
    .X(net5165));
 sg13g2_dlygate4sd3_1 hold2569 (.A(\soc_I.clint_I.mtime[37] ),
    .X(net5166));
 sg13g2_dlygate4sd3_1 hold2570 (.A(_01669_),
    .X(net5167));
 sg13g2_dlygate4sd3_1 hold2571 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[10] ),
    .X(net5168));
 sg13g2_dlygate4sd3_1 hold2572 (.A(\soc_I.clint_I.mtime[43] ),
    .X(net5169));
 sg13g2_dlygate4sd3_1 hold2573 (.A(_01676_),
    .X(net5170));
 sg13g2_dlygate4sd3_1 hold2574 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[20] ),
    .X(net5171));
 sg13g2_dlygate4sd3_1 hold2575 (.A(_05443_),
    .X(net5172));
 sg13g2_dlygate4sd3_1 hold2576 (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[18] ),
    .X(net5173));
 sg13g2_dlygate4sd3_1 hold2577 (.A(\soc_I.clint_I.mtime[50] ),
    .X(net5174));
 sg13g2_dlygate4sd3_1 hold2578 (.A(_06419_),
    .X(net5175));
 sg13g2_dlygate4sd3_1 hold2579 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[59] ),
    .X(net5176));
 sg13g2_dlygate4sd3_1 hold2580 (.A(\soc_I.rx_uart_i.wait_states[13] ),
    .X(net5177));
 sg13g2_dlygate4sd3_1 hold2581 (.A(_01855_),
    .X(net5178));
 sg13g2_dlygate4sd3_1 hold2582 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[45] ),
    .X(net5179));
 sg13g2_dlygate4sd3_1 hold2583 (.A(\soc_I.qqspi_I.spi_buf[27] ),
    .X(net5180));
 sg13g2_dlygate4sd3_1 hold2584 (.A(_07330_),
    .X(net5181));
 sg13g2_dlygate4sd3_1 hold2585 (.A(\soc_I.qqspi_I.xfer_cycles[3] ),
    .X(net5182));
 sg13g2_dlygate4sd3_1 hold2586 (.A(\soc_I.rx_uart_i.fifo_i.wr_ptr[3] ),
    .X(net5183));
 sg13g2_dlygate4sd3_1 hold2587 (.A(_06950_),
    .X(net5184));
 sg13g2_dlygate4sd3_1 hold2588 (.A(\soc_I.clint_I.div[6] ),
    .X(net5185));
 sg13g2_dlygate4sd3_1 hold2589 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[24] ),
    .X(net5186));
 sg13g2_dlygate4sd3_1 hold2590 (.A(_01257_),
    .X(net5187));
 sg13g2_dlygate4sd3_1 hold2591 (.A(\soc_I.clint_I.mtime[12] ),
    .X(net5188));
 sg13g2_dlygate4sd3_1 hold2592 (.A(_01644_),
    .X(net5189));
 sg13g2_dlygate4sd3_1 hold2593 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[27] ),
    .X(net5190));
 sg13g2_dlygate4sd3_1 hold2594 (.A(\soc_I.qqspi_I.spi_buf[8] ),
    .X(net5191));
 sg13g2_dlygate4sd3_1 hold2595 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[25] ),
    .X(net5192));
 sg13g2_dlygate4sd3_1 hold2596 (.A(_02183_),
    .X(net5193));
 sg13g2_dlygate4sd3_1 hold2597 (.A(\soc_I.clint_I.mtime[26] ),
    .X(net5194));
 sg13g2_dlygate4sd3_1 hold2598 (.A(_06361_),
    .X(net5195));
 sg13g2_dlygate4sd3_1 hold2599 (.A(_01658_),
    .X(net5196));
 sg13g2_dlygate4sd3_1 hold2600 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[7] ),
    .X(net5197));
 sg13g2_dlygate4sd3_1 hold2601 (.A(\soc_I.qqspi_I.spi_buf[5] ),
    .X(net5198));
 sg13g2_dlygate4sd3_1 hold2602 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[37] ),
    .X(net5199));
 sg13g2_dlygate4sd3_1 hold2603 (.A(_04745_),
    .X(net5200));
 sg13g2_dlygate4sd3_1 hold2604 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[2] ),
    .X(net5201));
 sg13g2_dlygate4sd3_1 hold2605 (.A(_02206_),
    .X(net5202));
 sg13g2_dlygate4sd3_1 hold2606 (.A(\soc_I.rx_uart_i.fifo_i.cnt[1] ),
    .X(net5203));
 sg13g2_dlygate4sd3_1 hold2607 (.A(_06653_),
    .X(net5204));
 sg13g2_dlygate4sd3_1 hold2608 (.A(_01783_),
    .X(net5205));
 sg13g2_dlygate4sd3_1 hold2609 (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[23] ),
    .X(net5206));
 sg13g2_dlygate4sd3_1 hold2610 (.A(\soc_I.tx_uart_i.tx_out ),
    .X(net5207));
 sg13g2_dlygate4sd3_1 hold2611 (.A(_01871_),
    .X(net5208));
 sg13g2_dlygate4sd3_1 hold2612 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[21] ),
    .X(net5209));
 sg13g2_dlygate4sd3_1 hold2613 (.A(\soc_I.spi0_I.div[1] ),
    .X(net5210));
 sg13g2_dlygate4sd3_1 hold2614 (.A(\led[1] ),
    .X(net5211));
 sg13g2_dlygate4sd3_1 hold2615 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[19] ),
    .X(net5212));
 sg13g2_dlygate4sd3_1 hold2616 (.A(_01220_),
    .X(net5213));
 sg13g2_dlygate4sd3_1 hold2617 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[3] ),
    .X(net5214));
 sg13g2_dlygate4sd3_1 hold2618 (.A(\soc_I.rx_uart_i.ready ),
    .X(net5215));
 sg13g2_dlygate4sd3_1 hold2619 (.A(_01795_),
    .X(net5216));
 sg13g2_dlygate4sd3_1 hold2620 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[29] ),
    .X(net5217));
 sg13g2_dlygate4sd3_1 hold2621 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtval[1] ),
    .X(net5218));
 sg13g2_dlygate4sd3_1 hold2622 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[30] ),
    .X(net5219));
 sg13g2_dlygate4sd3_1 hold2623 (.A(\soc_I.rx_uart_i.wait_states[0] ),
    .X(net5220));
 sg13g2_dlygate4sd3_1 hold2624 (.A(_01842_),
    .X(net5221));
 sg13g2_dlygate4sd3_1 hold2625 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[28] ),
    .X(net5222));
 sg13g2_dlygate4sd3_1 hold2626 (.A(_01229_),
    .X(net5223));
 sg13g2_dlygate4sd3_1 hold2627 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[10] ),
    .X(net5224));
 sg13g2_dlygate4sd3_1 hold2628 (.A(_01211_),
    .X(net5225));
 sg13g2_dlygate4sd3_1 hold2629 (.A(\led[0] ),
    .X(net5226));
 sg13g2_dlygate4sd3_1 hold2630 (.A(_01455_),
    .X(net5227));
 sg13g2_dlygate4sd3_1 hold2631 (.A(\soc_I.rx_uart_i.wait_states[11] ),
    .X(net5228));
 sg13g2_dlygate4sd3_1 hold2632 (.A(_06921_),
    .X(net5229));
 sg13g2_dlygate4sd3_1 hold2633 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[8] ),
    .X(net5230));
 sg13g2_dlygate4sd3_1 hold2634 (.A(_01209_),
    .X(net5231));
 sg13g2_dlygate4sd3_1 hold2635 (.A(\soc_I.div_reg[11] ),
    .X(net5232));
 sg13g2_dlygate4sd3_1 hold2636 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[8] ),
    .X(net5233));
 sg13g2_dlygate4sd3_1 hold2637 (.A(\soc_I.spi0_I.div[10] ),
    .X(net5234));
 sg13g2_dlygate4sd3_1 hold2638 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[10] ),
    .X(net5235));
 sg13g2_dlygate4sd3_1 hold2639 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[12] ),
    .X(net5236));
 sg13g2_dlygate4sd3_1 hold2640 (.A(\soc_I.kianv_I.Instr[27] ),
    .X(net5237));
 sg13g2_dlygate4sd3_1 hold2641 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[28] ),
    .X(net5238));
 sg13g2_dlygate4sd3_1 hold2642 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[2] ),
    .X(net5239));
 sg13g2_dlygate4sd3_1 hold2643 (.A(_05323_),
    .X(net5240));
 sg13g2_dlygate4sd3_1 hold2644 (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[5] ),
    .X(net5241));
 sg13g2_dlygate4sd3_1 hold2645 (.A(_01444_),
    .X(net5242));
 sg13g2_dlygate4sd3_1 hold2646 (.A(\soc_I.clint_I.mtime[14] ),
    .X(net5243));
 sg13g2_dlygate4sd3_1 hold2647 (.A(_01646_),
    .X(net5244));
 sg13g2_dlygate4sd3_1 hold2648 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[27] ),
    .X(net5245));
 sg13g2_dlygate4sd3_1 hold2649 (.A(\soc_I.rx_uart_i.wait_states[1] ),
    .X(net5246));
 sg13g2_dlygate4sd3_1 hold2650 (.A(_01843_),
    .X(net5247));
 sg13g2_dlygate4sd3_1 hold2651 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[22] ),
    .X(net5248));
 sg13g2_dlygate4sd3_1 hold2652 (.A(_01223_),
    .X(net5249));
 sg13g2_dlygate4sd3_1 hold2653 (.A(\soc_I.div_reg[14] ),
    .X(net5250));
 sg13g2_dlygate4sd3_1 hold2654 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[23] ),
    .X(net5251));
 sg13g2_dlygate4sd3_1 hold2655 (.A(\soc_I.clint_I.div[9] ),
    .X(net5252));
 sg13g2_dlygate4sd3_1 hold2656 (.A(\soc_I.div_reg[10] ),
    .X(net5253));
 sg13g2_dlygate4sd3_1 hold2657 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[26] ),
    .X(net5254));
 sg13g2_dlygate4sd3_1 hold2658 (.A(\soc_I.PC[21] ),
    .X(net5255));
 sg13g2_dlygate4sd3_1 hold2659 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[6] ),
    .X(net5256));
 sg13g2_dlygate4sd3_1 hold2660 (.A(_01207_),
    .X(net5257));
 sg13g2_dlygate4sd3_1 hold2661 (.A(\soc_I.PC[23] ),
    .X(net5258));
 sg13g2_dlygate4sd3_1 hold2662 (.A(_01559_),
    .X(net5259));
 sg13g2_dlygate4sd3_1 hold2663 (.A(\soc_I.clint_I.div[13] ),
    .X(net5260));
 sg13g2_dlygate4sd3_1 hold2664 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[30] ),
    .X(net5261));
 sg13g2_dlygate4sd3_1 hold2665 (.A(_01231_),
    .X(net5262));
 sg13g2_dlygate4sd3_1 hold2666 (.A(\soc_I.PC[26] ),
    .X(net5263));
 sg13g2_dlygate4sd3_1 hold2667 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[15] ),
    .X(net5264));
 sg13g2_dlygate4sd3_1 hold2668 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[7] ),
    .X(net5265));
 sg13g2_dlygate4sd3_1 hold2669 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[11] ),
    .X(net5266));
 sg13g2_dlygate4sd3_1 hold2670 (.A(\soc_I.rx_uart_i.wait_states[5] ),
    .X(net5267));
 sg13g2_dlygate4sd3_1 hold2671 (.A(_06889_),
    .X(net5268));
 sg13g2_dlygate4sd3_1 hold2672 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[4] ),
    .X(net5269));
 sg13g2_dlygate4sd3_1 hold2673 (.A(\soc_I.clint_I.tick_cnt[9] ),
    .X(net5270));
 sg13g2_dlygate4sd3_1 hold2674 (.A(\soc_I.div_reg[8] ),
    .X(net5271));
 sg13g2_dlygate4sd3_1 hold2675 (.A(\soc_I.PC[6] ),
    .X(net5272));
 sg13g2_dlygate4sd3_1 hold2676 (.A(\soc_I.qqspi_I.spi_buf[16] ),
    .X(net5273));
 sg13g2_dlygate4sd3_1 hold2677 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[44] ),
    .X(net5274));
 sg13g2_dlygate4sd3_1 hold2678 (.A(_04763_),
    .X(net5275));
 sg13g2_dlygate4sd3_1 hold2679 (.A(\soc_I.spi0_I.div[14] ),
    .X(net5276));
 sg13g2_dlygate4sd3_1 hold2680 (.A(\soc_I.qqspi_I.spi_buf[15] ),
    .X(net5277));
 sg13g2_dlygate4sd3_1 hold2681 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[14] ),
    .X(net5278));
 sg13g2_dlygate4sd3_1 hold2682 (.A(\soc_I.PC[11] ),
    .X(net5279));
 sg13g2_dlygate4sd3_1 hold2683 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[5] ),
    .X(net5280));
 sg13g2_dlygate4sd3_1 hold2684 (.A(_05345_),
    .X(net5281));
 sg13g2_dlygate4sd3_1 hold2685 (.A(\soc_I.spi0_I.div[9] ),
    .X(net5282));
 sg13g2_dlygate4sd3_1 hold2686 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[7] ),
    .X(net5283));
 sg13g2_dlygate4sd3_1 hold2687 (.A(_01208_),
    .X(net5284));
 sg13g2_dlygate4sd3_1 hold2688 (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[17] ),
    .X(net5285));
 sg13g2_dlygate4sd3_1 hold2689 (.A(\soc_I.qqspi_I.spi_buf[18] ),
    .X(net5286));
 sg13g2_dlygate4sd3_1 hold2690 (.A(\soc_I.qqspi_I.spi_buf[4] ),
    .X(net5287));
 sg13g2_dlygate4sd3_1 hold2691 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[46] ),
    .X(net5288));
 sg13g2_dlygate4sd3_1 hold2692 (.A(\soc_I.tx_uart_i.return_state[1] ),
    .X(net5289));
 sg13g2_dlygate4sd3_1 hold2693 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[4] ),
    .X(net5290));
 sg13g2_dlygate4sd3_1 hold2694 (.A(_01205_),
    .X(net5291));
 sg13g2_dlygate4sd3_1 hold2695 (.A(\soc_I.clint_I.div[3] ),
    .X(net5292));
 sg13g2_dlygate4sd3_1 hold2696 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[3] ),
    .X(net5293));
 sg13g2_dlygate4sd3_1 hold2697 (.A(_05525_),
    .X(net5294));
 sg13g2_dlygate4sd3_1 hold2698 (.A(\soc_I.clint_I.mtimecmp[23] ),
    .X(net5295));
 sg13g2_dlygate4sd3_1 hold2699 (.A(\soc_I.PC[22] ),
    .X(net5296));
 sg13g2_dlygate4sd3_1 hold2700 (.A(\soc_I.clint_I.mtime[24] ),
    .X(net5297));
 sg13g2_dlygate4sd3_1 hold2701 (.A(_06355_),
    .X(net5298));
 sg13g2_dlygate4sd3_1 hold2702 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[21] ),
    .X(net5299));
 sg13g2_dlygate4sd3_1 hold2703 (.A(\soc_I.qqspi_I.spi_buf[17] ),
    .X(net5300));
 sg13g2_dlygate4sd3_1 hold2704 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[9] ),
    .X(net5301));
 sg13g2_dlygate4sd3_1 hold2705 (.A(\soc_I.kianv_I.control_unit_I.div_ready ),
    .X(net5302));
 sg13g2_dlygate4sd3_1 hold2706 (.A(_05645_),
    .X(net5303));
 sg13g2_dlygate4sd3_1 hold2707 (.A(\soc_I.spi0_I.div[13] ),
    .X(net5304));
 sg13g2_dlygate4sd3_1 hold2708 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[16] ),
    .X(net5305));
 sg13g2_dlygate4sd3_1 hold2709 (.A(_01217_),
    .X(net5306));
 sg13g2_dlygate4sd3_1 hold2710 (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[17] ),
    .X(net5307));
 sg13g2_dlygate4sd3_1 hold2711 (.A(\led[3] ),
    .X(net5308));
 sg13g2_dlygate4sd3_1 hold2712 (.A(_01458_),
    .X(net5309));
 sg13g2_dlygate4sd3_1 hold2713 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[8] ),
    .X(net5310));
 sg13g2_dlygate4sd3_1 hold2714 (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[25] ),
    .X(net5311));
 sg13g2_dlygate4sd3_1 hold2715 (.A(_01464_),
    .X(net5312));
 sg13g2_dlygate4sd3_1 hold2716 (.A(\soc_I.div_reg[13] ),
    .X(net5313));
 sg13g2_dlygate4sd3_1 hold2717 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[35] ),
    .X(net5314));
 sg13g2_dlygate4sd3_1 hold2718 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[25] ),
    .X(net5315));
 sg13g2_dlygate4sd3_1 hold2719 (.A(_01226_),
    .X(net5316));
 sg13g2_dlygate4sd3_1 hold2720 (.A(\soc_I.clint_I.mtime[41] ),
    .X(net5317));
 sg13g2_dlygate4sd3_1 hold2721 (.A(_01673_),
    .X(net5318));
 sg13g2_dlygate4sd3_1 hold2722 (.A(\soc_I.div_reg[7] ),
    .X(net5319));
 sg13g2_dlygate4sd3_1 hold2723 (.A(\soc_I.qqspi_I.spi_buf[6] ),
    .X(net5320));
 sg13g2_dlygate4sd3_1 hold2724 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[20] ),
    .X(net5321));
 sg13g2_dlygate4sd3_1 hold2725 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[25] ),
    .X(net5322));
 sg13g2_dlygate4sd3_1 hold2726 (.A(\soc_I.PC[5] ),
    .X(net5323));
 sg13g2_dlygate4sd3_1 hold2727 (.A(_01541_),
    .X(net5324));
 sg13g2_dlygate4sd3_1 hold2728 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[3] ),
    .X(net5325));
 sg13g2_dlygate4sd3_1 hold2729 (.A(_01204_),
    .X(net5326));
 sg13g2_dlygate4sd3_1 hold2730 (.A(\soc_I.div_reg[6] ),
    .X(net5327));
 sg13g2_dlygate4sd3_1 hold2731 (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[8] ),
    .X(net5328));
 sg13g2_dlygate4sd3_1 hold2732 (.A(_01447_),
    .X(net5329));
 sg13g2_dlygate4sd3_1 hold2733 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[9] ),
    .X(net5330));
 sg13g2_dlygate4sd3_1 hold2734 (.A(_01545_),
    .X(net5331));
 sg13g2_dlygate4sd3_1 hold2735 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[11] ),
    .X(net5332));
 sg13g2_dlygate4sd3_1 hold2736 (.A(_05385_),
    .X(net5333));
 sg13g2_dlygate4sd3_1 hold2737 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[28] ),
    .X(net5334));
 sg13g2_dlygate4sd3_1 hold2738 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[31] ),
    .X(net5335));
 sg13g2_dlygate4sd3_1 hold2739 (.A(_02177_),
    .X(net5336));
 sg13g2_dlygate4sd3_1 hold2740 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[14] ),
    .X(net5337));
 sg13g2_dlygate4sd3_1 hold2741 (.A(_05406_),
    .X(net5338));
 sg13g2_dlygate4sd3_1 hold2742 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[3] ),
    .X(net5339));
 sg13g2_dlygate4sd3_1 hold2743 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[37] ),
    .X(net5340));
 sg13g2_dlygate4sd3_1 hold2744 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[34] ),
    .X(net5341));
 sg13g2_dlygate4sd3_1 hold2745 (.A(_01171_),
    .X(net5342));
 sg13g2_dlygate4sd3_1 hold2746 (.A(\soc_I.rx_uart_i.wait_states[12] ),
    .X(net5343));
 sg13g2_dlygate4sd3_1 hold2747 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[42] ),
    .X(net5344));
 sg13g2_dlygate4sd3_1 hold2748 (.A(_01179_),
    .X(net5345));
 sg13g2_dlygate4sd3_1 hold2749 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[11] ),
    .X(net5346));
 sg13g2_dlygate4sd3_1 hold2750 (.A(\soc_I.qqspi_I.spi_buf[13] ),
    .X(net5347));
 sg13g2_dlygate4sd3_1 hold2751 (.A(\soc_I.qqspi_I.spi_buf[7] ),
    .X(net5348));
 sg13g2_dlygate4sd3_1 hold2752 (.A(_02552_),
    .X(net5349));
 sg13g2_dlygate4sd3_1 hold2753 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[21] ),
    .X(net5350));
 sg13g2_dlygate4sd3_1 hold2754 (.A(\soc_I.qqspi_I.spi_buf[19] ),
    .X(net5351));
 sg13g2_dlygate4sd3_1 hold2755 (.A(\soc_I.rx_uart_i.fifo_i.din[5] ),
    .X(net5352));
 sg13g2_dlygate4sd3_1 hold2756 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[41] ),
    .X(net5353));
 sg13g2_dlygate4sd3_1 hold2757 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[5] ),
    .X(net5354));
 sg13g2_dlygate4sd3_1 hold2758 (.A(\soc_I.qqspi_I.spi_buf[12] ),
    .X(net5355));
 sg13g2_dlygate4sd3_1 hold2759 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[24] ),
    .X(net5356));
 sg13g2_dlygate4sd3_1 hold2760 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[51] ),
    .X(net5357));
 sg13g2_dlygate4sd3_1 hold2761 (.A(\soc_I.spi0_I.div[11] ),
    .X(net5358));
 sg13g2_dlygate4sd3_1 hold2762 (.A(\soc_I.div_reg[1] ),
    .X(net5359));
 sg13g2_dlygate4sd3_1 hold2763 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[18] ),
    .X(net5360));
 sg13g2_dlygate4sd3_1 hold2764 (.A(_00179_),
    .X(net5361));
 sg13g2_dlygate4sd3_1 hold2765 (.A(_05364_),
    .X(net5362));
 sg13g2_dlygate4sd3_1 hold2766 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[61] ),
    .X(net5363));
 sg13g2_dlygate4sd3_1 hold2767 (.A(\soc_I.spi0_I.div[15] ),
    .X(net5364));
 sg13g2_dlygate4sd3_1 hold2768 (.A(\soc_I.qqspi_I.spi_buf[10] ),
    .X(net5365));
 sg13g2_dlygate4sd3_1 hold2769 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[3] ),
    .X(net5366));
 sg13g2_dlygate4sd3_1 hold2770 (.A(\soc_I.div_reg[15] ),
    .X(net5367));
 sg13g2_dlygate4sd3_1 hold2771 (.A(\soc_I.rx_uart_i.wait_states[15] ),
    .X(net5368));
 sg13g2_dlygate4sd3_1 hold2772 (.A(_06941_),
    .X(net5369));
 sg13g2_dlygate4sd3_1 hold2773 (.A(\led[2] ),
    .X(net5370));
 sg13g2_dlygate4sd3_1 hold2774 (.A(_01457_),
    .X(net5371));
 sg13g2_dlygate4sd3_1 hold2775 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[40] ),
    .X(net5372));
 sg13g2_dlygate4sd3_1 hold2776 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[24] ),
    .X(net5373));
 sg13g2_dlygate4sd3_1 hold2777 (.A(_01225_),
    .X(net5374));
 sg13g2_dlygate4sd3_1 hold2778 (.A(\soc_I.clint_I.div[1] ),
    .X(net5375));
 sg13g2_dlygate4sd3_1 hold2779 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[6] ),
    .X(net5376));
 sg13g2_dlygate4sd3_1 hold2780 (.A(_05352_),
    .X(net5377));
 sg13g2_dlygate4sd3_1 hold2781 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[23] ),
    .X(net5378));
 sg13g2_dlygate4sd3_1 hold2782 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[42] ),
    .X(net5379));
 sg13g2_dlygate4sd3_1 hold2783 (.A(\soc_I.qqspi_I.spi_buf[14] ),
    .X(net5380));
 sg13g2_dlygate4sd3_1 hold2784 (.A(_00242_),
    .X(net5381));
 sg13g2_dlygate4sd3_1 hold2785 (.A(_01980_),
    .X(net5382));
 sg13g2_dlygate4sd3_1 hold2786 (.A(\soc_I.PC[25] ),
    .X(net5383));
 sg13g2_dlygate4sd3_1 hold2787 (.A(\soc_I.div_reg[9] ),
    .X(net5384));
 sg13g2_dlygate4sd3_1 hold2788 (.A(\soc_I.PC[13] ),
    .X(net5385));
 sg13g2_dlygate4sd3_1 hold2789 (.A(_06017_),
    .X(net5386));
 sg13g2_dlygate4sd3_1 hold2790 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[19] ),
    .X(net5387));
 sg13g2_dlygate4sd3_1 hold2791 (.A(_04697_),
    .X(net5388));
 sg13g2_dlygate4sd3_1 hold2792 (.A(\soc_I.PC[7] ),
    .X(net5389));
 sg13g2_dlygate4sd3_1 hold2793 (.A(\soc_I.clint_I.mtime[18] ),
    .X(net5390));
 sg13g2_dlygate4sd3_1 hold2794 (.A(_06337_),
    .X(net5391));
 sg13g2_dlygate4sd3_1 hold2795 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[21] ),
    .X(net5392));
 sg13g2_dlygate4sd3_1 hold2796 (.A(_01222_),
    .X(net5393));
 sg13g2_dlygate4sd3_1 hold2797 (.A(_00150_),
    .X(net5394));
 sg13g2_dlygate4sd3_1 hold2798 (.A(_01981_),
    .X(net5395));
 sg13g2_dlygate4sd3_1 hold2799 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[17] ),
    .X(net5396));
 sg13g2_dlygate4sd3_1 hold2800 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[17] ),
    .X(net5397));
 sg13g2_dlygate4sd3_1 hold2801 (.A(\soc_I.div_reg[0] ),
    .X(net5398));
 sg13g2_dlygate4sd3_1 hold2802 (.A(\soc_I.PC[15] ),
    .X(net5399));
 sg13g2_dlygate4sd3_1 hold2803 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[23] ),
    .X(net5400));
 sg13g2_dlygate4sd3_1 hold2804 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[45] ),
    .X(net5401));
 sg13g2_dlygate4sd3_1 hold2805 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[2] ),
    .X(net5402));
 sg13g2_dlygate4sd3_1 hold2806 (.A(_01203_),
    .X(net5403));
 sg13g2_dlygate4sd3_1 hold2807 (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[20] ),
    .X(net5404));
 sg13g2_dlygate4sd3_1 hold2808 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[34] ),
    .X(net5405));
 sg13g2_dlygate4sd3_1 hold2809 (.A(\soc_I.qqspi_I.spi_buf[20] ),
    .X(net5406));
 sg13g2_dlygate4sd3_1 hold2810 (.A(\soc_I.qqspi_I.spi_buf[11] ),
    .X(net5407));
 sg13g2_dlygate4sd3_1 hold2811 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[47] ),
    .X(net5408));
 sg13g2_dlygate4sd3_1 hold2812 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[29] ),
    .X(net5409));
 sg13g2_dlygate4sd3_1 hold2813 (.A(_01230_),
    .X(net5410));
 sg13g2_dlygate4sd3_1 hold2814 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[31] ),
    .X(net5411));
 sg13g2_dlygate4sd3_1 hold2815 (.A(_04731_),
    .X(net5412));
 sg13g2_dlygate4sd3_1 hold2816 (.A(\soc_I.qqspi_I.spi_buf[3] ),
    .X(net5413));
 sg13g2_dlygate4sd3_1 hold2817 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[1] ),
    .X(net5414));
 sg13g2_dlygate4sd3_1 hold2818 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[26] ),
    .X(net5415));
 sg13g2_dlygate4sd3_1 hold2819 (.A(\soc_I.clint_I.div[5] ),
    .X(net5416));
 sg13g2_dlygate4sd3_1 hold2820 (.A(\soc_I.qqspi_I.spi_buf[26] ),
    .X(net5417));
 sg13g2_dlygate4sd3_1 hold2821 (.A(_02024_),
    .X(net5418));
 sg13g2_dlygate4sd3_1 hold2822 (.A(\soc_I.qqspi_I.spi_buf[22] ),
    .X(net5419));
 sg13g2_dlygate4sd3_1 hold2823 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[21] ),
    .X(net5420));
 sg13g2_dlygate4sd3_1 hold2824 (.A(\soc_I.div_reg[4] ),
    .X(net5421));
 sg13g2_dlygate4sd3_1 hold2825 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[5] ),
    .X(net5422));
 sg13g2_dlygate4sd3_1 hold2826 (.A(_04454_),
    .X(net5423));
 sg13g2_dlygate4sd3_1 hold2827 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[38] ),
    .X(net5424));
 sg13g2_dlygate4sd3_1 hold2828 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[11] ),
    .X(net5425));
 sg13g2_dlygate4sd3_1 hold2829 (.A(\soc_I.PC[4] ),
    .X(net5426));
 sg13g2_dlygate4sd3_1 hold2830 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[29] ),
    .X(net5427));
 sg13g2_dlygate4sd3_1 hold2831 (.A(\soc_I.clint_I.mtime[16] ),
    .X(net5428));
 sg13g2_dlygate4sd3_1 hold2832 (.A(_01648_),
    .X(net5429));
 sg13g2_dlygate4sd3_1 hold2833 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[36] ),
    .X(net5430));
 sg13g2_dlygate4sd3_1 hold2834 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[32] ),
    .X(net5431));
 sg13g2_dlygate4sd3_1 hold2835 (.A(_02176_),
    .X(net5432));
 sg13g2_dlygate4sd3_1 hold2836 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[18] ),
    .X(net5433));
 sg13g2_dlygate4sd3_1 hold2837 (.A(\soc_I.div_reg[3] ),
    .X(net5434));
 sg13g2_dlygate4sd3_1 hold2838 (.A(\soc_I.qqspi_I.spi_buf[9] ),
    .X(net5435));
 sg13g2_dlygate4sd3_1 hold2839 (.A(\soc_I.div_reg[2] ),
    .X(net5436));
 sg13g2_dlygate4sd3_1 hold2840 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[14] ),
    .X(net5437));
 sg13g2_dlygate4sd3_1 hold2841 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[16] ),
    .X(net5438));
 sg13g2_dlygate4sd3_1 hold2842 (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[12] ),
    .X(net5439));
 sg13g2_dlygate4sd3_1 hold2843 (.A(_01451_),
    .X(net5440));
 sg13g2_dlygate4sd3_1 hold2844 (.A(\soc_I.PC[10] ),
    .X(net5441));
 sg13g2_dlygate4sd3_1 hold2845 (.A(\soc_I.qqspi_I.spi_buf[30] ),
    .X(net5442));
 sg13g2_dlygate4sd3_1 hold2846 (.A(_07348_),
    .X(net5443));
 sg13g2_dlygate4sd3_1 hold2847 (.A(\soc_I.clint_I.mtime[49] ),
    .X(net5444));
 sg13g2_dlygate4sd3_1 hold2848 (.A(_01682_),
    .X(net5445));
 sg13g2_dlygate4sd3_1 hold2849 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[15] ),
    .X(net5446));
 sg13g2_dlygate4sd3_1 hold2850 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[5] ),
    .X(net5447));
 sg13g2_dlygate4sd3_1 hold2851 (.A(_01206_),
    .X(net5448));
 sg13g2_dlygate4sd3_1 hold2852 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[32] ),
    .X(net5449));
 sg13g2_dlygate4sd3_1 hold2853 (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[9] ),
    .X(net5450));
 sg13g2_dlygate4sd3_1 hold2854 (.A(_01448_),
    .X(net5451));
 sg13g2_dlygate4sd3_1 hold2855 (.A(\soc_I.kianv_I.control_unit_I.main_fsm_I.mstatus[3] ),
    .X(net5452));
 sg13g2_dlygate4sd3_1 hold2856 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[41] ),
    .X(net5453));
 sg13g2_dlygate4sd3_1 hold2857 (.A(\soc_I.qqspi_I.spi_buf[29] ),
    .X(net5454));
 sg13g2_dlygate4sd3_1 hold2858 (.A(_07342_),
    .X(net5455));
 sg13g2_dlygate4sd3_1 hold2859 (.A(\soc_I.PC[12] ),
    .X(net5456));
 sg13g2_dlygate4sd3_1 hold2860 (.A(\soc_I.clint_I.div[0] ),
    .X(net5457));
 sg13g2_dlygate4sd3_1 hold2861 (.A(\soc_I.PC[28] ),
    .X(net5458));
 sg13g2_dlygate4sd3_1 hold2862 (.A(\soc_I.qqspi_I.spi_buf[2] ),
    .X(net5459));
 sg13g2_dlygate4sd3_1 hold2863 (.A(\soc_I.kianv_I.Instr[19] ),
    .X(net5460));
 sg13g2_dlygate4sd3_1 hold2864 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[44] ),
    .X(net5461));
 sg13g2_dlygate4sd3_1 hold2865 (.A(\soc_I.qqspi_I.spi_buf[23] ),
    .X(net5462));
 sg13g2_dlygate4sd3_1 hold2866 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[20] ),
    .X(net5463));
 sg13g2_dlygate4sd3_1 hold2867 (.A(_01221_),
    .X(net5464));
 sg13g2_dlygate4sd3_1 hold2868 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.exception_next_pc[10] ),
    .X(net5465));
 sg13g2_dlygate4sd3_1 hold2869 (.A(\soc_I.qqspi_I.spi_buf[0] ),
    .X(net5466));
 sg13g2_dlygate4sd3_1 hold2870 (.A(\soc_I.div_reg[5] ),
    .X(net5467));
 sg13g2_dlygate4sd3_1 hold2871 (.A(\soc_I.qqspi_I.spi_buf[1] ),
    .X(net5468));
 sg13g2_dlygate4sd3_1 hold2872 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.bit_idx[3] ),
    .X(net5469));
 sg13g2_dlygate4sd3_1 hold2873 (.A(_01371_),
    .X(net5470));
 sg13g2_dlygate4sd3_1 hold2874 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.state[0] ),
    .X(net5471));
 sg13g2_dlygate4sd3_1 hold2875 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[36] ),
    .X(net5472));
 sg13g2_dlygate4sd3_1 hold2876 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[12] ),
    .X(net5473));
 sg13g2_dlygate4sd3_1 hold2877 (.A(\soc_I.clint_I.mtime[28] ),
    .X(net5474));
 sg13g2_dlygate4sd3_1 hold2878 (.A(_06366_),
    .X(net5475));
 sg13g2_dlygate4sd3_1 hold2879 (.A(\soc_I.rx_uart_i.fifo_i.wr_ptr[2] ),
    .X(net5476));
 sg13g2_dlygate4sd3_1 hold2880 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[31] ),
    .X(net5477));
 sg13g2_dlygate4sd3_1 hold2881 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[17] ),
    .X(net5478));
 sg13g2_dlygate4sd3_1 hold2882 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[47] ),
    .X(net5479));
 sg13g2_dlygate4sd3_1 hold2883 (.A(_01184_),
    .X(net5480));
 sg13g2_dlygate4sd3_1 hold2884 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[50] ),
    .X(net5481));
 sg13g2_dlygate4sd3_1 hold2885 (.A(\soc_I.clint_I.mtime[38] ),
    .X(net5482));
 sg13g2_dlygate4sd3_1 hold2886 (.A(_01670_),
    .X(net5483));
 sg13g2_dlygate4sd3_1 hold2887 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[43] ),
    .X(net5484));
 sg13g2_dlygate4sd3_1 hold2888 (.A(\soc_I.qqspi_I.spi_buf[21] ),
    .X(net5485));
 sg13g2_dlygate4sd3_1 hold2889 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[27] ),
    .X(net5486));
 sg13g2_dlygate4sd3_1 hold2890 (.A(\soc_I.kianv_I.Instr[30] ),
    .X(net5487));
 sg13g2_dlygate4sd3_1 hold2891 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[17] ),
    .X(net5488));
 sg13g2_dlygate4sd3_1 hold2892 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[49] ),
    .X(net5489));
 sg13g2_dlygate4sd3_1 hold2893 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_state[0] ),
    .X(net5490));
 sg13g2_dlygate4sd3_1 hold2894 (.A(\soc_I.kianv_I.Instr[5] ),
    .X(net5491));
 sg13g2_dlygate4sd3_1 hold2895 (.A(\soc_I.kianv_I.Instr[26] ),
    .X(net5492));
 sg13g2_dlygate4sd3_1 hold2896 (.A(\soc_I.rx_uart_i.fifo_i.din[3] ),
    .X(net5493));
 sg13g2_dlygate4sd3_1 hold2897 (.A(\soc_I.kianv_I.Instr[4] ),
    .X(net5494));
 sg13g2_dlygate4sd3_1 hold2898 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[6] ),
    .X(net5495));
 sg13g2_dlygate4sd3_1 hold2899 (.A(_04671_),
    .X(net5496));
 sg13g2_dlygate4sd3_1 hold2900 (.A(_01143_),
    .X(net5497));
 sg13g2_dlygate4sd3_1 hold2901 (.A(\soc_I.clint_I.mtime[45] ),
    .X(net5498));
 sg13g2_dlygate4sd3_1 hold2902 (.A(_06406_),
    .X(net5499));
 sg13g2_dlygate4sd3_1 hold2903 (.A(_01677_),
    .X(net5500));
 sg13g2_dlygate4sd3_1 hold2904 (.A(\soc_I.PC[8] ),
    .X(net5501));
 sg13g2_dlygate4sd3_1 hold2905 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[11] ),
    .X(net5502));
 sg13g2_dlygate4sd3_1 hold2906 (.A(\soc_I.kianv_I.Instr[31] ),
    .X(net5503));
 sg13g2_dlygate4sd3_1 hold2907 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[26] ),
    .X(net5504));
 sg13g2_dlygate4sd3_1 hold2908 (.A(_01227_),
    .X(net5505));
 sg13g2_dlygate4sd3_1 hold2909 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[46] ),
    .X(net5506));
 sg13g2_dlygate4sd3_1 hold2910 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[51] ),
    .X(net5507));
 sg13g2_dlygate4sd3_1 hold2911 (.A(uio_out[7]),
    .X(net5508));
 sg13g2_dlygate4sd3_1 hold2912 (.A(\soc_I.clint_I.mtime[31] ),
    .X(net5509));
 sg13g2_dlygate4sd3_1 hold2913 (.A(_06378_),
    .X(net5510));
 sg13g2_dlygate4sd3_1 hold2914 (.A(\soc_I.clint_I.mtime[22] ),
    .X(net5511));
 sg13g2_dlygate4sd3_1 hold2915 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[27] ),
    .X(net5512));
 sg13g2_dlygate4sd3_1 hold2916 (.A(uio_out[6]),
    .X(net5513));
 sg13g2_dlygate4sd3_1 hold2917 (.A(_01982_),
    .X(net5514));
 sg13g2_dlygate4sd3_1 hold2918 (.A(\soc_I.clint_I.mtime[2] ),
    .X(net5515));
 sg13g2_dlygate4sd3_1 hold2919 (.A(_01634_),
    .X(net5516));
 sg13g2_dlygate4sd3_1 hold2920 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mtvec[24] ),
    .X(net5517));
 sg13g2_dlygate4sd3_1 hold2921 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.bit_idx[2] ),
    .X(net5518));
 sg13g2_dlygate4sd3_1 hold2922 (.A(_01370_),
    .X(net5519));
 sg13g2_dlygate4sd3_1 hold2923 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[13] ),
    .X(net5520));
 sg13g2_dlygate4sd3_1 hold2924 (.A(\soc_I.rx_uart_i.data_rd ),
    .X(net5521));
 sg13g2_dlygate4sd3_1 hold2925 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mepc[21] ),
    .X(net5522));
 sg13g2_dlygate4sd3_1 hold2926 (.A(\soc_I.kianv_I.Instr[6] ),
    .X(net5523));
 sg13g2_dlygate4sd3_1 hold2927 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[20] ),
    .X(net5524));
 sg13g2_dlygate4sd3_1 hold2928 (.A(_04699_),
    .X(net5525));
 sg13g2_dlygate4sd3_1 hold2929 (.A(\soc_I.kianv_I.Instr[14] ),
    .X(net5526));
 sg13g2_dlygate4sd3_1 hold2930 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[39] ),
    .X(net5527));
 sg13g2_dlygate4sd3_1 hold2931 (.A(\soc_I.rx_uart_i.fifo_i.din[7] ),
    .X(net5528));
 sg13g2_dlygate4sd3_1 hold2932 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[24] ),
    .X(net5529));
 sg13g2_dlygate4sd3_1 hold2933 (.A(\soc_I.qqspi_I.spi_buf[28] ),
    .X(net5530));
 sg13g2_dlygate4sd3_1 hold2934 (.A(_02026_),
    .X(net5531));
 sg13g2_dlygate4sd3_1 hold2935 (.A(\soc_I.clint_I.mtime[61] ),
    .X(net5532));
 sg13g2_dlygate4sd3_1 hold2936 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[35] ),
    .X(net5533));
 sg13g2_dlygate4sd3_1 hold2937 (.A(_00291_),
    .X(net5534));
 sg13g2_dlygate4sd3_1 hold2938 (.A(_01979_),
    .X(net5535));
 sg13g2_dlygate4sd3_1 hold2939 (.A(\soc_I.clint_I.mtime[34] ),
    .X(net5536));
 sg13g2_dlygate4sd3_1 hold2940 (.A(_06386_),
    .X(net5537));
 sg13g2_dlygate4sd3_1 hold2941 (.A(_01667_),
    .X(net5538));
 sg13g2_dlygate4sd3_1 hold2942 (.A(\soc_I.kianv_I.Instr[9] ),
    .X(net5539));
 sg13g2_dlygate4sd3_1 hold2943 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[5] ),
    .X(net5540));
 sg13g2_dlygate4sd3_1 hold2944 (.A(\soc_I.kianv_I.datapath_unit_I.OldPC[13] ),
    .X(net5541));
 sg13g2_dlygate4sd3_1 hold2945 (.A(\soc_I.kianv_I.Instr[2] ),
    .X(net5542));
 sg13g2_dlygate4sd3_1 hold2946 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[13] ),
    .X(net5543));
 sg13g2_dlygate4sd3_1 hold2947 (.A(\soc_I.kianv_I.Instr[28] ),
    .X(net5544));
 sg13g2_dlygate4sd3_1 hold2948 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[26] ),
    .X(net5545));
 sg13g2_dlygate4sd3_1 hold2949 (.A(\soc_I.clint_I.mtime[36] ),
    .X(net5546));
 sg13g2_dlygate4sd3_1 hold2950 (.A(_01668_),
    .X(net5547));
 sg13g2_dlygate4sd3_1 hold2951 (.A(\soc_I.kianv_I.Instr[13] ),
    .X(net5548));
 sg13g2_dlygate4sd3_1 hold2952 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[53] ),
    .X(net5549));
 sg13g2_dlygate4sd3_1 hold2953 (.A(\soc_I.spi0_I.div[0] ),
    .X(net5550));
 sg13g2_dlygate4sd3_1 hold2954 (.A(\soc_I.kianv_I.Instr[25] ),
    .X(net5551));
 sg13g2_dlygate4sd3_1 hold2955 (.A(\soc_I.clint_I.mtime[46] ),
    .X(net5552));
 sg13g2_dlygate4sd3_1 hold2956 (.A(_01678_),
    .X(net5553));
 sg13g2_dlygate4sd3_1 hold2957 (.A(\soc_I.kianv_I.datapath_unit_I.mul_I.rslt[33] ),
    .X(net5554));
 sg13g2_dlygate4sd3_1 hold2958 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[33] ),
    .X(net5555));
 sg13g2_dlygate4sd3_1 hold2959 (.A(\soc_I.kianv_I.Instr[8] ),
    .X(net5556));
 sg13g2_dlygate4sd3_1 hold2960 (.A(\soc_I.kianv_I.Instr[7] ),
    .X(net5557));
 sg13g2_dlygate4sd3_1 hold2961 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.instr_cnt_I.q[25] ),
    .X(net5558));
 sg13g2_dlygate4sd3_1 hold2962 (.A(\soc_I.kianv_I.Instr[11] ),
    .X(net5559));
 sg13g2_dlygate4sd3_1 hold2963 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[0] ),
    .X(net5560));
 sg13g2_dlygate4sd3_1 hold2964 (.A(\soc_I.spi_div_ready ),
    .X(net5561));
 sg13g2_dlygate4sd3_1 hold2965 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[31] ),
    .X(net5562));
 sg13g2_dlygate4sd3_1 hold2966 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][19] ),
    .X(net5563));
 sg13g2_dlygate4sd3_1 hold2967 (.A(\soc_I.kianv_I.Instr[12] ),
    .X(net5564));
 sg13g2_dlygate4sd3_1 hold2968 (.A(\soc_I.kianv_I.datapath_unit_I.AMOTmpData_I.q[0] ),
    .X(net5565));
 sg13g2_dlygate4sd3_1 hold2969 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[26] ),
    .X(net5566));
 sg13g2_dlygate4sd3_1 hold2970 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[13] ),
    .X(net5567));
 sg13g2_dlygate4sd3_1 hold2971 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.rem_rslt[31] ),
    .X(net5568));
 sg13g2_dlygate4sd3_1 hold2972 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[39] ),
    .X(net5569));
 sg13g2_dlygate4sd3_1 hold2973 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.cycle_cnt_I.q[59] ),
    .X(net5570));
 sg13g2_dlygate4sd3_1 hold2974 (.A(\soc_I.clint_I.tick_cnt[9] ),
    .X(net5571));
 sg13g2_dlygate4sd3_1 hold2975 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[16] ),
    .X(net5572));
 sg13g2_dlygate4sd3_1 hold2976 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[14] ),
    .X(net5573));
 sg13g2_dlygate4sd3_1 hold2977 (.A(\soc_I.rx_uart_i.fifo_i.cnt[2] ),
    .X(net5574));
 sg13g2_dlygate4sd3_1 hold2978 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][28] ),
    .X(net5575));
 sg13g2_dlygate4sd3_1 hold2979 (.A(_03635_),
    .X(net5576));
 sg13g2_dlygate4sd3_1 hold2980 (.A(\soc_I.kianv_I.datapath_unit_I.csr_exception_handler_I.mscratch[0] ),
    .X(net5577));
 sg13g2_dlygate4sd3_1 hold2981 (.A(\soc_I.qqspi_I.spi_buf[28] ),
    .X(net5578));
 sg13g2_dlygate4sd3_1 hold2982 (.A(\soc_I.kianv_I.datapath_unit_I.register_file_I.bank0[9][29] ),
    .X(net5579));
 sg13g2_dlygate4sd3_1 hold2983 (.A(\soc_I.kianv_I.datapath_unit_I.div_I.div_rslt[14] ),
    .X(net5580));
 sg13g2_antennanp ANTENNA_1 (.A(_00187_));
 sg13g2_antennanp ANTENNA_2 (.A(_00187_));
 sg13g2_antennanp ANTENNA_3 (.A(_00187_));
 sg13g2_antennanp ANTENNA_4 (.A(_00187_));
 sg13g2_antennanp ANTENNA_5 (.A(_00225_));
 sg13g2_antennanp ANTENNA_6 (.A(_00229_));
 sg13g2_antennanp ANTENNA_7 (.A(_00230_));
 sg13g2_antennanp ANTENNA_8 (.A(_00231_));
 sg13g2_antennanp ANTENNA_9 (.A(_00232_));
 sg13g2_antennanp ANTENNA_10 (.A(_00233_));
 sg13g2_antennanp ANTENNA_11 (.A(_00235_));
 sg13g2_antennanp ANTENNA_12 (.A(_00292_));
 sg13g2_antennanp ANTENNA_13 (.A(_00292_));
 sg13g2_antennanp ANTENNA_14 (.A(_00292_));
 sg13g2_antennanp ANTENNA_15 (.A(_00292_));
 sg13g2_antennanp ANTENNA_16 (.A(_00292_));
 sg13g2_antennanp ANTENNA_17 (.A(_00292_));
 sg13g2_antennanp ANTENNA_18 (.A(_00742_));
 sg13g2_antennanp ANTENNA_19 (.A(_00743_));
 sg13g2_antennanp ANTENNA_20 (.A(_00751_));
 sg13g2_antennanp ANTENNA_21 (.A(_00752_));
 sg13g2_antennanp ANTENNA_22 (.A(_00758_));
 sg13g2_antennanp ANTENNA_23 (.A(_00758_));
 sg13g2_antennanp ANTENNA_24 (.A(_00762_));
 sg13g2_antennanp ANTENNA_25 (.A(_00772_));
 sg13g2_antennanp ANTENNA_26 (.A(_01001_));
 sg13g2_antennanp ANTENNA_27 (.A(_01002_));
 sg13g2_antennanp ANTENNA_28 (.A(_02684_));
 sg13g2_antennanp ANTENNA_29 (.A(_02691_));
 sg13g2_antennanp ANTENNA_30 (.A(_02698_));
 sg13g2_antennanp ANTENNA_31 (.A(_02701_));
 sg13g2_antennanp ANTENNA_32 (.A(_02707_));
 sg13g2_antennanp ANTENNA_33 (.A(_02708_));
 sg13g2_antennanp ANTENNA_34 (.A(_02902_));
 sg13g2_antennanp ANTENNA_35 (.A(_03370_));
 sg13g2_antennanp ANTENNA_36 (.A(_10388_));
 sg13g2_antennanp ANTENNA_37 (.A(_10856_));
 sg13g2_antennanp ANTENNA_38 (.A(_10856_));
 sg13g2_antennanp ANTENNA_39 (.A(_10856_));
 sg13g2_antennanp ANTENNA_40 (.A(_10856_));
 sg13g2_antennanp ANTENNA_41 (.A(_10856_));
 sg13g2_antennanp ANTENNA_42 (.A(_10856_));
 sg13g2_antennanp ANTENNA_43 (.A(_10856_));
 sg13g2_antennanp ANTENNA_44 (.A(_10856_));
 sg13g2_antennanp ANTENNA_45 (.A(_10856_));
 sg13g2_antennanp ANTENNA_46 (.A(_10856_));
 sg13g2_antennanp ANTENNA_47 (.A(_10856_));
 sg13g2_antennanp ANTENNA_48 (.A(_10856_));
 sg13g2_antennanp ANTENNA_49 (.A(_10856_));
 sg13g2_antennanp ANTENNA_50 (.A(_10856_));
 sg13g2_antennanp ANTENNA_51 (.A(_10856_));
 sg13g2_antennanp ANTENNA_52 (.A(_10856_));
 sg13g2_antennanp ANTENNA_53 (.A(_10856_));
 sg13g2_antennanp ANTENNA_54 (.A(_10856_));
 sg13g2_antennanp ANTENNA_55 (.A(_12499_));
 sg13g2_antennanp ANTENNA_56 (.A(_12499_));
 sg13g2_antennanp ANTENNA_57 (.A(_12499_));
 sg13g2_antennanp ANTENNA_58 (.A(_12499_));
 sg13g2_antennanp ANTENNA_59 (.A(_12787_));
 sg13g2_antennanp ANTENNA_60 (.A(_12795_));
 sg13g2_antennanp ANTENNA_61 (.A(_12893_));
 sg13g2_antennanp ANTENNA_62 (.A(_12893_));
 sg13g2_antennanp ANTENNA_63 (.A(_12893_));
 sg13g2_antennanp ANTENNA_64 (.A(_12893_));
 sg13g2_antennanp ANTENNA_65 (.A(_13330_));
 sg13g2_antennanp ANTENNA_66 (.A(_13330_));
 sg13g2_antennanp ANTENNA_67 (.A(_13330_));
 sg13g2_antennanp ANTENNA_68 (.A(_13330_));
 sg13g2_antennanp ANTENNA_69 (.A(_13836_));
 sg13g2_antennanp ANTENNA_70 (.A(_13836_));
 sg13g2_antennanp ANTENNA_71 (.A(_13836_));
 sg13g2_antennanp ANTENNA_72 (.A(_13836_));
 sg13g2_antennanp ANTENNA_73 (.A(_13974_));
 sg13g2_antennanp ANTENNA_74 (.A(_13974_));
 sg13g2_antennanp ANTENNA_75 (.A(_13984_));
 sg13g2_antennanp ANTENNA_76 (.A(_13984_));
 sg13g2_antennanp ANTENNA_77 (.A(_14046_));
 sg13g2_antennanp ANTENNA_78 (.A(_14046_));
 sg13g2_antennanp ANTENNA_79 (.A(_14046_));
 sg13g2_antennanp ANTENNA_80 (.A(_14046_));
 sg13g2_antennanp ANTENNA_81 (.A(_14046_));
 sg13g2_antennanp ANTENNA_82 (.A(_14046_));
 sg13g2_antennanp ANTENNA_83 (.A(_14046_));
 sg13g2_antennanp ANTENNA_84 (.A(_14046_));
 sg13g2_antennanp ANTENNA_85 (.A(_14046_));
 sg13g2_antennanp ANTENNA_86 (.A(_14046_));
 sg13g2_antennanp ANTENNA_87 (.A(_14046_));
 sg13g2_antennanp ANTENNA_88 (.A(_14059_));
 sg13g2_antennanp ANTENNA_89 (.A(_14065_));
 sg13g2_antennanp ANTENNA_90 (.A(_14065_));
 sg13g2_antennanp ANTENNA_91 (.A(_14065_));
 sg13g2_antennanp ANTENNA_92 (.A(_14065_));
 sg13g2_antennanp ANTENNA_93 (.A(_14065_));
 sg13g2_antennanp ANTENNA_94 (.A(_14065_));
 sg13g2_antennanp ANTENNA_95 (.A(_14065_));
 sg13g2_antennanp ANTENNA_96 (.A(_14065_));
 sg13g2_antennanp ANTENNA_97 (.A(_14080_));
 sg13g2_antennanp ANTENNA_98 (.A(_14086_));
 sg13g2_antennanp ANTENNA_99 (.A(_14090_));
 sg13g2_antennanp ANTENNA_100 (.A(_14097_));
 sg13g2_antennanp ANTENNA_101 (.A(_14109_));
 sg13g2_antennanp ANTENNA_102 (.A(clk));
 sg13g2_antennanp ANTENNA_103 (.A(clk));
 sg13g2_antennanp ANTENNA_104 (.A(\soc_I.clint_I.addr[1] ));
 sg13g2_antennanp ANTENNA_105 (.A(\soc_I.clint_I.addr[1] ));
 sg13g2_antennanp ANTENNA_106 (.A(\soc_I.clint_I.addr[1] ));
 sg13g2_antennanp ANTENNA_107 (.A(\soc_I.clint_I.addr[1] ));
 sg13g2_antennanp ANTENNA_108 (.A(\soc_I.clint_I.addr[1] ));
 sg13g2_antennanp ANTENNA_109 (.A(\soc_I.clint_I.addr[1] ));
 sg13g2_antennanp ANTENNA_110 (.A(\soc_I.clint_I.addr[1] ));
 sg13g2_antennanp ANTENNA_111 (.A(\soc_I.kianv_I.datapath_unit_I.A1[13] ));
 sg13g2_antennanp ANTENNA_112 (.A(\soc_I.kianv_I.datapath_unit_I.A1[20] ));
 sg13g2_antennanp ANTENNA_113 (.A(\soc_I.kianv_I.datapath_unit_I.A1[22] ));
 sg13g2_antennanp ANTENNA_114 (.A(\soc_I.kianv_I.datapath_unit_I.A1[26] ));
 sg13g2_antennanp ANTENNA_115 (.A(\soc_I.kianv_I.datapath_unit_I.A1[3] ));
 sg13g2_antennanp ANTENNA_116 (.A(\soc_I.kianv_I.datapath_unit_I.A1[4] ));
 sg13g2_antennanp ANTENNA_117 (.A(\soc_I.kianv_I.datapath_unit_I.A1[9] ));
 sg13g2_antennanp ANTENNA_118 (.A(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[13] ));
 sg13g2_antennanp ANTENNA_119 (.A(\soc_I.kianv_I.datapath_unit_I.Data[13] ));
 sg13g2_antennanp ANTENNA_120 (.A(\soc_I.kianv_I.datapath_unit_I.Data[13] ));
 sg13g2_antennanp ANTENNA_121 (.A(\soc_I.kianv_I.datapath_unit_I.Data[8] ));
 sg13g2_antennanp ANTENNA_122 (.A(\soc_I.kianv_I.datapath_unit_I.Data[8] ));
 sg13g2_antennanp ANTENNA_123 (.A(\soc_I.kianv_I.datapath_unit_I.MULExtResult[16] ));
 sg13g2_antennanp ANTENNA_124 (.A(uio_oe[1]));
 sg13g2_antennanp ANTENNA_125 (.A(uio_oe[1]));
 sg13g2_antennanp ANTENNA_126 (.A(uio_out[0]));
 sg13g2_antennanp ANTENNA_127 (.A(uio_out[0]));
 sg13g2_antennanp ANTENNA_128 (.A(uio_out[6]));
 sg13g2_antennanp ANTENNA_129 (.A(uio_out[6]));
 sg13g2_antennanp ANTENNA_130 (.A(uio_out[7]));
 sg13g2_antennanp ANTENNA_131 (.A(uio_out[7]));
 sg13g2_antennanp ANTENNA_132 (.A(net7490));
 sg13g2_antennanp ANTENNA_133 (.A(net7490));
 sg13g2_antennanp ANTENNA_134 (.A(net7490));
 sg13g2_antennanp ANTENNA_135 (.A(net7490));
 sg13g2_antennanp ANTENNA_136 (.A(net7510));
 sg13g2_antennanp ANTENNA_137 (.A(net7510));
 sg13g2_antennanp ANTENNA_138 (.A(net7510));
 sg13g2_antennanp ANTENNA_139 (.A(net7510));
 sg13g2_antennanp ANTENNA_140 (.A(net7533));
 sg13g2_antennanp ANTENNA_141 (.A(net7533));
 sg13g2_antennanp ANTENNA_142 (.A(net7533));
 sg13g2_antennanp ANTENNA_143 (.A(net7533));
 sg13g2_antennanp ANTENNA_144 (.A(net7533));
 sg13g2_antennanp ANTENNA_145 (.A(net7533));
 sg13g2_antennanp ANTENNA_146 (.A(net7533));
 sg13g2_antennanp ANTENNA_147 (.A(net7533));
 sg13g2_antennanp ANTENNA_148 (.A(net7533));
 sg13g2_antennanp ANTENNA_149 (.A(net7618));
 sg13g2_antennanp ANTENNA_150 (.A(net7618));
 sg13g2_antennanp ANTENNA_151 (.A(net7618));
 sg13g2_antennanp ANTENNA_152 (.A(net7618));
 sg13g2_antennanp ANTENNA_153 (.A(net7618));
 sg13g2_antennanp ANTENNA_154 (.A(net7618));
 sg13g2_antennanp ANTENNA_155 (.A(net7618));
 sg13g2_antennanp ANTENNA_156 (.A(net7618));
 sg13g2_antennanp ANTENNA_157 (.A(net7618));
 sg13g2_antennanp ANTENNA_158 (.A(net7618));
 sg13g2_antennanp ANTENNA_159 (.A(net7618));
 sg13g2_antennanp ANTENNA_160 (.A(net7618));
 sg13g2_antennanp ANTENNA_161 (.A(net7618));
 sg13g2_antennanp ANTENNA_162 (.A(net7618));
 sg13g2_antennanp ANTENNA_163 (.A(net7618));
 sg13g2_antennanp ANTENNA_164 (.A(net7618));
 sg13g2_antennanp ANTENNA_165 (.A(net7618));
 sg13g2_antennanp ANTENNA_166 (.A(net7618));
 sg13g2_antennanp ANTENNA_167 (.A(net7618));
 sg13g2_antennanp ANTENNA_168 (.A(net7618));
 sg13g2_antennanp ANTENNA_169 (.A(net7618));
 sg13g2_antennanp ANTENNA_170 (.A(net7647));
 sg13g2_antennanp ANTENNA_171 (.A(net7647));
 sg13g2_antennanp ANTENNA_172 (.A(net7647));
 sg13g2_antennanp ANTENNA_173 (.A(net7647));
 sg13g2_antennanp ANTENNA_174 (.A(net7647));
 sg13g2_antennanp ANTENNA_175 (.A(net7647));
 sg13g2_antennanp ANTENNA_176 (.A(net7647));
 sg13g2_antennanp ANTENNA_177 (.A(net7668));
 sg13g2_antennanp ANTENNA_178 (.A(net7668));
 sg13g2_antennanp ANTENNA_179 (.A(net7668));
 sg13g2_antennanp ANTENNA_180 (.A(net7668));
 sg13g2_antennanp ANTENNA_181 (.A(net8597));
 sg13g2_antennanp ANTENNA_182 (.A(net8597));
 sg13g2_antennanp ANTENNA_183 (.A(net8597));
 sg13g2_antennanp ANTENNA_184 (.A(net8597));
 sg13g2_antennanp ANTENNA_185 (.A(net8597));
 sg13g2_antennanp ANTENNA_186 (.A(net8597));
 sg13g2_antennanp ANTENNA_187 (.A(net8597));
 sg13g2_antennanp ANTENNA_188 (.A(net8597));
 sg13g2_antennanp ANTENNA_189 (.A(net8597));
 sg13g2_antennanp ANTENNA_190 (.A(net8597));
 sg13g2_antennanp ANTENNA_191 (.A(net8597));
 sg13g2_antennanp ANTENNA_192 (.A(net8597));
 sg13g2_antennanp ANTENNA_193 (.A(net8597));
 sg13g2_antennanp ANTENNA_194 (.A(net8674));
 sg13g2_antennanp ANTENNA_195 (.A(net8674));
 sg13g2_antennanp ANTENNA_196 (.A(net8674));
 sg13g2_antennanp ANTENNA_197 (.A(net8674));
 sg13g2_antennanp ANTENNA_198 (.A(net8674));
 sg13g2_antennanp ANTENNA_199 (.A(net8674));
 sg13g2_antennanp ANTENNA_200 (.A(net8674));
 sg13g2_antennanp ANTENNA_201 (.A(net8674));
 sg13g2_antennanp ANTENNA_202 (.A(net8922));
 sg13g2_antennanp ANTENNA_203 (.A(net8922));
 sg13g2_antennanp ANTENNA_204 (.A(net8922));
 sg13g2_antennanp ANTENNA_205 (.A(net8922));
 sg13g2_antennanp ANTENNA_206 (.A(net8922));
 sg13g2_antennanp ANTENNA_207 (.A(net8922));
 sg13g2_antennanp ANTENNA_208 (.A(net8922));
 sg13g2_antennanp ANTENNA_209 (.A(net8922));
 sg13g2_antennanp ANTENNA_210 (.A(net8962));
 sg13g2_antennanp ANTENNA_211 (.A(net8962));
 sg13g2_antennanp ANTENNA_212 (.A(net8962));
 sg13g2_antennanp ANTENNA_213 (.A(net8962));
 sg13g2_antennanp ANTENNA_214 (.A(net8962));
 sg13g2_antennanp ANTENNA_215 (.A(net8962));
 sg13g2_antennanp ANTENNA_216 (.A(net8962));
 sg13g2_antennanp ANTENNA_217 (.A(net8962));
 sg13g2_antennanp ANTENNA_218 (.A(net8962));
 sg13g2_antennanp ANTENNA_219 (.A(net8962));
 sg13g2_antennanp ANTENNA_220 (.A(net8962));
 sg13g2_antennanp ANTENNA_221 (.A(net8962));
 sg13g2_antennanp ANTENNA_222 (.A(net8962));
 sg13g2_antennanp ANTENNA_223 (.A(net8962));
 sg13g2_antennanp ANTENNA_224 (.A(net9110));
 sg13g2_antennanp ANTENNA_225 (.A(net9110));
 sg13g2_antennanp ANTENNA_226 (.A(net9110));
 sg13g2_antennanp ANTENNA_227 (.A(net9110));
 sg13g2_antennanp ANTENNA_228 (.A(net9110));
 sg13g2_antennanp ANTENNA_229 (.A(net9110));
 sg13g2_antennanp ANTENNA_230 (.A(net9110));
 sg13g2_antennanp ANTENNA_231 (.A(net9110));
 sg13g2_antennanp ANTENNA_232 (.A(net9110));
 sg13g2_antennanp ANTENNA_233 (.A(net9110));
 sg13g2_antennanp ANTENNA_234 (.A(net9110));
 sg13g2_antennanp ANTENNA_235 (.A(net9110));
 sg13g2_antennanp ANTENNA_236 (.A(net9110));
 sg13g2_antennanp ANTENNA_237 (.A(net9110));
 sg13g2_antennanp ANTENNA_238 (.A(net9110));
 sg13g2_antennanp ANTENNA_239 (.A(net9110));
 sg13g2_antennanp ANTENNA_240 (.A(net9110));
 sg13g2_antennanp ANTENNA_241 (.A(net9110));
 sg13g2_antennanp ANTENNA_242 (.A(net9110));
 sg13g2_antennanp ANTENNA_243 (.A(net9110));
 sg13g2_antennanp ANTENNA_244 (.A(net9439));
 sg13g2_antennanp ANTENNA_245 (.A(net9439));
 sg13g2_antennanp ANTENNA_246 (.A(net9439));
 sg13g2_antennanp ANTENNA_247 (.A(net9439));
 sg13g2_antennanp ANTENNA_248 (.A(net9439));
 sg13g2_antennanp ANTENNA_249 (.A(net9439));
 sg13g2_antennanp ANTENNA_250 (.A(net9439));
 sg13g2_antennanp ANTENNA_251 (.A(net9439));
 sg13g2_antennanp ANTENNA_252 (.A(net9439));
 sg13g2_antennanp ANTENNA_253 (.A(net9545));
 sg13g2_antennanp ANTENNA_254 (.A(net9545));
 sg13g2_antennanp ANTENNA_255 (.A(net9545));
 sg13g2_antennanp ANTENNA_256 (.A(net9545));
 sg13g2_antennanp ANTENNA_257 (.A(net10));
 sg13g2_antennanp ANTENNA_258 (.A(net13));
 sg13g2_antennanp ANTENNA_259 (.A(net13));
 sg13g2_antennanp ANTENNA_260 (.A(net13));
 sg13g2_antennanp ANTENNA_261 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_262 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_263 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_264 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_265 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_266 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_267 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_268 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_269 (.A(clknet_2_2_0_clk));
 sg13g2_antennanp ANTENNA_270 (.A(clknet_2_2_0_clk));
 sg13g2_antennanp ANTENNA_271 (.A(clknet_2_2_0_clk));
 sg13g2_antennanp ANTENNA_272 (.A(clknet_2_2_0_clk));
 sg13g2_antennanp ANTENNA_273 (.A(clknet_2_2_0_clk));
 sg13g2_antennanp ANTENNA_274 (.A(clknet_2_2_0_clk));
 sg13g2_antennanp ANTENNA_275 (.A(clknet_2_2_0_clk));
 sg13g2_antennanp ANTENNA_276 (.A(clknet_2_2_0_clk));
 sg13g2_antennanp ANTENNA_277 (.A(clknet_2_2_0_clk));
 sg13g2_antennanp ANTENNA_278 (.A(clknet_2_2_0_clk));
 sg13g2_antennanp ANTENNA_279 (.A(clknet_2_2_0_clk));
 sg13g2_antennanp ANTENNA_280 (.A(clknet_2_2_0_clk));
 sg13g2_antennanp ANTENNA_281 (.A(clknet_2_2_0_clk));
 sg13g2_antennanp ANTENNA_282 (.A(clknet_2_2_0_clk));
 sg13g2_antennanp ANTENNA_283 (.A(clknet_2_2_0_clk));
 sg13g2_antennanp ANTENNA_284 (.A(clknet_2_2_0_clk));
 sg13g2_antennanp ANTENNA_285 (.A(clknet_2_2_0_clk));
 sg13g2_antennanp ANTENNA_286 (.A(clknet_2_2_0_clk));
 sg13g2_antennanp ANTENNA_287 (.A(clknet_2_2_0_clk));
 sg13g2_antennanp ANTENNA_288 (.A(clknet_2_2_0_clk));
 sg13g2_antennanp ANTENNA_289 (.A(net5385));
 sg13g2_antennanp ANTENNA_290 (.A(_00187_));
 sg13g2_antennanp ANTENNA_291 (.A(_00187_));
 sg13g2_antennanp ANTENNA_292 (.A(_00187_));
 sg13g2_antennanp ANTENNA_293 (.A(_00187_));
 sg13g2_antennanp ANTENNA_294 (.A(_00225_));
 sg13g2_antennanp ANTENNA_295 (.A(_00229_));
 sg13g2_antennanp ANTENNA_296 (.A(_00230_));
 sg13g2_antennanp ANTENNA_297 (.A(_00231_));
 sg13g2_antennanp ANTENNA_298 (.A(_00232_));
 sg13g2_antennanp ANTENNA_299 (.A(_00233_));
 sg13g2_antennanp ANTENNA_300 (.A(_00235_));
 sg13g2_antennanp ANTENNA_301 (.A(_00742_));
 sg13g2_antennanp ANTENNA_302 (.A(_00743_));
 sg13g2_antennanp ANTENNA_303 (.A(_00750_));
 sg13g2_antennanp ANTENNA_304 (.A(_00751_));
 sg13g2_antennanp ANTENNA_305 (.A(_00752_));
 sg13g2_antennanp ANTENNA_306 (.A(_00754_));
 sg13g2_antennanp ANTENNA_307 (.A(_01001_));
 sg13g2_antennanp ANTENNA_308 (.A(_01002_));
 sg13g2_antennanp ANTENNA_309 (.A(_02689_));
 sg13g2_antennanp ANTENNA_310 (.A(_02690_));
 sg13g2_antennanp ANTENNA_311 (.A(_02698_));
 sg13g2_antennanp ANTENNA_312 (.A(_02707_));
 sg13g2_antennanp ANTENNA_313 (.A(_02708_));
 sg13g2_antennanp ANTENNA_314 (.A(_02710_));
 sg13g2_antennanp ANTENNA_315 (.A(_02902_));
 sg13g2_antennanp ANTENNA_316 (.A(_03370_));
 sg13g2_antennanp ANTENNA_317 (.A(_12499_));
 sg13g2_antennanp ANTENNA_318 (.A(_12499_));
 sg13g2_antennanp ANTENNA_319 (.A(_12499_));
 sg13g2_antennanp ANTENNA_320 (.A(_12499_));
 sg13g2_antennanp ANTENNA_321 (.A(_12787_));
 sg13g2_antennanp ANTENNA_322 (.A(_12795_));
 sg13g2_antennanp ANTENNA_323 (.A(_12893_));
 sg13g2_antennanp ANTENNA_324 (.A(_12893_));
 sg13g2_antennanp ANTENNA_325 (.A(_12893_));
 sg13g2_antennanp ANTENNA_326 (.A(_12893_));
 sg13g2_antennanp ANTENNA_327 (.A(_13836_));
 sg13g2_antennanp ANTENNA_328 (.A(_13836_));
 sg13g2_antennanp ANTENNA_329 (.A(_13836_));
 sg13g2_antennanp ANTENNA_330 (.A(_13836_));
 sg13g2_antennanp ANTENNA_331 (.A(_13974_));
 sg13g2_antennanp ANTENNA_332 (.A(_13974_));
 sg13g2_antennanp ANTENNA_333 (.A(_13974_));
 sg13g2_antennanp ANTENNA_334 (.A(_13974_));
 sg13g2_antennanp ANTENNA_335 (.A(_13984_));
 sg13g2_antennanp ANTENNA_336 (.A(_13984_));
 sg13g2_antennanp ANTENNA_337 (.A(_14059_));
 sg13g2_antennanp ANTENNA_338 (.A(_14065_));
 sg13g2_antennanp ANTENNA_339 (.A(_14065_));
 sg13g2_antennanp ANTENNA_340 (.A(_14065_));
 sg13g2_antennanp ANTENNA_341 (.A(_14065_));
 sg13g2_antennanp ANTENNA_342 (.A(_14065_));
 sg13g2_antennanp ANTENNA_343 (.A(_14065_));
 sg13g2_antennanp ANTENNA_344 (.A(_14080_));
 sg13g2_antennanp ANTENNA_345 (.A(_14086_));
 sg13g2_antennanp ANTENNA_346 (.A(_14090_));
 sg13g2_antennanp ANTENNA_347 (.A(_14097_));
 sg13g2_antennanp ANTENNA_348 (.A(_14109_));
 sg13g2_antennanp ANTENNA_349 (.A(clk));
 sg13g2_antennanp ANTENNA_350 (.A(clk));
 sg13g2_antennanp ANTENNA_351 (.A(\soc_I.PC[6] ));
 sg13g2_antennanp ANTENNA_352 (.A(\soc_I.PC[6] ));
 sg13g2_antennanp ANTENNA_353 (.A(\soc_I.PC[6] ));
 sg13g2_antennanp ANTENNA_354 (.A(\soc_I.PC[6] ));
 sg13g2_antennanp ANTENNA_355 (.A(\soc_I.clint_I.addr[1] ));
 sg13g2_antennanp ANTENNA_356 (.A(\soc_I.clint_I.addr[1] ));
 sg13g2_antennanp ANTENNA_357 (.A(\soc_I.clint_I.addr[1] ));
 sg13g2_antennanp ANTENNA_358 (.A(\soc_I.clint_I.addr[1] ));
 sg13g2_antennanp ANTENNA_359 (.A(\soc_I.clint_I.addr[1] ));
 sg13g2_antennanp ANTENNA_360 (.A(\soc_I.clint_I.addr[1] ));
 sg13g2_antennanp ANTENNA_361 (.A(\soc_I.clint_I.addr[1] ));
 sg13g2_antennanp ANTENNA_362 (.A(\soc_I.clint_I.addr[1] ));
 sg13g2_antennanp ANTENNA_363 (.A(\soc_I.clint_I.addr[1] ));
 sg13g2_antennanp ANTENNA_364 (.A(\soc_I.kianv_I.datapath_unit_I.A1[13] ));
 sg13g2_antennanp ANTENNA_365 (.A(\soc_I.kianv_I.datapath_unit_I.A1[20] ));
 sg13g2_antennanp ANTENNA_366 (.A(\soc_I.kianv_I.datapath_unit_I.A1[22] ));
 sg13g2_antennanp ANTENNA_367 (.A(\soc_I.kianv_I.datapath_unit_I.A1[26] ));
 sg13g2_antennanp ANTENNA_368 (.A(\soc_I.kianv_I.datapath_unit_I.A1[3] ));
 sg13g2_antennanp ANTENNA_369 (.A(\soc_I.kianv_I.datapath_unit_I.A1[4] ));
 sg13g2_antennanp ANTENNA_370 (.A(\soc_I.kianv_I.datapath_unit_I.A1[9] ));
 sg13g2_antennanp ANTENNA_371 (.A(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[13] ));
 sg13g2_antennanp ANTENNA_372 (.A(\soc_I.kianv_I.datapath_unit_I.Data[4] ));
 sg13g2_antennanp ANTENNA_373 (.A(\soc_I.kianv_I.datapath_unit_I.Data[4] ));
 sg13g2_antennanp ANTENNA_374 (.A(\soc_I.kianv_I.datapath_unit_I.Data[4] ));
 sg13g2_antennanp ANTENNA_375 (.A(\soc_I.kianv_I.datapath_unit_I.Data[4] ));
 sg13g2_antennanp ANTENNA_376 (.A(\soc_I.kianv_I.datapath_unit_I.Data[8] ));
 sg13g2_antennanp ANTENNA_377 (.A(\soc_I.kianv_I.datapath_unit_I.Data[8] ));
 sg13g2_antennanp ANTENNA_378 (.A(\soc_I.kianv_I.datapath_unit_I.Data[9] ));
 sg13g2_antennanp ANTENNA_379 (.A(\soc_I.kianv_I.datapath_unit_I.Data[9] ));
 sg13g2_antennanp ANTENNA_380 (.A(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[17] ));
 sg13g2_antennanp ANTENNA_381 (.A(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[21] ));
 sg13g2_antennanp ANTENNA_382 (.A(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[8] ));
 sg13g2_antennanp ANTENNA_383 (.A(\soc_I.kianv_I.datapath_unit_I.MULExtResult[16] ));
 sg13g2_antennanp ANTENNA_384 (.A(\soc_I.kianv_I.datapath_unit_I.MULExtResult[25] ));
 sg13g2_antennanp ANTENNA_385 (.A(\soc_I.kianv_I.datapath_unit_I.MULExtResult[27] ));
 sg13g2_antennanp ANTENNA_386 (.A(\soc_I.kianv_I.datapath_unit_I.MULExtResult[28] ));
 sg13g2_antennanp ANTENNA_387 (.A(\soc_I.kianv_I.datapath_unit_I.MULExtResult[31] ));
 sg13g2_antennanp ANTENNA_388 (.A(uio_oe[1]));
 sg13g2_antennanp ANTENNA_389 (.A(uio_oe[1]));
 sg13g2_antennanp ANTENNA_390 (.A(uio_out[0]));
 sg13g2_antennanp ANTENNA_391 (.A(uio_out[0]));
 sg13g2_antennanp ANTENNA_392 (.A(uio_out[6]));
 sg13g2_antennanp ANTENNA_393 (.A(uio_out[6]));
 sg13g2_antennanp ANTENNA_394 (.A(uio_out[7]));
 sg13g2_antennanp ANTENNA_395 (.A(uio_out[7]));
 sg13g2_antennanp ANTENNA_396 (.A(net7490));
 sg13g2_antennanp ANTENNA_397 (.A(net7490));
 sg13g2_antennanp ANTENNA_398 (.A(net7490));
 sg13g2_antennanp ANTENNA_399 (.A(net7490));
 sg13g2_antennanp ANTENNA_400 (.A(net7510));
 sg13g2_antennanp ANTENNA_401 (.A(net7510));
 sg13g2_antennanp ANTENNA_402 (.A(net7510));
 sg13g2_antennanp ANTENNA_403 (.A(net7510));
 sg13g2_antennanp ANTENNA_404 (.A(net7533));
 sg13g2_antennanp ANTENNA_405 (.A(net7533));
 sg13g2_antennanp ANTENNA_406 (.A(net7533));
 sg13g2_antennanp ANTENNA_407 (.A(net7533));
 sg13g2_antennanp ANTENNA_408 (.A(net7533));
 sg13g2_antennanp ANTENNA_409 (.A(net7533));
 sg13g2_antennanp ANTENNA_410 (.A(net7618));
 sg13g2_antennanp ANTENNA_411 (.A(net7618));
 sg13g2_antennanp ANTENNA_412 (.A(net7618));
 sg13g2_antennanp ANTENNA_413 (.A(net7618));
 sg13g2_antennanp ANTENNA_414 (.A(net7618));
 sg13g2_antennanp ANTENNA_415 (.A(net7618));
 sg13g2_antennanp ANTENNA_416 (.A(net7618));
 sg13g2_antennanp ANTENNA_417 (.A(net7618));
 sg13g2_antennanp ANTENNA_418 (.A(net7618));
 sg13g2_antennanp ANTENNA_419 (.A(net7618));
 sg13g2_antennanp ANTENNA_420 (.A(net7618));
 sg13g2_antennanp ANTENNA_421 (.A(net7618));
 sg13g2_antennanp ANTENNA_422 (.A(net7618));
 sg13g2_antennanp ANTENNA_423 (.A(net7618));
 sg13g2_antennanp ANTENNA_424 (.A(net7618));
 sg13g2_antennanp ANTENNA_425 (.A(net7618));
 sg13g2_antennanp ANTENNA_426 (.A(net8597));
 sg13g2_antennanp ANTENNA_427 (.A(net8597));
 sg13g2_antennanp ANTENNA_428 (.A(net8597));
 sg13g2_antennanp ANTENNA_429 (.A(net8597));
 sg13g2_antennanp ANTENNA_430 (.A(net8597));
 sg13g2_antennanp ANTENNA_431 (.A(net8597));
 sg13g2_antennanp ANTENNA_432 (.A(net8597));
 sg13g2_antennanp ANTENNA_433 (.A(net8597));
 sg13g2_antennanp ANTENNA_434 (.A(net8597));
 sg13g2_antennanp ANTENNA_435 (.A(net8597));
 sg13g2_antennanp ANTENNA_436 (.A(net8597));
 sg13g2_antennanp ANTENNA_437 (.A(net8597));
 sg13g2_antennanp ANTENNA_438 (.A(net8597));
 sg13g2_antennanp ANTENNA_439 (.A(net8674));
 sg13g2_antennanp ANTENNA_440 (.A(net8674));
 sg13g2_antennanp ANTENNA_441 (.A(net8674));
 sg13g2_antennanp ANTENNA_442 (.A(net8674));
 sg13g2_antennanp ANTENNA_443 (.A(net8674));
 sg13g2_antennanp ANTENNA_444 (.A(net8674));
 sg13g2_antennanp ANTENNA_445 (.A(net8674));
 sg13g2_antennanp ANTENNA_446 (.A(net8674));
 sg13g2_antennanp ANTENNA_447 (.A(net8922));
 sg13g2_antennanp ANTENNA_448 (.A(net8922));
 sg13g2_antennanp ANTENNA_449 (.A(net8922));
 sg13g2_antennanp ANTENNA_450 (.A(net8922));
 sg13g2_antennanp ANTENNA_451 (.A(net8922));
 sg13g2_antennanp ANTENNA_452 (.A(net8922));
 sg13g2_antennanp ANTENNA_453 (.A(net8922));
 sg13g2_antennanp ANTENNA_454 (.A(net8922));
 sg13g2_antennanp ANTENNA_455 (.A(net8962));
 sg13g2_antennanp ANTENNA_456 (.A(net8962));
 sg13g2_antennanp ANTENNA_457 (.A(net8962));
 sg13g2_antennanp ANTENNA_458 (.A(net8962));
 sg13g2_antennanp ANTENNA_459 (.A(net8962));
 sg13g2_antennanp ANTENNA_460 (.A(net8962));
 sg13g2_antennanp ANTENNA_461 (.A(net8962));
 sg13g2_antennanp ANTENNA_462 (.A(net8962));
 sg13g2_antennanp ANTENNA_463 (.A(net8962));
 sg13g2_antennanp ANTENNA_464 (.A(net8962));
 sg13g2_antennanp ANTENNA_465 (.A(net8962));
 sg13g2_antennanp ANTENNA_466 (.A(net8962));
 sg13g2_antennanp ANTENNA_467 (.A(net8962));
 sg13g2_antennanp ANTENNA_468 (.A(net8962));
 sg13g2_antennanp ANTENNA_469 (.A(net8962));
 sg13g2_antennanp ANTENNA_470 (.A(net9001));
 sg13g2_antennanp ANTENNA_471 (.A(net9001));
 sg13g2_antennanp ANTENNA_472 (.A(net9001));
 sg13g2_antennanp ANTENNA_473 (.A(net9001));
 sg13g2_antennanp ANTENNA_474 (.A(net9001));
 sg13g2_antennanp ANTENNA_475 (.A(net9001));
 sg13g2_antennanp ANTENNA_476 (.A(net9001));
 sg13g2_antennanp ANTENNA_477 (.A(net9001));
 sg13g2_antennanp ANTENNA_478 (.A(net9001));
 sg13g2_antennanp ANTENNA_479 (.A(net9001));
 sg13g2_antennanp ANTENNA_480 (.A(net9001));
 sg13g2_antennanp ANTENNA_481 (.A(net9001));
 sg13g2_antennanp ANTENNA_482 (.A(net9001));
 sg13g2_antennanp ANTENNA_483 (.A(net9001));
 sg13g2_antennanp ANTENNA_484 (.A(net9001));
 sg13g2_antennanp ANTENNA_485 (.A(net9001));
 sg13g2_antennanp ANTENNA_486 (.A(net9439));
 sg13g2_antennanp ANTENNA_487 (.A(net9439));
 sg13g2_antennanp ANTENNA_488 (.A(net9439));
 sg13g2_antennanp ANTENNA_489 (.A(net9439));
 sg13g2_antennanp ANTENNA_490 (.A(net9439));
 sg13g2_antennanp ANTENNA_491 (.A(net9439));
 sg13g2_antennanp ANTENNA_492 (.A(net9439));
 sg13g2_antennanp ANTENNA_493 (.A(net9439));
 sg13g2_antennanp ANTENNA_494 (.A(net9439));
 sg13g2_antennanp ANTENNA_495 (.A(net9545));
 sg13g2_antennanp ANTENNA_496 (.A(net9545));
 sg13g2_antennanp ANTENNA_497 (.A(net9545));
 sg13g2_antennanp ANTENNA_498 (.A(net9545));
 sg13g2_antennanp ANTENNA_499 (.A(net10));
 sg13g2_antennanp ANTENNA_500 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_501 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_502 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_503 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_504 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_505 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_506 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_507 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_508 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_509 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_510 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_511 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_512 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_513 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_514 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_515 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_516 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_517 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_518 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_519 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_520 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_521 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_522 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_523 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_524 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_525 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_526 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_527 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_528 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_529 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_530 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_531 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_532 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_533 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_534 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_535 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_536 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_537 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_538 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_539 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_540 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_541 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_542 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_543 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_544 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_545 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_546 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_547 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_548 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_549 (.A(clknet_2_1_0_clk));
 sg13g2_antennanp ANTENNA_550 (.A(net5385));
 sg13g2_antennanp ANTENNA_551 (.A(_00187_));
 sg13g2_antennanp ANTENNA_552 (.A(_00187_));
 sg13g2_antennanp ANTENNA_553 (.A(_00187_));
 sg13g2_antennanp ANTENNA_554 (.A(_00187_));
 sg13g2_antennanp ANTENNA_555 (.A(_00225_));
 sg13g2_antennanp ANTENNA_556 (.A(_00229_));
 sg13g2_antennanp ANTENNA_557 (.A(_00230_));
 sg13g2_antennanp ANTENNA_558 (.A(_00231_));
 sg13g2_antennanp ANTENNA_559 (.A(_00232_));
 sg13g2_antennanp ANTENNA_560 (.A(_00233_));
 sg13g2_antennanp ANTENNA_561 (.A(_00235_));
 sg13g2_antennanp ANTENNA_562 (.A(_00742_));
 sg13g2_antennanp ANTENNA_563 (.A(_00743_));
 sg13g2_antennanp ANTENNA_564 (.A(_00750_));
 sg13g2_antennanp ANTENNA_565 (.A(_00751_));
 sg13g2_antennanp ANTENNA_566 (.A(_00752_));
 sg13g2_antennanp ANTENNA_567 (.A(_00754_));
 sg13g2_antennanp ANTENNA_568 (.A(_00762_));
 sg13g2_antennanp ANTENNA_569 (.A(_01001_));
 sg13g2_antennanp ANTENNA_570 (.A(_01002_));
 sg13g2_antennanp ANTENNA_571 (.A(_02684_));
 sg13g2_antennanp ANTENNA_572 (.A(_02690_));
 sg13g2_antennanp ANTENNA_573 (.A(_02691_));
 sg13g2_antennanp ANTENNA_574 (.A(_02698_));
 sg13g2_antennanp ANTENNA_575 (.A(_02701_));
 sg13g2_antennanp ANTENNA_576 (.A(_02707_));
 sg13g2_antennanp ANTENNA_577 (.A(_02710_));
 sg13g2_antennanp ANTENNA_578 (.A(_03370_));
 sg13g2_antennanp ANTENNA_579 (.A(_12499_));
 sg13g2_antennanp ANTENNA_580 (.A(_12499_));
 sg13g2_antennanp ANTENNA_581 (.A(_12499_));
 sg13g2_antennanp ANTENNA_582 (.A(_12499_));
 sg13g2_antennanp ANTENNA_583 (.A(_12787_));
 sg13g2_antennanp ANTENNA_584 (.A(_12795_));
 sg13g2_antennanp ANTENNA_585 (.A(_12893_));
 sg13g2_antennanp ANTENNA_586 (.A(_12893_));
 sg13g2_antennanp ANTENNA_587 (.A(_12893_));
 sg13g2_antennanp ANTENNA_588 (.A(_12893_));
 sg13g2_antennanp ANTENNA_589 (.A(_13836_));
 sg13g2_antennanp ANTENNA_590 (.A(_13836_));
 sg13g2_antennanp ANTENNA_591 (.A(_13836_));
 sg13g2_antennanp ANTENNA_592 (.A(_13836_));
 sg13g2_antennanp ANTENNA_593 (.A(_13974_));
 sg13g2_antennanp ANTENNA_594 (.A(_13974_));
 sg13g2_antennanp ANTENNA_595 (.A(_13974_));
 sg13g2_antennanp ANTENNA_596 (.A(_13974_));
 sg13g2_antennanp ANTENNA_597 (.A(_14059_));
 sg13g2_antennanp ANTENNA_598 (.A(_14080_));
 sg13g2_antennanp ANTENNA_599 (.A(_14086_));
 sg13g2_antennanp ANTENNA_600 (.A(_14090_));
 sg13g2_antennanp ANTENNA_601 (.A(_14097_));
 sg13g2_antennanp ANTENNA_602 (.A(_14109_));
 sg13g2_antennanp ANTENNA_603 (.A(clk));
 sg13g2_antennanp ANTENNA_604 (.A(clk));
 sg13g2_antennanp ANTENNA_605 (.A(\soc_I.clint_I.addr[1] ));
 sg13g2_antennanp ANTENNA_606 (.A(\soc_I.clint_I.addr[1] ));
 sg13g2_antennanp ANTENNA_607 (.A(\soc_I.clint_I.addr[1] ));
 sg13g2_antennanp ANTENNA_608 (.A(\soc_I.clint_I.addr[1] ));
 sg13g2_antennanp ANTENNA_609 (.A(\soc_I.clint_I.addr[1] ));
 sg13g2_antennanp ANTENNA_610 (.A(\soc_I.clint_I.addr[1] ));
 sg13g2_antennanp ANTENNA_611 (.A(\soc_I.clint_I.addr[1] ));
 sg13g2_antennanp ANTENNA_612 (.A(\soc_I.clint_I.addr[1] ));
 sg13g2_antennanp ANTENNA_613 (.A(\soc_I.clint_I.addr[1] ));
 sg13g2_antennanp ANTENNA_614 (.A(\soc_I.kianv_I.datapath_unit_I.A1[13] ));
 sg13g2_antennanp ANTENNA_615 (.A(\soc_I.kianv_I.datapath_unit_I.A1[20] ));
 sg13g2_antennanp ANTENNA_616 (.A(\soc_I.kianv_I.datapath_unit_I.A1[22] ));
 sg13g2_antennanp ANTENNA_617 (.A(\soc_I.kianv_I.datapath_unit_I.A1[26] ));
 sg13g2_antennanp ANTENNA_618 (.A(\soc_I.kianv_I.datapath_unit_I.A1[3] ));
 sg13g2_antennanp ANTENNA_619 (.A(\soc_I.kianv_I.datapath_unit_I.A1[4] ));
 sg13g2_antennanp ANTENNA_620 (.A(\soc_I.kianv_I.datapath_unit_I.A1[9] ));
 sg13g2_antennanp ANTENNA_621 (.A(\soc_I.kianv_I.datapath_unit_I.CSRDataOut[13] ));
 sg13g2_antennanp ANTENNA_622 (.A(\soc_I.kianv_I.datapath_unit_I.Data[9] ));
 sg13g2_antennanp ANTENNA_623 (.A(\soc_I.kianv_I.datapath_unit_I.Data[9] ));
 sg13g2_antennanp ANTENNA_624 (.A(\soc_I.kianv_I.datapath_unit_I.MULExtResultOut[8] ));
 sg13g2_antennanp ANTENNA_625 (.A(\soc_I.kianv_I.datapath_unit_I.MULExtResult[16] ));
 sg13g2_antennanp ANTENNA_626 (.A(\soc_I.kianv_I.datapath_unit_I.MULExtResult[28] ));
 sg13g2_antennanp ANTENNA_627 (.A(\soc_I.kianv_I.datapath_unit_I.MULExtResult[31] ));
 sg13g2_antennanp ANTENNA_628 (.A(uio_oe[1]));
 sg13g2_antennanp ANTENNA_629 (.A(uio_oe[1]));
 sg13g2_antennanp ANTENNA_630 (.A(uio_out[0]));
 sg13g2_antennanp ANTENNA_631 (.A(uio_out[0]));
 sg13g2_antennanp ANTENNA_632 (.A(uio_out[6]));
 sg13g2_antennanp ANTENNA_633 (.A(uio_out[6]));
 sg13g2_antennanp ANTENNA_634 (.A(uio_out[7]));
 sg13g2_antennanp ANTENNA_635 (.A(uio_out[7]));
 sg13g2_antennanp ANTENNA_636 (.A(net7490));
 sg13g2_antennanp ANTENNA_637 (.A(net7490));
 sg13g2_antennanp ANTENNA_638 (.A(net7490));
 sg13g2_antennanp ANTENNA_639 (.A(net7490));
 sg13g2_antennanp ANTENNA_640 (.A(net7510));
 sg13g2_antennanp ANTENNA_641 (.A(net7510));
 sg13g2_antennanp ANTENNA_642 (.A(net7510));
 sg13g2_antennanp ANTENNA_643 (.A(net7510));
 sg13g2_antennanp ANTENNA_644 (.A(net7618));
 sg13g2_antennanp ANTENNA_645 (.A(net7618));
 sg13g2_antennanp ANTENNA_646 (.A(net7618));
 sg13g2_antennanp ANTENNA_647 (.A(net7618));
 sg13g2_antennanp ANTENNA_648 (.A(net7618));
 sg13g2_antennanp ANTENNA_649 (.A(net7618));
 sg13g2_antennanp ANTENNA_650 (.A(net7618));
 sg13g2_antennanp ANTENNA_651 (.A(net7618));
 sg13g2_antennanp ANTENNA_652 (.A(net7618));
 sg13g2_antennanp ANTENNA_653 (.A(net7618));
 sg13g2_antennanp ANTENNA_654 (.A(net7618));
 sg13g2_antennanp ANTENNA_655 (.A(net7618));
 sg13g2_antennanp ANTENNA_656 (.A(net7618));
 sg13g2_antennanp ANTENNA_657 (.A(net7618));
 sg13g2_antennanp ANTENNA_658 (.A(net7618));
 sg13g2_antennanp ANTENNA_659 (.A(net7618));
 sg13g2_antennanp ANTENNA_660 (.A(net8674));
 sg13g2_antennanp ANTENNA_661 (.A(net8674));
 sg13g2_antennanp ANTENNA_662 (.A(net8674));
 sg13g2_antennanp ANTENNA_663 (.A(net8674));
 sg13g2_antennanp ANTENNA_664 (.A(net8674));
 sg13g2_antennanp ANTENNA_665 (.A(net8674));
 sg13g2_antennanp ANTENNA_666 (.A(net8674));
 sg13g2_antennanp ANTENNA_667 (.A(net8674));
 sg13g2_antennanp ANTENNA_668 (.A(net8962));
 sg13g2_antennanp ANTENNA_669 (.A(net8962));
 sg13g2_antennanp ANTENNA_670 (.A(net8962));
 sg13g2_antennanp ANTENNA_671 (.A(net8962));
 sg13g2_antennanp ANTENNA_672 (.A(net8962));
 sg13g2_antennanp ANTENNA_673 (.A(net8962));
 sg13g2_antennanp ANTENNA_674 (.A(net8962));
 sg13g2_antennanp ANTENNA_675 (.A(net8962));
 sg13g2_antennanp ANTENNA_676 (.A(net8962));
 sg13g2_antennanp ANTENNA_677 (.A(net8962));
 sg13g2_antennanp ANTENNA_678 (.A(net8962));
 sg13g2_antennanp ANTENNA_679 (.A(net8962));
 sg13g2_antennanp ANTENNA_680 (.A(net8962));
 sg13g2_antennanp ANTENNA_681 (.A(net8962));
 sg13g2_antennanp ANTENNA_682 (.A(net8962));
 sg13g2_antennanp ANTENNA_683 (.A(net9001));
 sg13g2_antennanp ANTENNA_684 (.A(net9001));
 sg13g2_antennanp ANTENNA_685 (.A(net9001));
 sg13g2_antennanp ANTENNA_686 (.A(net9001));
 sg13g2_antennanp ANTENNA_687 (.A(net9001));
 sg13g2_antennanp ANTENNA_688 (.A(net9001));
 sg13g2_antennanp ANTENNA_689 (.A(net9001));
 sg13g2_antennanp ANTENNA_690 (.A(net9001));
 sg13g2_antennanp ANTENNA_691 (.A(net9001));
 sg13g2_antennanp ANTENNA_692 (.A(net9001));
 sg13g2_antennanp ANTENNA_693 (.A(net9001));
 sg13g2_antennanp ANTENNA_694 (.A(net9001));
 sg13g2_antennanp ANTENNA_695 (.A(net9001));
 sg13g2_antennanp ANTENNA_696 (.A(net9001));
 sg13g2_antennanp ANTENNA_697 (.A(net9001));
 sg13g2_antennanp ANTENNA_698 (.A(net9001));
 sg13g2_antennanp ANTENNA_699 (.A(net10));
 sg13g2_antennanp ANTENNA_700 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_701 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_702 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_703 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_704 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_705 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_706 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_707 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_708 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_709 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_710 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_711 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_712 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_713 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_714 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_715 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_716 (.A(net5385));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_fill_2 FILLER_0_21 ();
 sg13g2_decap_4 FILLER_0_95 ();
 sg13g2_fill_2 FILLER_0_99 ();
 sg13g2_decap_4 FILLER_0_127 ();
 sg13g2_decap_8 FILLER_0_157 ();
 sg13g2_decap_4 FILLER_0_164 ();
 sg13g2_fill_1 FILLER_0_198 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_fill_2 FILLER_0_210 ();
 sg13g2_fill_1 FILLER_0_212 ();
 sg13g2_fill_2 FILLER_0_232 ();
 sg13g2_decap_4 FILLER_0_243 ();
 sg13g2_fill_1 FILLER_0_247 ();
 sg13g2_decap_8 FILLER_0_274 ();
 sg13g2_fill_2 FILLER_0_281 ();
 sg13g2_fill_1 FILLER_0_283 ();
 sg13g2_fill_1 FILLER_0_293 ();
 sg13g2_fill_1 FILLER_0_308 ();
 sg13g2_decap_4 FILLER_0_337 ();
 sg13g2_fill_1 FILLER_0_341 ();
 sg13g2_fill_2 FILLER_0_346 ();
 sg13g2_fill_1 FILLER_0_348 ();
 sg13g2_decap_8 FILLER_0_362 ();
 sg13g2_decap_4 FILLER_0_369 ();
 sg13g2_fill_2 FILLER_0_373 ();
 sg13g2_decap_4 FILLER_0_380 ();
 sg13g2_fill_1 FILLER_0_384 ();
 sg13g2_decap_8 FILLER_0_415 ();
 sg13g2_decap_4 FILLER_0_422 ();
 sg13g2_fill_2 FILLER_0_448 ();
 sg13g2_fill_2 FILLER_0_455 ();
 sg13g2_fill_1 FILLER_0_457 ();
 sg13g2_decap_4 FILLER_0_466 ();
 sg13g2_fill_2 FILLER_0_470 ();
 sg13g2_fill_2 FILLER_0_502 ();
 sg13g2_fill_1 FILLER_0_504 ();
 sg13g2_fill_2 FILLER_0_510 ();
 sg13g2_fill_1 FILLER_0_512 ();
 sg13g2_decap_8 FILLER_0_517 ();
 sg13g2_decap_8 FILLER_0_524 ();
 sg13g2_fill_2 FILLER_0_536 ();
 sg13g2_fill_1 FILLER_0_538 ();
 sg13g2_decap_8 FILLER_0_543 ();
 sg13g2_decap_4 FILLER_0_550 ();
 sg13g2_fill_1 FILLER_0_554 ();
 sg13g2_fill_2 FILLER_0_563 ();
 sg13g2_fill_1 FILLER_0_565 ();
 sg13g2_fill_2 FILLER_0_571 ();
 sg13g2_fill_1 FILLER_0_573 ();
 sg13g2_decap_8 FILLER_0_578 ();
 sg13g2_fill_2 FILLER_0_585 ();
 sg13g2_decap_4 FILLER_0_592 ();
 sg13g2_fill_2 FILLER_0_596 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_fill_1 FILLER_0_616 ();
 sg13g2_fill_1 FILLER_0_643 ();
 sg13g2_fill_2 FILLER_0_649 ();
 sg13g2_fill_1 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_656 ();
 sg13g2_decap_8 FILLER_0_663 ();
 sg13g2_fill_2 FILLER_0_670 ();
 sg13g2_fill_1 FILLER_0_672 ();
 sg13g2_fill_1 FILLER_0_682 ();
 sg13g2_decap_4 FILLER_0_692 ();
 sg13g2_fill_1 FILLER_0_696 ();
 sg13g2_fill_1 FILLER_0_701 ();
 sg13g2_decap_8 FILLER_0_720 ();
 sg13g2_decap_4 FILLER_0_727 ();
 sg13g2_decap_4 FILLER_0_739 ();
 sg13g2_fill_1 FILLER_0_743 ();
 sg13g2_fill_2 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_4 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_792 ();
 sg13g2_fill_2 FILLER_0_799 ();
 sg13g2_fill_1 FILLER_0_801 ();
 sg13g2_fill_2 FILLER_0_807 ();
 sg13g2_fill_1 FILLER_0_809 ();
 sg13g2_decap_8 FILLER_0_814 ();
 sg13g2_decap_8 FILLER_0_821 ();
 sg13g2_decap_4 FILLER_0_828 ();
 sg13g2_fill_2 FILLER_0_837 ();
 sg13g2_fill_1 FILLER_0_839 ();
 sg13g2_decap_8 FILLER_0_844 ();
 sg13g2_fill_2 FILLER_0_851 ();
 sg13g2_decap_8 FILLER_0_858 ();
 sg13g2_decap_8 FILLER_0_869 ();
 sg13g2_decap_8 FILLER_0_876 ();
 sg13g2_fill_2 FILLER_0_883 ();
 sg13g2_fill_1 FILLER_0_890 ();
 sg13g2_fill_2 FILLER_0_899 ();
 sg13g2_fill_2 FILLER_0_918 ();
 sg13g2_fill_1 FILLER_0_925 ();
 sg13g2_decap_8 FILLER_0_931 ();
 sg13g2_decap_8 FILLER_0_938 ();
 sg13g2_fill_2 FILLER_0_945 ();
 sg13g2_fill_1 FILLER_0_947 ();
 sg13g2_fill_2 FILLER_0_956 ();
 sg13g2_fill_1 FILLER_0_958 ();
 sg13g2_decap_8 FILLER_0_963 ();
 sg13g2_decap_4 FILLER_0_970 ();
 sg13g2_fill_1 FILLER_0_974 ();
 sg13g2_fill_2 FILLER_0_980 ();
 sg13g2_fill_1 FILLER_0_982 ();
 sg13g2_decap_8 FILLER_0_991 ();
 sg13g2_decap_4 FILLER_0_998 ();
 sg13g2_decap_4 FILLER_0_1032 ();
 sg13g2_decap_8 FILLER_0_1062 ();
 sg13g2_decap_4 FILLER_0_1069 ();
 sg13g2_decap_8 FILLER_0_1086 ();
 sg13g2_fill_1 FILLER_0_1093 ();
 sg13g2_decap_8 FILLER_0_1120 ();
 sg13g2_fill_2 FILLER_0_1127 ();
 sg13g2_fill_2 FILLER_0_1134 ();
 sg13g2_fill_2 FILLER_0_1144 ();
 sg13g2_fill_2 FILLER_0_1160 ();
 sg13g2_decap_4 FILLER_0_1170 ();
 sg13g2_fill_1 FILLER_0_1174 ();
 sg13g2_fill_2 FILLER_0_1209 ();
 sg13g2_fill_2 FILLER_0_1216 ();
 sg13g2_fill_1 FILLER_0_1218 ();
 sg13g2_decap_8 FILLER_0_1223 ();
 sg13g2_fill_1 FILLER_0_1230 ();
 sg13g2_fill_2 FILLER_0_1239 ();
 sg13g2_fill_2 FILLER_0_1245 ();
 sg13g2_fill_1 FILLER_0_1247 ();
 sg13g2_decap_4 FILLER_0_1261 ();
 sg13g2_decap_4 FILLER_0_1270 ();
 sg13g2_fill_2 FILLER_0_1278 ();
 sg13g2_fill_1 FILLER_0_1280 ();
 sg13g2_fill_2 FILLER_0_1295 ();
 sg13g2_decap_8 FILLER_0_1323 ();
 sg13g2_decap_8 FILLER_0_1330 ();
 sg13g2_decap_4 FILLER_0_1337 ();
 sg13g2_fill_2 FILLER_0_1341 ();
 sg13g2_fill_1 FILLER_0_1348 ();
 sg13g2_fill_2 FILLER_0_1353 ();
 sg13g2_fill_1 FILLER_0_1355 ();
 sg13g2_fill_1 FILLER_0_1360 ();
 sg13g2_decap_8 FILLER_0_1370 ();
 sg13g2_fill_1 FILLER_0_1377 ();
 sg13g2_fill_2 FILLER_0_1383 ();
 sg13g2_decap_8 FILLER_0_1389 ();
 sg13g2_fill_1 FILLER_0_1396 ();
 sg13g2_fill_2 FILLER_0_1431 ();
 sg13g2_fill_2 FILLER_0_1438 ();
 sg13g2_fill_2 FILLER_0_1448 ();
 sg13g2_decap_4 FILLER_0_1459 ();
 sg13g2_fill_2 FILLER_0_1463 ();
 sg13g2_fill_2 FILLER_0_1470 ();
 sg13g2_decap_4 FILLER_0_1476 ();
 sg13g2_fill_1 FILLER_0_1489 ();
 sg13g2_fill_2 FILLER_0_1495 ();
 sg13g2_fill_1 FILLER_0_1497 ();
 sg13g2_fill_2 FILLER_0_1506 ();
 sg13g2_decap_4 FILLER_0_1517 ();
 sg13g2_fill_1 FILLER_0_1521 ();
 sg13g2_fill_1 FILLER_0_1527 ();
 sg13g2_fill_2 FILLER_0_1532 ();
 sg13g2_fill_2 FILLER_0_1543 ();
 sg13g2_fill_1 FILLER_0_1545 ();
 sg13g2_fill_1 FILLER_0_1551 ();
 sg13g2_decap_8 FILLER_0_1556 ();
 sg13g2_decap_4 FILLER_0_1563 ();
 sg13g2_fill_1 FILLER_0_1567 ();
 sg13g2_fill_2 FILLER_0_1598 ();
 sg13g2_fill_2 FILLER_0_1604 ();
 sg13g2_fill_2 FILLER_0_1619 ();
 sg13g2_fill_1 FILLER_0_1621 ();
 sg13g2_decap_4 FILLER_0_1627 ();
 sg13g2_fill_1 FILLER_0_1631 ();
 sg13g2_decap_4 FILLER_0_1636 ();
 sg13g2_fill_1 FILLER_0_1640 ();
 sg13g2_decap_8 FILLER_0_1646 ();
 sg13g2_decap_4 FILLER_0_1653 ();
 sg13g2_fill_1 FILLER_0_1657 ();
 sg13g2_decap_4 FILLER_0_1667 ();
 sg13g2_fill_1 FILLER_0_1671 ();
 sg13g2_decap_8 FILLER_0_1702 ();
 sg13g2_fill_2 FILLER_0_1709 ();
 sg13g2_fill_1 FILLER_0_1711 ();
 sg13g2_fill_2 FILLER_0_1716 ();
 sg13g2_decap_4 FILLER_0_1731 ();
 sg13g2_fill_2 FILLER_0_1735 ();
 sg13g2_fill_2 FILLER_0_1746 ();
 sg13g2_fill_1 FILLER_0_1748 ();
 sg13g2_fill_2 FILLER_0_1767 ();
 sg13g2_fill_1 FILLER_0_1773 ();
 sg13g2_fill_1 FILLER_0_1783 ();
 sg13g2_decap_8 FILLER_0_1797 ();
 sg13g2_fill_2 FILLER_0_1804 ();
 sg13g2_fill_2 FILLER_0_1815 ();
 sg13g2_decap_8 FILLER_0_1843 ();
 sg13g2_decap_8 FILLER_0_1850 ();
 sg13g2_decap_8 FILLER_0_1861 ();
 sg13g2_decap_8 FILLER_0_1868 ();
 sg13g2_fill_2 FILLER_0_1879 ();
 sg13g2_fill_2 FILLER_0_1885 ();
 sg13g2_fill_1 FILLER_0_1887 ();
 sg13g2_decap_8 FILLER_0_1906 ();
 sg13g2_fill_1 FILLER_0_1913 ();
 sg13g2_decap_4 FILLER_0_1932 ();
 sg13g2_fill_1 FILLER_0_1940 ();
 sg13g2_decap_8 FILLER_0_1950 ();
 sg13g2_fill_2 FILLER_0_1957 ();
 sg13g2_fill_1 FILLER_0_1959 ();
 sg13g2_decap_8 FILLER_0_1977 ();
 sg13g2_fill_2 FILLER_0_1984 ();
 sg13g2_fill_1 FILLER_0_1986 ();
 sg13g2_fill_2 FILLER_0_1992 ();
 sg13g2_decap_8 FILLER_0_2007 ();
 sg13g2_fill_2 FILLER_0_2014 ();
 sg13g2_decap_8 FILLER_0_2021 ();
 sg13g2_fill_1 FILLER_0_2028 ();
 sg13g2_decap_8 FILLER_0_2033 ();
 sg13g2_decap_8 FILLER_0_2040 ();
 sg13g2_fill_2 FILLER_0_2047 ();
 sg13g2_fill_1 FILLER_0_2049 ();
 sg13g2_decap_8 FILLER_0_2076 ();
 sg13g2_decap_4 FILLER_0_2083 ();
 sg13g2_fill_1 FILLER_0_2087 ();
 sg13g2_fill_1 FILLER_0_2096 ();
 sg13g2_decap_4 FILLER_0_2128 ();
 sg13g2_fill_1 FILLER_0_2132 ();
 sg13g2_fill_2 FILLER_0_2163 ();
 sg13g2_decap_8 FILLER_0_2195 ();
 sg13g2_decap_8 FILLER_0_2202 ();
 sg13g2_decap_8 FILLER_0_2209 ();
 sg13g2_fill_2 FILLER_0_2216 ();
 sg13g2_fill_1 FILLER_0_2218 ();
 sg13g2_decap_8 FILLER_0_2224 ();
 sg13g2_decap_4 FILLER_0_2231 ();
 sg13g2_fill_2 FILLER_0_2235 ();
 sg13g2_fill_1 FILLER_0_2241 ();
 sg13g2_decap_8 FILLER_0_2246 ();
 sg13g2_decap_8 FILLER_0_2253 ();
 sg13g2_fill_2 FILLER_0_2260 ();
 sg13g2_fill_1 FILLER_0_2267 ();
 sg13g2_decap_8 FILLER_0_2272 ();
 sg13g2_fill_2 FILLER_0_2279 ();
 sg13g2_fill_1 FILLER_0_2281 ();
 sg13g2_fill_2 FILLER_0_2308 ();
 sg13g2_fill_1 FILLER_0_2310 ();
 sg13g2_decap_4 FILLER_0_2337 ();
 sg13g2_fill_2 FILLER_0_2341 ();
 sg13g2_fill_2 FILLER_0_2348 ();
 sg13g2_fill_1 FILLER_0_2350 ();
 sg13g2_decap_8 FILLER_0_2355 ();
 sg13g2_fill_2 FILLER_0_2362 ();
 sg13g2_decap_4 FILLER_0_2368 ();
 sg13g2_fill_1 FILLER_0_2372 ();
 sg13g2_decap_8 FILLER_0_2387 ();
 sg13g2_decap_8 FILLER_0_2398 ();
 sg13g2_decap_8 FILLER_0_2405 ();
 sg13g2_decap_8 FILLER_0_2412 ();
 sg13g2_decap_8 FILLER_0_2419 ();
 sg13g2_decap_4 FILLER_0_2426 ();
 sg13g2_decap_8 FILLER_0_2434 ();
 sg13g2_decap_4 FILLER_0_2441 ();
 sg13g2_fill_1 FILLER_0_2445 ();
 sg13g2_fill_2 FILLER_0_2451 ();
 sg13g2_fill_1 FILLER_0_2453 ();
 sg13g2_fill_1 FILLER_0_2458 ();
 sg13g2_decap_8 FILLER_0_2467 ();
 sg13g2_decap_4 FILLER_0_2474 ();
 sg13g2_decap_8 FILLER_0_2500 ();
 sg13g2_fill_2 FILLER_0_2507 ();
 sg13g2_fill_1 FILLER_0_2509 ();
 sg13g2_decap_4 FILLER_0_2519 ();
 sg13g2_fill_1 FILLER_0_2523 ();
 sg13g2_fill_1 FILLER_0_2537 ();
 sg13g2_fill_2 FILLER_0_2542 ();
 sg13g2_fill_1 FILLER_0_2544 ();
 sg13g2_decap_4 FILLER_0_2554 ();
 sg13g2_fill_2 FILLER_0_2558 ();
 sg13g2_fill_2 FILLER_0_2590 ();
 sg13g2_decap_4 FILLER_0_2596 ();
 sg13g2_decap_8 FILLER_0_2613 ();
 sg13g2_decap_8 FILLER_0_2620 ();
 sg13g2_decap_8 FILLER_0_2627 ();
 sg13g2_decap_8 FILLER_0_2634 ();
 sg13g2_decap_8 FILLER_0_2641 ();
 sg13g2_decap_8 FILLER_0_2648 ();
 sg13g2_decap_8 FILLER_0_2655 ();
 sg13g2_decap_8 FILLER_0_2662 ();
 sg13g2_fill_2 FILLER_0_2669 ();
 sg13g2_fill_1 FILLER_0_2675 ();
 sg13g2_decap_4 FILLER_0_2681 ();
 sg13g2_fill_1 FILLER_0_2685 ();
 sg13g2_decap_8 FILLER_0_2690 ();
 sg13g2_fill_2 FILLER_0_2697 ();
 sg13g2_fill_2 FILLER_0_2704 ();
 sg13g2_decap_8 FILLER_0_2710 ();
 sg13g2_decap_4 FILLER_0_2717 ();
 sg13g2_fill_1 FILLER_0_2721 ();
 sg13g2_decap_8 FILLER_0_2735 ();
 sg13g2_decap_4 FILLER_0_2742 ();
 sg13g2_fill_1 FILLER_0_2746 ();
 sg13g2_decap_8 FILLER_0_2777 ();
 sg13g2_decap_8 FILLER_0_2784 ();
 sg13g2_decap_8 FILLER_0_2791 ();
 sg13g2_decap_8 FILLER_0_2798 ();
 sg13g2_decap_8 FILLER_0_2805 ();
 sg13g2_decap_8 FILLER_0_2812 ();
 sg13g2_decap_8 FILLER_0_2819 ();
 sg13g2_decap_8 FILLER_0_2826 ();
 sg13g2_decap_8 FILLER_0_2833 ();
 sg13g2_decap_8 FILLER_0_2840 ();
 sg13g2_decap_8 FILLER_0_2847 ();
 sg13g2_decap_8 FILLER_0_2854 ();
 sg13g2_decap_8 FILLER_0_2861 ();
 sg13g2_decap_8 FILLER_0_2868 ();
 sg13g2_decap_8 FILLER_0_2875 ();
 sg13g2_decap_8 FILLER_0_2882 ();
 sg13g2_decap_8 FILLER_0_2889 ();
 sg13g2_decap_8 FILLER_0_2896 ();
 sg13g2_decap_8 FILLER_0_2903 ();
 sg13g2_decap_8 FILLER_0_2910 ();
 sg13g2_decap_8 FILLER_0_2917 ();
 sg13g2_decap_8 FILLER_0_2924 ();
 sg13g2_decap_8 FILLER_0_2931 ();
 sg13g2_decap_8 FILLER_0_2938 ();
 sg13g2_decap_8 FILLER_0_2945 ();
 sg13g2_decap_8 FILLER_0_2952 ();
 sg13g2_decap_8 FILLER_0_2959 ();
 sg13g2_decap_8 FILLER_0_2966 ();
 sg13g2_decap_8 FILLER_0_2973 ();
 sg13g2_decap_8 FILLER_0_2980 ();
 sg13g2_decap_8 FILLER_0_2987 ();
 sg13g2_decap_8 FILLER_0_2994 ();
 sg13g2_decap_8 FILLER_0_3001 ();
 sg13g2_decap_8 FILLER_0_3008 ();
 sg13g2_decap_8 FILLER_0_3015 ();
 sg13g2_decap_8 FILLER_0_3022 ();
 sg13g2_decap_8 FILLER_0_3029 ();
 sg13g2_decap_8 FILLER_0_3036 ();
 sg13g2_decap_8 FILLER_0_3043 ();
 sg13g2_decap_8 FILLER_0_3050 ();
 sg13g2_decap_8 FILLER_0_3057 ();
 sg13g2_decap_8 FILLER_0_3064 ();
 sg13g2_decap_8 FILLER_0_3071 ();
 sg13g2_decap_8 FILLER_0_3078 ();
 sg13g2_decap_8 FILLER_0_3085 ();
 sg13g2_decap_8 FILLER_0_3092 ();
 sg13g2_decap_8 FILLER_0_3099 ();
 sg13g2_decap_8 FILLER_0_3106 ();
 sg13g2_decap_8 FILLER_0_3113 ();
 sg13g2_decap_8 FILLER_0_3120 ();
 sg13g2_decap_8 FILLER_0_3127 ();
 sg13g2_decap_8 FILLER_0_3134 ();
 sg13g2_decap_8 FILLER_0_3141 ();
 sg13g2_decap_8 FILLER_0_3148 ();
 sg13g2_decap_8 FILLER_0_3155 ();
 sg13g2_decap_8 FILLER_0_3162 ();
 sg13g2_decap_8 FILLER_0_3169 ();
 sg13g2_decap_8 FILLER_0_3176 ();
 sg13g2_decap_8 FILLER_0_3183 ();
 sg13g2_decap_8 FILLER_0_3190 ();
 sg13g2_decap_8 FILLER_0_3197 ();
 sg13g2_decap_8 FILLER_0_3204 ();
 sg13g2_decap_8 FILLER_0_3211 ();
 sg13g2_decap_8 FILLER_0_3218 ();
 sg13g2_decap_8 FILLER_0_3225 ();
 sg13g2_decap_8 FILLER_0_3232 ();
 sg13g2_decap_8 FILLER_0_3239 ();
 sg13g2_decap_8 FILLER_0_3246 ();
 sg13g2_decap_8 FILLER_0_3253 ();
 sg13g2_decap_8 FILLER_0_3260 ();
 sg13g2_decap_8 FILLER_0_3267 ();
 sg13g2_decap_8 FILLER_0_3274 ();
 sg13g2_decap_8 FILLER_0_3281 ();
 sg13g2_decap_8 FILLER_0_3288 ();
 sg13g2_decap_8 FILLER_0_3295 ();
 sg13g2_decap_8 FILLER_0_3302 ();
 sg13g2_decap_8 FILLER_0_3309 ();
 sg13g2_decap_8 FILLER_0_3316 ();
 sg13g2_decap_8 FILLER_0_3323 ();
 sg13g2_decap_8 FILLER_0_3330 ();
 sg13g2_decap_8 FILLER_0_3337 ();
 sg13g2_decap_8 FILLER_0_3344 ();
 sg13g2_decap_8 FILLER_0_3351 ();
 sg13g2_decap_8 FILLER_0_3358 ();
 sg13g2_decap_8 FILLER_0_3365 ();
 sg13g2_decap_8 FILLER_0_3372 ();
 sg13g2_decap_8 FILLER_0_3379 ();
 sg13g2_decap_8 FILLER_0_3386 ();
 sg13g2_decap_8 FILLER_0_3393 ();
 sg13g2_decap_8 FILLER_0_3400 ();
 sg13g2_decap_8 FILLER_0_3407 ();
 sg13g2_decap_8 FILLER_0_3414 ();
 sg13g2_decap_8 FILLER_0_3421 ();
 sg13g2_decap_8 FILLER_0_3428 ();
 sg13g2_decap_8 FILLER_0_3435 ();
 sg13g2_decap_8 FILLER_0_3442 ();
 sg13g2_decap_8 FILLER_0_3449 ();
 sg13g2_decap_8 FILLER_0_3456 ();
 sg13g2_decap_8 FILLER_0_3463 ();
 sg13g2_decap_8 FILLER_0_3470 ();
 sg13g2_decap_8 FILLER_0_3477 ();
 sg13g2_decap_8 FILLER_0_3484 ();
 sg13g2_decap_8 FILLER_0_3491 ();
 sg13g2_decap_8 FILLER_0_3498 ();
 sg13g2_decap_8 FILLER_0_3505 ();
 sg13g2_decap_8 FILLER_0_3512 ();
 sg13g2_decap_8 FILLER_0_3519 ();
 sg13g2_decap_8 FILLER_0_3526 ();
 sg13g2_decap_8 FILLER_0_3533 ();
 sg13g2_decap_8 FILLER_0_3540 ();
 sg13g2_decap_8 FILLER_0_3547 ();
 sg13g2_decap_8 FILLER_0_3554 ();
 sg13g2_decap_8 FILLER_0_3561 ();
 sg13g2_decap_8 FILLER_0_3568 ();
 sg13g2_decap_4 FILLER_0_3575 ();
 sg13g2_fill_1 FILLER_0_3579 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_4 FILLER_1_14 ();
 sg13g2_fill_1 FILLER_1_18 ();
 sg13g2_decap_8 FILLER_1_76 ();
 sg13g2_fill_2 FILLER_1_83 ();
 sg13g2_fill_1 FILLER_1_85 ();
 sg13g2_decap_8 FILLER_1_96 ();
 sg13g2_fill_2 FILLER_1_103 ();
 sg13g2_fill_2 FILLER_1_115 ();
 sg13g2_decap_4 FILLER_1_149 ();
 sg13g2_fill_2 FILLER_1_153 ();
 sg13g2_fill_2 FILLER_1_214 ();
 sg13g2_decap_8 FILLER_1_265 ();
 sg13g2_fill_2 FILLER_1_272 ();
 sg13g2_fill_2 FILLER_1_388 ();
 sg13g2_fill_1 FILLER_1_404 ();
 sg13g2_fill_2 FILLER_1_444 ();
 sg13g2_fill_1 FILLER_1_446 ();
 sg13g2_fill_2 FILLER_1_478 ();
 sg13g2_fill_1 FILLER_1_480 ();
 sg13g2_fill_2 FILLER_1_485 ();
 sg13g2_fill_2 FILLER_1_500 ();
 sg13g2_fill_2 FILLER_1_554 ();
 sg13g2_fill_1 FILLER_1_712 ();
 sg13g2_fill_2 FILLER_1_753 ();
 sg13g2_fill_2 FILLER_1_826 ();
 sg13g2_decap_4 FILLER_1_906 ();
 sg13g2_fill_2 FILLER_1_910 ();
 sg13g2_fill_2 FILLER_1_1012 ();
 sg13g2_fill_2 FILLER_1_1045 ();
 sg13g2_fill_2 FILLER_1_1064 ();
 sg13g2_fill_1 FILLER_1_1066 ();
 sg13g2_decap_8 FILLER_1_1115 ();
 sg13g2_fill_2 FILLER_1_1122 ();
 sg13g2_fill_1 FILLER_1_1124 ();
 sg13g2_fill_2 FILLER_1_1191 ();
 sg13g2_fill_2 FILLER_1_1206 ();
 sg13g2_fill_1 FILLER_1_1234 ();
 sg13g2_fill_2 FILLER_1_1287 ();
 sg13g2_decap_8 FILLER_1_1329 ();
 sg13g2_fill_1 FILLER_1_1336 ();
 sg13g2_decap_4 FILLER_1_1455 ();
 sg13g2_fill_1 FILLER_1_1459 ();
 sg13g2_fill_1 FILLER_1_1486 ();
 sg13g2_fill_2 FILLER_1_1574 ();
 sg13g2_fill_1 FILLER_1_1576 ();
 sg13g2_fill_1 FILLER_1_1591 ();
 sg13g2_decap_8 FILLER_1_1670 ();
 sg13g2_decap_4 FILLER_1_1677 ();
 sg13g2_fill_2 FILLER_1_1681 ();
 sg13g2_fill_2 FILLER_1_1817 ();
 sg13g2_fill_1 FILLER_1_1819 ();
 sg13g2_fill_1 FILLER_1_1846 ();
 sg13g2_fill_1 FILLER_1_1925 ();
 sg13g2_decap_4 FILLER_1_2044 ();
 sg13g2_fill_2 FILLER_1_2057 ();
 sg13g2_fill_1 FILLER_1_2059 ();
 sg13g2_fill_1 FILLER_1_2064 ();
 sg13g2_decap_8 FILLER_1_2074 ();
 sg13g2_decap_4 FILLER_1_2081 ();
 sg13g2_fill_1 FILLER_1_2085 ();
 sg13g2_fill_1 FILLER_1_2112 ();
 sg13g2_fill_2 FILLER_1_2139 ();
 sg13g2_fill_1 FILLER_1_2141 ();
 sg13g2_fill_2 FILLER_1_2169 ();
 sg13g2_fill_1 FILLER_1_2171 ();
 sg13g2_fill_2 FILLER_1_2177 ();
 sg13g2_fill_1 FILLER_1_2179 ();
 sg13g2_fill_1 FILLER_1_2309 ();
 sg13g2_fill_1 FILLER_1_2323 ();
 sg13g2_fill_2 FILLER_1_2333 ();
 sg13g2_fill_1 FILLER_1_2418 ();
 sg13g2_fill_1 FILLER_1_2471 ();
 sg13g2_decap_8 FILLER_1_2498 ();
 sg13g2_fill_2 FILLER_1_2566 ();
 sg13g2_fill_2 FILLER_1_2572 ();
 sg13g2_fill_1 FILLER_1_2574 ();
 sg13g2_decap_8 FILLER_1_2641 ();
 sg13g2_decap_8 FILLER_1_2648 ();
 sg13g2_decap_4 FILLER_1_2655 ();
 sg13g2_fill_1 FILLER_1_2659 ();
 sg13g2_fill_2 FILLER_1_2747 ();
 sg13g2_decap_4 FILLER_1_2781 ();
 sg13g2_decap_4 FILLER_1_2815 ();
 sg13g2_decap_8 FILLER_1_2828 ();
 sg13g2_fill_2 FILLER_1_2835 ();
 sg13g2_decap_8 FILLER_1_2846 ();
 sg13g2_decap_8 FILLER_1_2853 ();
 sg13g2_decap_8 FILLER_1_2860 ();
 sg13g2_decap_8 FILLER_1_2867 ();
 sg13g2_decap_8 FILLER_1_2874 ();
 sg13g2_decap_8 FILLER_1_2881 ();
 sg13g2_decap_8 FILLER_1_2888 ();
 sg13g2_decap_8 FILLER_1_2895 ();
 sg13g2_decap_8 FILLER_1_2902 ();
 sg13g2_decap_8 FILLER_1_2909 ();
 sg13g2_decap_8 FILLER_1_2916 ();
 sg13g2_decap_8 FILLER_1_2923 ();
 sg13g2_decap_8 FILLER_1_2930 ();
 sg13g2_decap_8 FILLER_1_2937 ();
 sg13g2_decap_8 FILLER_1_2944 ();
 sg13g2_decap_8 FILLER_1_2951 ();
 sg13g2_decap_8 FILLER_1_2958 ();
 sg13g2_decap_8 FILLER_1_2965 ();
 sg13g2_decap_8 FILLER_1_2972 ();
 sg13g2_decap_8 FILLER_1_2979 ();
 sg13g2_decap_8 FILLER_1_2986 ();
 sg13g2_decap_8 FILLER_1_2993 ();
 sg13g2_decap_8 FILLER_1_3000 ();
 sg13g2_decap_8 FILLER_1_3007 ();
 sg13g2_decap_8 FILLER_1_3014 ();
 sg13g2_decap_8 FILLER_1_3021 ();
 sg13g2_decap_8 FILLER_1_3028 ();
 sg13g2_decap_8 FILLER_1_3035 ();
 sg13g2_decap_8 FILLER_1_3042 ();
 sg13g2_decap_8 FILLER_1_3049 ();
 sg13g2_decap_8 FILLER_1_3056 ();
 sg13g2_decap_8 FILLER_1_3063 ();
 sg13g2_decap_8 FILLER_1_3070 ();
 sg13g2_decap_8 FILLER_1_3077 ();
 sg13g2_decap_8 FILLER_1_3084 ();
 sg13g2_decap_8 FILLER_1_3091 ();
 sg13g2_decap_8 FILLER_1_3098 ();
 sg13g2_decap_8 FILLER_1_3105 ();
 sg13g2_decap_8 FILLER_1_3112 ();
 sg13g2_decap_8 FILLER_1_3119 ();
 sg13g2_decap_8 FILLER_1_3126 ();
 sg13g2_decap_8 FILLER_1_3133 ();
 sg13g2_decap_8 FILLER_1_3140 ();
 sg13g2_decap_8 FILLER_1_3147 ();
 sg13g2_decap_8 FILLER_1_3154 ();
 sg13g2_decap_8 FILLER_1_3161 ();
 sg13g2_decap_8 FILLER_1_3168 ();
 sg13g2_decap_8 FILLER_1_3175 ();
 sg13g2_decap_8 FILLER_1_3182 ();
 sg13g2_decap_8 FILLER_1_3189 ();
 sg13g2_decap_8 FILLER_1_3196 ();
 sg13g2_decap_8 FILLER_1_3203 ();
 sg13g2_decap_8 FILLER_1_3210 ();
 sg13g2_decap_8 FILLER_1_3217 ();
 sg13g2_decap_8 FILLER_1_3224 ();
 sg13g2_decap_8 FILLER_1_3231 ();
 sg13g2_decap_8 FILLER_1_3238 ();
 sg13g2_decap_8 FILLER_1_3245 ();
 sg13g2_decap_8 FILLER_1_3252 ();
 sg13g2_decap_8 FILLER_1_3259 ();
 sg13g2_decap_8 FILLER_1_3266 ();
 sg13g2_decap_8 FILLER_1_3273 ();
 sg13g2_decap_8 FILLER_1_3280 ();
 sg13g2_decap_8 FILLER_1_3287 ();
 sg13g2_decap_8 FILLER_1_3294 ();
 sg13g2_decap_8 FILLER_1_3301 ();
 sg13g2_decap_8 FILLER_1_3308 ();
 sg13g2_decap_8 FILLER_1_3315 ();
 sg13g2_decap_8 FILLER_1_3322 ();
 sg13g2_decap_8 FILLER_1_3329 ();
 sg13g2_decap_8 FILLER_1_3336 ();
 sg13g2_decap_8 FILLER_1_3343 ();
 sg13g2_decap_8 FILLER_1_3350 ();
 sg13g2_decap_8 FILLER_1_3357 ();
 sg13g2_decap_8 FILLER_1_3364 ();
 sg13g2_decap_8 FILLER_1_3371 ();
 sg13g2_decap_8 FILLER_1_3378 ();
 sg13g2_decap_8 FILLER_1_3385 ();
 sg13g2_decap_8 FILLER_1_3392 ();
 sg13g2_decap_8 FILLER_1_3399 ();
 sg13g2_decap_8 FILLER_1_3406 ();
 sg13g2_decap_8 FILLER_1_3413 ();
 sg13g2_decap_8 FILLER_1_3420 ();
 sg13g2_decap_8 FILLER_1_3427 ();
 sg13g2_decap_8 FILLER_1_3434 ();
 sg13g2_decap_8 FILLER_1_3441 ();
 sg13g2_decap_8 FILLER_1_3448 ();
 sg13g2_decap_8 FILLER_1_3455 ();
 sg13g2_decap_8 FILLER_1_3462 ();
 sg13g2_decap_8 FILLER_1_3469 ();
 sg13g2_decap_8 FILLER_1_3476 ();
 sg13g2_decap_8 FILLER_1_3483 ();
 sg13g2_decap_8 FILLER_1_3490 ();
 sg13g2_decap_8 FILLER_1_3497 ();
 sg13g2_decap_8 FILLER_1_3504 ();
 sg13g2_decap_8 FILLER_1_3511 ();
 sg13g2_decap_8 FILLER_1_3518 ();
 sg13g2_decap_8 FILLER_1_3525 ();
 sg13g2_decap_8 FILLER_1_3532 ();
 sg13g2_decap_8 FILLER_1_3539 ();
 sg13g2_decap_8 FILLER_1_3546 ();
 sg13g2_decap_8 FILLER_1_3553 ();
 sg13g2_decap_8 FILLER_1_3560 ();
 sg13g2_decap_8 FILLER_1_3567 ();
 sg13g2_decap_4 FILLER_1_3574 ();
 sg13g2_fill_2 FILLER_1_3578 ();
 sg13g2_decap_4 FILLER_2_0 ();
 sg13g2_fill_2 FILLER_2_48 ();
 sg13g2_fill_1 FILLER_2_50 ();
 sg13g2_fill_2 FILLER_2_87 ();
 sg13g2_decap_8 FILLER_2_131 ();
 sg13g2_decap_4 FILLER_2_138 ();
 sg13g2_fill_2 FILLER_2_142 ();
 sg13g2_fill_2 FILLER_2_179 ();
 sg13g2_fill_1 FILLER_2_181 ();
 sg13g2_fill_1 FILLER_2_201 ();
 sg13g2_decap_8 FILLER_2_234 ();
 sg13g2_fill_2 FILLER_2_289 ();
 sg13g2_fill_1 FILLER_2_291 ();
 sg13g2_fill_2 FILLER_2_302 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_fill_2 FILLER_2_357 ();
 sg13g2_fill_1 FILLER_2_363 ();
 sg13g2_fill_2 FILLER_2_373 ();
 sg13g2_fill_1 FILLER_2_375 ();
 sg13g2_fill_2 FILLER_2_397 ();
 sg13g2_decap_8 FILLER_2_425 ();
 sg13g2_fill_2 FILLER_2_462 ();
 sg13g2_fill_1 FILLER_2_464 ();
 sg13g2_fill_2 FILLER_2_495 ();
 sg13g2_fill_2 FILLER_2_502 ();
 sg13g2_fill_2 FILLER_2_544 ();
 sg13g2_fill_1 FILLER_2_555 ();
 sg13g2_fill_2 FILLER_2_565 ();
 sg13g2_fill_2 FILLER_2_598 ();
 sg13g2_fill_1 FILLER_2_600 ();
 sg13g2_decap_8 FILLER_2_624 ();
 sg13g2_decap_4 FILLER_2_631 ();
 sg13g2_fill_2 FILLER_2_635 ();
 sg13g2_fill_1 FILLER_2_655 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_fill_1 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_677 ();
 sg13g2_decap_8 FILLER_2_684 ();
 sg13g2_decap_8 FILLER_2_722 ();
 sg13g2_fill_1 FILLER_2_729 ();
 sg13g2_decap_4 FILLER_2_756 ();
 sg13g2_fill_1 FILLER_2_760 ();
 sg13g2_fill_2 FILLER_2_774 ();
 sg13g2_fill_2 FILLER_2_780 ();
 sg13g2_fill_1 FILLER_2_782 ();
 sg13g2_decap_8 FILLER_2_797 ();
 sg13g2_fill_1 FILLER_2_804 ();
 sg13g2_fill_2 FILLER_2_809 ();
 sg13g2_fill_2 FILLER_2_825 ();
 sg13g2_fill_1 FILLER_2_836 ();
 sg13g2_decap_4 FILLER_2_841 ();
 sg13g2_fill_1 FILLER_2_845 ();
 sg13g2_decap_4 FILLER_2_864 ();
 sg13g2_decap_4 FILLER_2_881 ();
 sg13g2_fill_1 FILLER_2_885 ();
 sg13g2_fill_1 FILLER_2_891 ();
 sg13g2_decap_8 FILLER_2_896 ();
 sg13g2_decap_4 FILLER_2_912 ();
 sg13g2_fill_1 FILLER_2_916 ();
 sg13g2_fill_2 FILLER_2_926 ();
 sg13g2_fill_1 FILLER_2_928 ();
 sg13g2_decap_8 FILLER_2_942 ();
 sg13g2_fill_2 FILLER_2_949 ();
 sg13g2_fill_1 FILLER_2_951 ();
 sg13g2_fill_1 FILLER_2_957 ();
 sg13g2_decap_4 FILLER_2_962 ();
 sg13g2_fill_2 FILLER_2_980 ();
 sg13g2_fill_2 FILLER_2_990 ();
 sg13g2_fill_1 FILLER_2_992 ();
 sg13g2_fill_2 FILLER_2_998 ();
 sg13g2_fill_1 FILLER_2_1000 ();
 sg13g2_fill_1 FILLER_2_1032 ();
 sg13g2_fill_1 FILLER_2_1086 ();
 sg13g2_fill_2 FILLER_2_1132 ();
 sg13g2_fill_2 FILLER_2_1139 ();
 sg13g2_decap_8 FILLER_2_1145 ();
 sg13g2_decap_4 FILLER_2_1152 ();
 sg13g2_fill_1 FILLER_2_1187 ();
 sg13g2_fill_2 FILLER_2_1196 ();
 sg13g2_fill_1 FILLER_2_1198 ();
 sg13g2_decap_8 FILLER_2_1211 ();
 sg13g2_fill_2 FILLER_2_1226 ();
 sg13g2_fill_1 FILLER_2_1237 ();
 sg13g2_decap_4 FILLER_2_1243 ();
 sg13g2_fill_2 FILLER_2_1255 ();
 sg13g2_fill_1 FILLER_2_1257 ();
 sg13g2_fill_1 FILLER_2_1271 ();
 sg13g2_decap_8 FILLER_2_1276 ();
 sg13g2_fill_2 FILLER_2_1283 ();
 sg13g2_decap_8 FILLER_2_1353 ();
 sg13g2_fill_1 FILLER_2_1360 ();
 sg13g2_decap_4 FILLER_2_1365 ();
 sg13g2_fill_1 FILLER_2_1369 ();
 sg13g2_decap_8 FILLER_2_1387 ();
 sg13g2_fill_2 FILLER_2_1394 ();
 sg13g2_decap_4 FILLER_2_1431 ();
 sg13g2_fill_1 FILLER_2_1435 ();
 sg13g2_fill_1 FILLER_2_1441 ();
 sg13g2_decap_8 FILLER_2_1477 ();
 sg13g2_decap_8 FILLER_2_1484 ();
 sg13g2_fill_1 FILLER_2_1491 ();
 sg13g2_fill_1 FILLER_2_1518 ();
 sg13g2_fill_1 FILLER_2_1524 ();
 sg13g2_decap_4 FILLER_2_1529 ();
 sg13g2_fill_2 FILLER_2_1533 ();
 sg13g2_decap_8 FILLER_2_1542 ();
 sg13g2_fill_1 FILLER_2_1549 ();
 sg13g2_decap_8 FILLER_2_1554 ();
 sg13g2_fill_2 FILLER_2_1561 ();
 sg13g2_fill_1 FILLER_2_1563 ();
 sg13g2_fill_2 FILLER_2_1609 ();
 sg13g2_fill_1 FILLER_2_1633 ();
 sg13g2_fill_1 FILLER_2_1643 ();
 sg13g2_decap_4 FILLER_2_1695 ();
 sg13g2_fill_1 FILLER_2_1699 ();
 sg13g2_decap_4 FILLER_2_1704 ();
 sg13g2_fill_1 FILLER_2_1708 ();
 sg13g2_decap_8 FILLER_2_1722 ();
 sg13g2_fill_2 FILLER_2_1729 ();
 sg13g2_decap_4 FILLER_2_1735 ();
 sg13g2_fill_2 FILLER_2_1739 ();
 sg13g2_decap_8 FILLER_2_1758 ();
 sg13g2_fill_2 FILLER_2_1765 ();
 sg13g2_decap_8 FILLER_2_1776 ();
 sg13g2_decap_4 FILLER_2_1783 ();
 sg13g2_fill_2 FILLER_2_1787 ();
 sg13g2_decap_8 FILLER_2_1794 ();
 sg13g2_fill_1 FILLER_2_1801 ();
 sg13g2_decap_4 FILLER_2_1837 ();
 sg13g2_fill_1 FILLER_2_1841 ();
 sg13g2_decap_8 FILLER_2_1887 ();
 sg13g2_decap_4 FILLER_2_1894 ();
 sg13g2_fill_2 FILLER_2_1903 ();
 sg13g2_decap_8 FILLER_2_1909 ();
 sg13g2_decap_4 FILLER_2_1916 ();
 sg13g2_decap_4 FILLER_2_1946 ();
 sg13g2_decap_8 FILLER_2_1954 ();
 sg13g2_fill_1 FILLER_2_1974 ();
 sg13g2_fill_2 FILLER_2_1988 ();
 sg13g2_decap_4 FILLER_2_2026 ();
 sg13g2_decap_8 FILLER_2_2096 ();
 sg13g2_decap_4 FILLER_2_2103 ();
 sg13g2_decap_8 FILLER_2_2116 ();
 sg13g2_fill_2 FILLER_2_2123 ();
 sg13g2_decap_4 FILLER_2_2129 ();
 sg13g2_fill_2 FILLER_2_2142 ();
 sg13g2_fill_1 FILLER_2_2144 ();
 sg13g2_decap_8 FILLER_2_2176 ();
 sg13g2_decap_8 FILLER_2_2183 ();
 sg13g2_fill_2 FILLER_2_2204 ();
 sg13g2_fill_2 FILLER_2_2215 ();
 sg13g2_fill_1 FILLER_2_2217 ();
 sg13g2_fill_2 FILLER_2_2240 ();
 sg13g2_fill_1 FILLER_2_2242 ();
 sg13g2_fill_1 FILLER_2_2273 ();
 sg13g2_fill_2 FILLER_2_2302 ();
 sg13g2_decap_8 FILLER_2_2335 ();
 sg13g2_decap_4 FILLER_2_2342 ();
 sg13g2_fill_1 FILLER_2_2346 ();
 sg13g2_decap_4 FILLER_2_2351 ();
 sg13g2_fill_2 FILLER_2_2373 ();
 sg13g2_decap_8 FILLER_2_2392 ();
 sg13g2_decap_8 FILLER_2_2408 ();
 sg13g2_decap_8 FILLER_2_2415 ();
 sg13g2_fill_2 FILLER_2_2422 ();
 sg13g2_fill_1 FILLER_2_2429 ();
 sg13g2_fill_2 FILLER_2_2439 ();
 sg13g2_fill_2 FILLER_2_2450 ();
 sg13g2_fill_1 FILLER_2_2452 ();
 sg13g2_fill_2 FILLER_2_2462 ();
 sg13g2_fill_1 FILLER_2_2464 ();
 sg13g2_fill_2 FILLER_2_2479 ();
 sg13g2_fill_1 FILLER_2_2481 ();
 sg13g2_fill_2 FILLER_2_2490 ();
 sg13g2_fill_1 FILLER_2_2492 ();
 sg13g2_decap_8 FILLER_2_2498 ();
 sg13g2_decap_4 FILLER_2_2505 ();
 sg13g2_fill_1 FILLER_2_2509 ();
 sg13g2_fill_1 FILLER_2_2515 ();
 sg13g2_fill_2 FILLER_2_2520 ();
 sg13g2_fill_1 FILLER_2_2522 ();
 sg13g2_decap_8 FILLER_2_2527 ();
 sg13g2_decap_4 FILLER_2_2534 ();
 sg13g2_fill_1 FILLER_2_2538 ();
 sg13g2_decap_8 FILLER_2_2588 ();
 sg13g2_decap_4 FILLER_2_2595 ();
 sg13g2_fill_2 FILLER_2_2609 ();
 sg13g2_fill_1 FILLER_2_2611 ();
 sg13g2_decap_4 FILLER_2_2616 ();
 sg13g2_fill_1 FILLER_2_2620 ();
 sg13g2_fill_2 FILLER_2_2639 ();
 sg13g2_fill_1 FILLER_2_2641 ();
 sg13g2_fill_2 FILLER_2_2647 ();
 sg13g2_decap_8 FILLER_2_2654 ();
 sg13g2_decap_8 FILLER_2_2661 ();
 sg13g2_decap_4 FILLER_2_2668 ();
 sg13g2_fill_2 FILLER_2_2703 ();
 sg13g2_fill_1 FILLER_2_2705 ();
 sg13g2_fill_2 FILLER_2_2710 ();
 sg13g2_fill_1 FILLER_2_2712 ();
 sg13g2_fill_1 FILLER_2_2735 ();
 sg13g2_fill_2 FILLER_2_2750 ();
 sg13g2_decap_8 FILLER_2_2778 ();
 sg13g2_fill_2 FILLER_2_2785 ();
 sg13g2_fill_2 FILLER_2_2796 ();
 sg13g2_fill_1 FILLER_2_2811 ();
 sg13g2_fill_2 FILLER_2_2821 ();
 sg13g2_fill_1 FILLER_2_2823 ();
 sg13g2_decap_8 FILLER_2_2850 ();
 sg13g2_decap_8 FILLER_2_2857 ();
 sg13g2_fill_2 FILLER_2_2864 ();
 sg13g2_fill_1 FILLER_2_2866 ();
 sg13g2_decap_8 FILLER_2_2871 ();
 sg13g2_decap_4 FILLER_2_2878 ();
 sg13g2_decap_8 FILLER_2_2887 ();
 sg13g2_fill_1 FILLER_2_2894 ();
 sg13g2_decap_4 FILLER_2_2899 ();
 sg13g2_decap_8 FILLER_2_2921 ();
 sg13g2_decap_8 FILLER_2_2928 ();
 sg13g2_decap_4 FILLER_2_2935 ();
 sg13g2_decap_8 FILLER_2_2973 ();
 sg13g2_decap_4 FILLER_2_2980 ();
 sg13g2_fill_2 FILLER_2_2984 ();
 sg13g2_decap_8 FILLER_2_2991 ();
 sg13g2_fill_1 FILLER_2_3024 ();
 sg13g2_decap_8 FILLER_2_3051 ();
 sg13g2_decap_8 FILLER_2_3058 ();
 sg13g2_decap_8 FILLER_2_3065 ();
 sg13g2_decap_8 FILLER_2_3072 ();
 sg13g2_decap_8 FILLER_2_3079 ();
 sg13g2_decap_8 FILLER_2_3086 ();
 sg13g2_decap_8 FILLER_2_3093 ();
 sg13g2_decap_8 FILLER_2_3100 ();
 sg13g2_decap_8 FILLER_2_3107 ();
 sg13g2_decap_8 FILLER_2_3114 ();
 sg13g2_decap_8 FILLER_2_3121 ();
 sg13g2_decap_8 FILLER_2_3128 ();
 sg13g2_decap_8 FILLER_2_3135 ();
 sg13g2_decap_8 FILLER_2_3142 ();
 sg13g2_fill_2 FILLER_2_3149 ();
 sg13g2_fill_2 FILLER_2_3155 ();
 sg13g2_fill_1 FILLER_2_3161 ();
 sg13g2_decap_8 FILLER_2_3171 ();
 sg13g2_decap_8 FILLER_2_3178 ();
 sg13g2_decap_8 FILLER_2_3185 ();
 sg13g2_decap_8 FILLER_2_3192 ();
 sg13g2_decap_8 FILLER_2_3199 ();
 sg13g2_decap_8 FILLER_2_3206 ();
 sg13g2_decap_8 FILLER_2_3213 ();
 sg13g2_fill_2 FILLER_2_3220 ();
 sg13g2_decap_8 FILLER_2_3227 ();
 sg13g2_decap_8 FILLER_2_3234 ();
 sg13g2_decap_4 FILLER_2_3241 ();
 sg13g2_fill_1 FILLER_2_3245 ();
 sg13g2_decap_8 FILLER_2_3250 ();
 sg13g2_decap_8 FILLER_2_3257 ();
 sg13g2_decap_8 FILLER_2_3264 ();
 sg13g2_decap_8 FILLER_2_3271 ();
 sg13g2_decap_8 FILLER_2_3278 ();
 sg13g2_decap_8 FILLER_2_3285 ();
 sg13g2_decap_8 FILLER_2_3292 ();
 sg13g2_fill_2 FILLER_2_3299 ();
 sg13g2_decap_8 FILLER_2_3306 ();
 sg13g2_decap_8 FILLER_2_3313 ();
 sg13g2_decap_8 FILLER_2_3320 ();
 sg13g2_decap_8 FILLER_2_3327 ();
 sg13g2_decap_8 FILLER_2_3334 ();
 sg13g2_decap_8 FILLER_2_3341 ();
 sg13g2_decap_8 FILLER_2_3348 ();
 sg13g2_decap_8 FILLER_2_3355 ();
 sg13g2_decap_8 FILLER_2_3362 ();
 sg13g2_decap_8 FILLER_2_3369 ();
 sg13g2_decap_8 FILLER_2_3376 ();
 sg13g2_decap_8 FILLER_2_3383 ();
 sg13g2_decap_8 FILLER_2_3390 ();
 sg13g2_decap_8 FILLER_2_3397 ();
 sg13g2_decap_8 FILLER_2_3404 ();
 sg13g2_decap_8 FILLER_2_3411 ();
 sg13g2_decap_8 FILLER_2_3418 ();
 sg13g2_decap_8 FILLER_2_3425 ();
 sg13g2_decap_8 FILLER_2_3432 ();
 sg13g2_decap_8 FILLER_2_3439 ();
 sg13g2_decap_8 FILLER_2_3446 ();
 sg13g2_decap_8 FILLER_2_3453 ();
 sg13g2_decap_8 FILLER_2_3460 ();
 sg13g2_decap_8 FILLER_2_3467 ();
 sg13g2_decap_8 FILLER_2_3474 ();
 sg13g2_decap_8 FILLER_2_3481 ();
 sg13g2_decap_8 FILLER_2_3488 ();
 sg13g2_decap_8 FILLER_2_3495 ();
 sg13g2_decap_8 FILLER_2_3502 ();
 sg13g2_decap_8 FILLER_2_3509 ();
 sg13g2_decap_8 FILLER_2_3516 ();
 sg13g2_decap_8 FILLER_2_3523 ();
 sg13g2_decap_8 FILLER_2_3530 ();
 sg13g2_decap_8 FILLER_2_3537 ();
 sg13g2_decap_8 FILLER_2_3544 ();
 sg13g2_decap_8 FILLER_2_3551 ();
 sg13g2_decap_8 FILLER_2_3558 ();
 sg13g2_decap_8 FILLER_2_3565 ();
 sg13g2_decap_8 FILLER_2_3572 ();
 sg13g2_fill_1 FILLER_2_3579 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_fill_1 FILLER_3_31 ();
 sg13g2_decap_8 FILLER_3_62 ();
 sg13g2_fill_2 FILLER_3_69 ();
 sg13g2_fill_1 FILLER_3_71 ();
 sg13g2_decap_8 FILLER_3_76 ();
 sg13g2_decap_4 FILLER_3_83 ();
 sg13g2_fill_1 FILLER_3_87 ();
 sg13g2_fill_1 FILLER_3_102 ();
 sg13g2_decap_4 FILLER_3_122 ();
 sg13g2_fill_2 FILLER_3_136 ();
 sg13g2_fill_1 FILLER_3_138 ();
 sg13g2_fill_2 FILLER_3_166 ();
 sg13g2_fill_1 FILLER_3_168 ();
 sg13g2_fill_2 FILLER_3_267 ();
 sg13g2_fill_2 FILLER_3_279 ();
 sg13g2_fill_1 FILLER_3_290 ();
 sg13g2_fill_2 FILLER_3_346 ();
 sg13g2_decap_8 FILLER_3_393 ();
 sg13g2_fill_2 FILLER_3_400 ();
 sg13g2_decap_4 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_423 ();
 sg13g2_fill_2 FILLER_3_440 ();
 sg13g2_fill_2 FILLER_3_480 ();
 sg13g2_fill_2 FILLER_3_621 ();
 sg13g2_decap_4 FILLER_3_679 ();
 sg13g2_fill_1 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_723 ();
 sg13g2_fill_2 FILLER_3_739 ();
 sg13g2_fill_1 FILLER_3_858 ();
 sg13g2_fill_2 FILLER_3_885 ();
 sg13g2_fill_2 FILLER_3_913 ();
 sg13g2_fill_1 FILLER_3_915 ();
 sg13g2_fill_2 FILLER_3_994 ();
 sg13g2_fill_1 FILLER_3_996 ();
 sg13g2_decap_4 FILLER_3_1005 ();
 sg13g2_decap_8 FILLER_3_1030 ();
 sg13g2_fill_1 FILLER_3_1037 ();
 sg13g2_fill_2 FILLER_3_1043 ();
 sg13g2_fill_1 FILLER_3_1045 ();
 sg13g2_fill_2 FILLER_3_1050 ();
 sg13g2_fill_1 FILLER_3_1052 ();
 sg13g2_decap_8 FILLER_3_1057 ();
 sg13g2_fill_2 FILLER_3_1064 ();
 sg13g2_fill_1 FILLER_3_1066 ();
 sg13g2_decap_4 FILLER_3_1102 ();
 sg13g2_fill_2 FILLER_3_1106 ();
 sg13g2_fill_2 FILLER_3_1116 ();
 sg13g2_fill_2 FILLER_3_1127 ();
 sg13g2_fill_1 FILLER_3_1129 ();
 sg13g2_decap_8 FILLER_3_1156 ();
 sg13g2_decap_8 FILLER_3_1163 ();
 sg13g2_fill_2 FILLER_3_1170 ();
 sg13g2_fill_2 FILLER_3_1180 ();
 sg13g2_fill_1 FILLER_3_1191 ();
 sg13g2_fill_2 FILLER_3_1201 ();
 sg13g2_decap_8 FILLER_3_1234 ();
 sg13g2_fill_1 FILLER_3_1241 ();
 sg13g2_decap_4 FILLER_3_1282 ();
 sg13g2_fill_2 FILLER_3_1286 ();
 sg13g2_decap_8 FILLER_3_1292 ();
 sg13g2_fill_1 FILLER_3_1339 ();
 sg13g2_fill_2 FILLER_3_1352 ();
 sg13g2_fill_1 FILLER_3_1354 ();
 sg13g2_fill_2 FILLER_3_1386 ();
 sg13g2_fill_1 FILLER_3_1388 ();
 sg13g2_decap_8 FILLER_3_1397 ();
 sg13g2_fill_2 FILLER_3_1404 ();
 sg13g2_fill_1 FILLER_3_1406 ();
 sg13g2_decap_8 FILLER_3_1442 ();
 sg13g2_fill_2 FILLER_3_1449 ();
 sg13g2_fill_1 FILLER_3_1451 ();
 sg13g2_fill_2 FILLER_3_1456 ();
 sg13g2_fill_1 FILLER_3_1476 ();
 sg13g2_decap_8 FILLER_3_1485 ();
 sg13g2_fill_1 FILLER_3_1492 ();
 sg13g2_decap_4 FILLER_3_1498 ();
 sg13g2_fill_2 FILLER_3_1510 ();
 sg13g2_fill_1 FILLER_3_1512 ();
 sg13g2_fill_2 FILLER_3_1522 ();
 sg13g2_decap_4 FILLER_3_1559 ();
 sg13g2_fill_1 FILLER_3_1563 ();
 sg13g2_decap_4 FILLER_3_1569 ();
 sg13g2_fill_2 FILLER_3_1578 ();
 sg13g2_decap_8 FILLER_3_1592 ();
 sg13g2_fill_2 FILLER_3_1599 ();
 sg13g2_fill_1 FILLER_3_1658 ();
 sg13g2_fill_2 FILLER_3_1681 ();
 sg13g2_fill_1 FILLER_3_1683 ();
 sg13g2_fill_2 FILLER_3_1719 ();
 sg13g2_fill_2 FILLER_3_1761 ();
 sg13g2_fill_2 FILLER_3_1815 ();
 sg13g2_decap_4 FILLER_3_1821 ();
 sg13g2_fill_2 FILLER_3_1851 ();
 sg13g2_fill_1 FILLER_3_1853 ();
 sg13g2_fill_2 FILLER_3_1867 ();
 sg13g2_fill_1 FILLER_3_1878 ();
 sg13g2_fill_2 FILLER_3_1944 ();
 sg13g2_fill_1 FILLER_3_1972 ();
 sg13g2_fill_2 FILLER_3_2094 ();
 sg13g2_decap_8 FILLER_3_2122 ();
 sg13g2_decap_4 FILLER_3_2129 ();
 sg13g2_fill_1 FILLER_3_2147 ();
 sg13g2_fill_1 FILLER_3_2161 ();
 sg13g2_decap_8 FILLER_3_2167 ();
 sg13g2_fill_1 FILLER_3_2174 ();
 sg13g2_fill_1 FILLER_3_2235 ();
 sg13g2_fill_2 FILLER_3_2272 ();
 sg13g2_fill_1 FILLER_3_2274 ();
 sg13g2_decap_8 FILLER_3_2301 ();
 sg13g2_fill_2 FILLER_3_2308 ();
 sg13g2_fill_1 FILLER_3_2310 ();
 sg13g2_fill_1 FILLER_3_2319 ();
 sg13g2_fill_2 FILLER_3_2328 ();
 sg13g2_fill_1 FILLER_3_2330 ();
 sg13g2_fill_1 FILLER_3_2357 ();
 sg13g2_fill_2 FILLER_3_2632 ();
 sg13g2_fill_1 FILLER_3_2634 ();
 sg13g2_decap_8 FILLER_3_2661 ();
 sg13g2_decap_8 FILLER_3_2668 ();
 sg13g2_fill_1 FILLER_3_2683 ();
 sg13g2_fill_2 FILLER_3_2701 ();
 sg13g2_fill_1 FILLER_3_2703 ();
 sg13g2_fill_2 FILLER_3_2735 ();
 sg13g2_fill_2 FILLER_3_2742 ();
 sg13g2_fill_1 FILLER_3_2744 ();
 sg13g2_decap_4 FILLER_3_2760 ();
 sg13g2_fill_2 FILLER_3_2764 ();
 sg13g2_fill_1 FILLER_3_2823 ();
 sg13g2_decap_4 FILLER_3_2829 ();
 sg13g2_fill_2 FILLER_3_2833 ();
 sg13g2_decap_8 FILLER_3_2839 ();
 sg13g2_decap_4 FILLER_3_2846 ();
 sg13g2_fill_2 FILLER_3_2850 ();
 sg13g2_fill_2 FILLER_3_2882 ();
 sg13g2_fill_2 FILLER_3_2910 ();
 sg13g2_decap_4 FILLER_3_2938 ();
 sg13g2_decap_8 FILLER_3_3048 ();
 sg13g2_decap_8 FILLER_3_3055 ();
 sg13g2_decap_8 FILLER_3_3062 ();
 sg13g2_decap_8 FILLER_3_3069 ();
 sg13g2_decap_8 FILLER_3_3076 ();
 sg13g2_decap_8 FILLER_3_3083 ();
 sg13g2_decap_8 FILLER_3_3090 ();
 sg13g2_decap_8 FILLER_3_3097 ();
 sg13g2_decap_8 FILLER_3_3104 ();
 sg13g2_decap_8 FILLER_3_3111 ();
 sg13g2_decap_8 FILLER_3_3118 ();
 sg13g2_fill_2 FILLER_3_3125 ();
 sg13g2_fill_1 FILLER_3_3127 ();
 sg13g2_decap_8 FILLER_3_3132 ();
 sg13g2_decap_8 FILLER_3_3139 ();
 sg13g2_decap_8 FILLER_3_3172 ();
 sg13g2_decap_8 FILLER_3_3179 ();
 sg13g2_decap_8 FILLER_3_3186 ();
 sg13g2_decap_8 FILLER_3_3193 ();
 sg13g2_decap_8 FILLER_3_3200 ();
 sg13g2_decap_8 FILLER_3_3207 ();
 sg13g2_decap_4 FILLER_3_3214 ();
 sg13g2_fill_1 FILLER_3_3218 ();
 sg13g2_fill_2 FILLER_3_3271 ();
 sg13g2_fill_1 FILLER_3_3273 ();
 sg13g2_fill_2 FILLER_3_3300 ();
 sg13g2_decap_8 FILLER_3_3328 ();
 sg13g2_decap_8 FILLER_3_3335 ();
 sg13g2_decap_8 FILLER_3_3342 ();
 sg13g2_decap_8 FILLER_3_3349 ();
 sg13g2_decap_8 FILLER_3_3356 ();
 sg13g2_decap_8 FILLER_3_3363 ();
 sg13g2_fill_2 FILLER_3_3370 ();
 sg13g2_decap_4 FILLER_3_3398 ();
 sg13g2_decap_8 FILLER_3_3428 ();
 sg13g2_decap_8 FILLER_3_3435 ();
 sg13g2_decap_8 FILLER_3_3442 ();
 sg13g2_decap_8 FILLER_3_3454 ();
 sg13g2_decap_4 FILLER_3_3461 ();
 sg13g2_decap_8 FILLER_3_3469 ();
 sg13g2_decap_8 FILLER_3_3476 ();
 sg13g2_decap_8 FILLER_3_3483 ();
 sg13g2_decap_8 FILLER_3_3490 ();
 sg13g2_decap_8 FILLER_3_3497 ();
 sg13g2_decap_8 FILLER_3_3504 ();
 sg13g2_decap_8 FILLER_3_3511 ();
 sg13g2_fill_2 FILLER_3_3518 ();
 sg13g2_decap_8 FILLER_3_3524 ();
 sg13g2_decap_8 FILLER_3_3531 ();
 sg13g2_decap_8 FILLER_3_3538 ();
 sg13g2_decap_8 FILLER_3_3545 ();
 sg13g2_decap_8 FILLER_3_3552 ();
 sg13g2_decap_8 FILLER_3_3559 ();
 sg13g2_decap_8 FILLER_3_3566 ();
 sg13g2_decap_8 FILLER_3_3573 ();
 sg13g2_decap_4 FILLER_4_0 ();
 sg13g2_fill_1 FILLER_4_4 ();
 sg13g2_fill_1 FILLER_4_31 ();
 sg13g2_decap_4 FILLER_4_55 ();
 sg13g2_fill_1 FILLER_4_59 ();
 sg13g2_decap_4 FILLER_4_90 ();
 sg13g2_fill_1 FILLER_4_120 ();
 sg13g2_fill_1 FILLER_4_126 ();
 sg13g2_fill_2 FILLER_4_132 ();
 sg13g2_fill_1 FILLER_4_179 ();
 sg13g2_decap_8 FILLER_4_193 ();
 sg13g2_fill_2 FILLER_4_213 ();
 sg13g2_fill_2 FILLER_4_257 ();
 sg13g2_fill_1 FILLER_4_259 ();
 sg13g2_fill_1 FILLER_4_278 ();
 sg13g2_decap_8 FILLER_4_284 ();
 sg13g2_decap_4 FILLER_4_291 ();
 sg13g2_fill_2 FILLER_4_295 ();
 sg13g2_decap_8 FILLER_4_346 ();
 sg13g2_decap_8 FILLER_4_353 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_fill_1 FILLER_4_371 ();
 sg13g2_decap_4 FILLER_4_398 ();
 sg13g2_fill_2 FILLER_4_402 ();
 sg13g2_fill_2 FILLER_4_409 ();
 sg13g2_fill_1 FILLER_4_411 ();
 sg13g2_fill_2 FILLER_4_438 ();
 sg13g2_fill_2 FILLER_4_487 ();
 sg13g2_decap_4 FILLER_4_495 ();
 sg13g2_decap_4 FILLER_4_525 ();
 sg13g2_fill_1 FILLER_4_529 ();
 sg13g2_fill_2 FILLER_4_538 ();
 sg13g2_fill_1 FILLER_4_545 ();
 sg13g2_decap_4 FILLER_4_549 ();
 sg13g2_fill_2 FILLER_4_566 ();
 sg13g2_fill_1 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_586 ();
 sg13g2_decap_8 FILLER_4_593 ();
 sg13g2_decap_4 FILLER_4_600 ();
 sg13g2_fill_2 FILLER_4_604 ();
 sg13g2_fill_2 FILLER_4_610 ();
 sg13g2_fill_1 FILLER_4_612 ();
 sg13g2_fill_2 FILLER_4_626 ();
 sg13g2_fill_1 FILLER_4_628 ();
 sg13g2_fill_2 FILLER_4_673 ();
 sg13g2_fill_2 FILLER_4_710 ();
 sg13g2_decap_8 FILLER_4_716 ();
 sg13g2_fill_1 FILLER_4_767 ();
 sg13g2_fill_1 FILLER_4_785 ();
 sg13g2_fill_2 FILLER_4_790 ();
 sg13g2_fill_1 FILLER_4_792 ();
 sg13g2_decap_4 FILLER_4_806 ();
 sg13g2_fill_2 FILLER_4_810 ();
 sg13g2_decap_4 FILLER_4_820 ();
 sg13g2_decap_8 FILLER_4_838 ();
 sg13g2_fill_2 FILLER_4_866 ();
 sg13g2_fill_2 FILLER_4_875 ();
 sg13g2_decap_4 FILLER_4_889 ();
 sg13g2_fill_1 FILLER_4_897 ();
 sg13g2_decap_4 FILLER_4_902 ();
 sg13g2_fill_1 FILLER_4_906 ();
 sg13g2_decap_8 FILLER_4_912 ();
 sg13g2_decap_4 FILLER_4_919 ();
 sg13g2_fill_2 FILLER_4_923 ();
 sg13g2_fill_1 FILLER_4_933 ();
 sg13g2_fill_2 FILLER_4_943 ();
 sg13g2_fill_2 FILLER_4_958 ();
 sg13g2_fill_2 FILLER_4_969 ();
 sg13g2_decap_4 FILLER_4_1030 ();
 sg13g2_fill_1 FILLER_4_1034 ();
 sg13g2_fill_2 FILLER_4_1061 ();
 sg13g2_decap_8 FILLER_4_1068 ();
 sg13g2_fill_2 FILLER_4_1075 ();
 sg13g2_fill_1 FILLER_4_1077 ();
 sg13g2_decap_4 FILLER_4_1103 ();
 sg13g2_decap_8 FILLER_4_1117 ();
 sg13g2_fill_1 FILLER_4_1124 ();
 sg13g2_decap_8 FILLER_4_1147 ();
 sg13g2_decap_8 FILLER_4_1159 ();
 sg13g2_decap_4 FILLER_4_1170 ();
 sg13g2_decap_8 FILLER_4_1240 ();
 sg13g2_fill_2 FILLER_4_1247 ();
 sg13g2_fill_2 FILLER_4_1275 ();
 sg13g2_decap_8 FILLER_4_1303 ();
 sg13g2_fill_1 FILLER_4_1310 ();
 sg13g2_fill_2 FILLER_4_1333 ();
 sg13g2_fill_1 FILLER_4_1340 ();
 sg13g2_fill_2 FILLER_4_1367 ();
 sg13g2_fill_1 FILLER_4_1369 ();
 sg13g2_decap_8 FILLER_4_1396 ();
 sg13g2_fill_2 FILLER_4_1416 ();
 sg13g2_decap_4 FILLER_4_1439 ();
 sg13g2_fill_2 FILLER_4_1443 ();
 sg13g2_fill_1 FILLER_4_1471 ();
 sg13g2_decap_4 FILLER_4_1477 ();
 sg13g2_fill_1 FILLER_4_1481 ();
 sg13g2_decap_8 FILLER_4_1494 ();
 sg13g2_decap_4 FILLER_4_1501 ();
 sg13g2_fill_1 FILLER_4_1505 ();
 sg13g2_fill_2 FILLER_4_1536 ();
 sg13g2_fill_1 FILLER_4_1538 ();
 sg13g2_decap_8 FILLER_4_1599 ();
 sg13g2_decap_4 FILLER_4_1606 ();
 sg13g2_decap_8 FILLER_4_1618 ();
 sg13g2_decap_4 FILLER_4_1625 ();
 sg13g2_fill_2 FILLER_4_1633 ();
 sg13g2_fill_1 FILLER_4_1635 ();
 sg13g2_decap_8 FILLER_4_1684 ();
 sg13g2_decap_8 FILLER_4_1691 ();
 sg13g2_fill_2 FILLER_4_1720 ();
 sg13g2_fill_1 FILLER_4_1722 ();
 sg13g2_fill_2 FILLER_4_1732 ();
 sg13g2_decap_4 FILLER_4_1739 ();
 sg13g2_fill_2 FILLER_4_1769 ();
 sg13g2_fill_2 FILLER_4_1789 ();
 sg13g2_decap_4 FILLER_4_1795 ();
 sg13g2_fill_2 FILLER_4_1817 ();
 sg13g2_fill_2 FILLER_4_1837 ();
 sg13g2_fill_2 FILLER_4_1852 ();
 sg13g2_fill_1 FILLER_4_1854 ();
 sg13g2_fill_2 FILLER_4_1859 ();
 sg13g2_fill_2 FILLER_4_1887 ();
 sg13g2_fill_1 FILLER_4_1889 ();
 sg13g2_fill_1 FILLER_4_1894 ();
 sg13g2_fill_2 FILLER_4_1908 ();
 sg13g2_fill_2 FILLER_4_1914 ();
 sg13g2_fill_2 FILLER_4_1939 ();
 sg13g2_fill_1 FILLER_4_1950 ();
 sg13g2_decap_8 FILLER_4_1964 ();
 sg13g2_decap_8 FILLER_4_1975 ();
 sg13g2_decap_4 FILLER_4_1982 ();
 sg13g2_decap_4 FILLER_4_1999 ();
 sg13g2_fill_1 FILLER_4_2003 ();
 sg13g2_decap_4 FILLER_4_2017 ();
 sg13g2_fill_1 FILLER_4_2021 ();
 sg13g2_decap_8 FILLER_4_2035 ();
 sg13g2_decap_8 FILLER_4_2042 ();
 sg13g2_fill_2 FILLER_4_2087 ();
 sg13g2_fill_1 FILLER_4_2089 ();
 sg13g2_fill_2 FILLER_4_2095 ();
 sg13g2_fill_1 FILLER_4_2102 ();
 sg13g2_fill_2 FILLER_4_2177 ();
 sg13g2_fill_1 FILLER_4_2192 ();
 sg13g2_fill_1 FILLER_4_2206 ();
 sg13g2_fill_1 FILLER_4_2211 ();
 sg13g2_fill_2 FILLER_4_2225 ();
 sg13g2_decap_8 FILLER_4_2267 ();
 sg13g2_fill_1 FILLER_4_2274 ();
 sg13g2_fill_1 FILLER_4_2279 ();
 sg13g2_fill_2 FILLER_4_2297 ();
 sg13g2_fill_1 FILLER_4_2299 ();
 sg13g2_decap_8 FILLER_4_2326 ();
 sg13g2_fill_2 FILLER_4_2333 ();
 sg13g2_fill_1 FILLER_4_2340 ();
 sg13g2_fill_1 FILLER_4_2345 ();
 sg13g2_decap_4 FILLER_4_2380 ();
 sg13g2_fill_2 FILLER_4_2384 ();
 sg13g2_fill_2 FILLER_4_2395 ();
 sg13g2_fill_2 FILLER_4_2401 ();
 sg13g2_fill_1 FILLER_4_2403 ();
 sg13g2_decap_4 FILLER_4_2413 ();
 sg13g2_fill_2 FILLER_4_2417 ();
 sg13g2_fill_2 FILLER_4_2433 ();
 sg13g2_decap_8 FILLER_4_2444 ();
 sg13g2_fill_2 FILLER_4_2455 ();
 sg13g2_fill_2 FILLER_4_2461 ();
 sg13g2_fill_1 FILLER_4_2481 ();
 sg13g2_decap_4 FILLER_4_2491 ();
 sg13g2_fill_1 FILLER_4_2499 ();
 sg13g2_fill_2 FILLER_4_2521 ();
 sg13g2_fill_1 FILLER_4_2541 ();
 sg13g2_fill_1 FILLER_4_2594 ();
 sg13g2_decap_4 FILLER_4_2608 ();
 sg13g2_fill_2 FILLER_4_2651 ();
 sg13g2_decap_4 FILLER_4_2670 ();
 sg13g2_fill_2 FILLER_4_2674 ();
 sg13g2_fill_1 FILLER_4_2684 ();
 sg13g2_fill_2 FILLER_4_2716 ();
 sg13g2_fill_2 FILLER_4_2731 ();
 sg13g2_fill_1 FILLER_4_2733 ();
 sg13g2_fill_2 FILLER_4_2760 ();
 sg13g2_fill_1 FILLER_4_2762 ();
 sg13g2_decap_4 FILLER_4_2772 ();
 sg13g2_fill_1 FILLER_4_2776 ();
 sg13g2_decap_4 FILLER_4_2790 ();
 sg13g2_fill_1 FILLER_4_2794 ();
 sg13g2_fill_2 FILLER_4_2817 ();
 sg13g2_fill_1 FILLER_4_2819 ();
 sg13g2_decap_8 FILLER_4_2855 ();
 sg13g2_fill_2 FILLER_4_2862 ();
 sg13g2_decap_4 FILLER_4_2899 ();
 sg13g2_decap_8 FILLER_4_2908 ();
 sg13g2_fill_2 FILLER_4_2915 ();
 sg13g2_fill_1 FILLER_4_2917 ();
 sg13g2_fill_1 FILLER_4_2922 ();
 sg13g2_fill_2 FILLER_4_2927 ();
 sg13g2_fill_1 FILLER_4_2947 ();
 sg13g2_decap_8 FILLER_4_2979 ();
 sg13g2_fill_2 FILLER_4_2986 ();
 sg13g2_fill_1 FILLER_4_2988 ();
 sg13g2_fill_1 FILLER_4_2993 ();
 sg13g2_fill_2 FILLER_4_2998 ();
 sg13g2_decap_8 FILLER_4_3066 ();
 sg13g2_decap_8 FILLER_4_3073 ();
 sg13g2_decap_8 FILLER_4_3080 ();
 sg13g2_decap_8 FILLER_4_3087 ();
 sg13g2_decap_8 FILLER_4_3094 ();
 sg13g2_decap_8 FILLER_4_3101 ();
 sg13g2_decap_8 FILLER_4_3108 ();
 sg13g2_fill_2 FILLER_4_3115 ();
 sg13g2_fill_1 FILLER_4_3117 ();
 sg13g2_decap_8 FILLER_4_3144 ();
 sg13g2_fill_1 FILLER_4_3181 ();
 sg13g2_decap_8 FILLER_4_3208 ();
 sg13g2_decap_8 FILLER_4_3215 ();
 sg13g2_fill_2 FILLER_4_3222 ();
 sg13g2_fill_1 FILLER_4_3224 ();
 sg13g2_fill_1 FILLER_4_3229 ();
 sg13g2_fill_2 FILLER_4_3234 ();
 sg13g2_fill_1 FILLER_4_3250 ();
 sg13g2_fill_2 FILLER_4_3256 ();
 sg13g2_fill_1 FILLER_4_3258 ();
 sg13g2_fill_1 FILLER_4_3272 ();
 sg13g2_fill_2 FILLER_4_3282 ();
 sg13g2_fill_1 FILLER_4_3284 ();
 sg13g2_fill_1 FILLER_4_3289 ();
 sg13g2_decap_4 FILLER_4_3299 ();
 sg13g2_fill_2 FILLER_4_3303 ();
 sg13g2_decap_4 FILLER_4_3309 ();
 sg13g2_decap_4 FILLER_4_3326 ();
 sg13g2_fill_2 FILLER_4_3330 ();
 sg13g2_decap_4 FILLER_4_3358 ();
 sg13g2_fill_1 FILLER_4_3362 ();
 sg13g2_fill_1 FILLER_4_3393 ();
 sg13g2_fill_1 FILLER_4_3412 ();
 sg13g2_decap_8 FILLER_4_3430 ();
 sg13g2_fill_2 FILLER_4_3437 ();
 sg13g2_fill_2 FILLER_4_3443 ();
 sg13g2_decap_4 FILLER_4_3450 ();
 sg13g2_decap_8 FILLER_4_3536 ();
 sg13g2_decap_8 FILLER_4_3543 ();
 sg13g2_decap_8 FILLER_4_3550 ();
 sg13g2_decap_8 FILLER_4_3557 ();
 sg13g2_decap_8 FILLER_4_3564 ();
 sg13g2_decap_8 FILLER_4_3571 ();
 sg13g2_fill_2 FILLER_4_3578 ();
 sg13g2_decap_4 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_4 ();
 sg13g2_fill_1 FILLER_5_50 ();
 sg13g2_fill_1 FILLER_5_82 ();
 sg13g2_decap_4 FILLER_5_96 ();
 sg13g2_fill_1 FILLER_5_104 ();
 sg13g2_decap_8 FILLER_5_109 ();
 sg13g2_decap_4 FILLER_5_116 ();
 sg13g2_fill_1 FILLER_5_120 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_4 FILLER_5_154 ();
 sg13g2_fill_2 FILLER_5_158 ();
 sg13g2_fill_1 FILLER_5_196 ();
 sg13g2_decap_4 FILLER_5_220 ();
 sg13g2_fill_2 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_241 ();
 sg13g2_fill_2 FILLER_5_274 ();
 sg13g2_fill_1 FILLER_5_322 ();
 sg13g2_fill_2 FILLER_5_380 ();
 sg13g2_fill_1 FILLER_5_382 ();
 sg13g2_fill_2 FILLER_5_422 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_fill_2 FILLER_5_448 ();
 sg13g2_fill_1 FILLER_5_450 ();
 sg13g2_decap_4 FILLER_5_461 ();
 sg13g2_fill_2 FILLER_5_465 ();
 sg13g2_decap_4 FILLER_5_473 ();
 sg13g2_fill_2 FILLER_5_477 ();
 sg13g2_decap_4 FILLER_5_505 ();
 sg13g2_fill_1 FILLER_5_509 ();
 sg13g2_decap_4 FILLER_5_531 ();
 sg13g2_fill_1 FILLER_5_535 ();
 sg13g2_decap_4 FILLER_5_592 ();
 sg13g2_fill_2 FILLER_5_609 ();
 sg13g2_fill_1 FILLER_5_611 ();
 sg13g2_fill_2 FILLER_5_638 ();
 sg13g2_fill_1 FILLER_5_666 ();
 sg13g2_decap_8 FILLER_5_689 ();
 sg13g2_decap_8 FILLER_5_727 ();
 sg13g2_decap_4 FILLER_5_738 ();
 sg13g2_fill_1 FILLER_5_750 ();
 sg13g2_decap_4 FILLER_5_761 ();
 sg13g2_fill_2 FILLER_5_804 ();
 sg13g2_fill_1 FILLER_5_806 ();
 sg13g2_fill_2 FILLER_5_833 ();
 sg13g2_fill_1 FILLER_5_835 ();
 sg13g2_fill_1 FILLER_5_858 ();
 sg13g2_fill_1 FILLER_5_888 ();
 sg13g2_fill_2 FILLER_5_935 ();
 sg13g2_fill_2 FILLER_5_942 ();
 sg13g2_decap_8 FILLER_5_956 ();
 sg13g2_fill_1 FILLER_5_963 ();
 sg13g2_fill_2 FILLER_5_969 ();
 sg13g2_fill_2 FILLER_5_976 ();
 sg13g2_decap_8 FILLER_5_999 ();
 sg13g2_decap_8 FILLER_5_1006 ();
 sg13g2_decap_4 FILLER_5_1013 ();
 sg13g2_fill_2 FILLER_5_1017 ();
 sg13g2_fill_2 FILLER_5_1045 ();
 sg13g2_fill_1 FILLER_5_1067 ();
 sg13g2_fill_1 FILLER_5_1073 ();
 sg13g2_fill_1 FILLER_5_1094 ();
 sg13g2_fill_1 FILLER_5_1105 ();
 sg13g2_fill_2 FILLER_5_1127 ();
 sg13g2_decap_8 FILLER_5_1181 ();
 sg13g2_decap_8 FILLER_5_1188 ();
 sg13g2_decap_4 FILLER_5_1195 ();
 sg13g2_fill_2 FILLER_5_1213 ();
 sg13g2_fill_1 FILLER_5_1215 ();
 sg13g2_fill_2 FILLER_5_1252 ();
 sg13g2_fill_2 FILLER_5_1266 ();
 sg13g2_fill_1 FILLER_5_1282 ();
 sg13g2_decap_8 FILLER_5_1302 ();
 sg13g2_decap_4 FILLER_5_1309 ();
 sg13g2_decap_4 FILLER_5_1339 ();
 sg13g2_fill_1 FILLER_5_1343 ();
 sg13g2_fill_2 FILLER_5_1349 ();
 sg13g2_fill_1 FILLER_5_1351 ();
 sg13g2_fill_2 FILLER_5_1373 ();
 sg13g2_fill_1 FILLER_5_1397 ();
 sg13g2_decap_8 FILLER_5_1429 ();
 sg13g2_fill_2 FILLER_5_1436 ();
 sg13g2_decap_4 FILLER_5_1443 ();
 sg13g2_fill_1 FILLER_5_1447 ();
 sg13g2_fill_2 FILLER_5_1452 ();
 sg13g2_fill_1 FILLER_5_1476 ();
 sg13g2_decap_4 FILLER_5_1503 ();
 sg13g2_fill_2 FILLER_5_1521 ();
 sg13g2_fill_2 FILLER_5_1546 ();
 sg13g2_fill_2 FILLER_5_1558 ();
 sg13g2_fill_1 FILLER_5_1573 ();
 sg13g2_decap_4 FILLER_5_1596 ();
 sg13g2_fill_2 FILLER_5_1647 ();
 sg13g2_fill_2 FILLER_5_1653 ();
 sg13g2_fill_1 FILLER_5_1660 ();
 sg13g2_decap_8 FILLER_5_1665 ();
 sg13g2_fill_2 FILLER_5_1672 ();
 sg13g2_fill_1 FILLER_5_1674 ();
 sg13g2_decap_8 FILLER_5_1680 ();
 sg13g2_decap_8 FILLER_5_1687 ();
 sg13g2_decap_4 FILLER_5_1694 ();
 sg13g2_fill_1 FILLER_5_1729 ();
 sg13g2_fill_2 FILLER_5_1756 ();
 sg13g2_fill_2 FILLER_5_1762 ();
 sg13g2_decap_8 FILLER_5_1782 ();
 sg13g2_fill_2 FILLER_5_1789 ();
 sg13g2_decap_8 FILLER_5_1799 ();
 sg13g2_decap_8 FILLER_5_1806 ();
 sg13g2_decap_4 FILLER_5_1844 ();
 sg13g2_fill_2 FILLER_5_1848 ();
 sg13g2_decap_4 FILLER_5_1881 ();
 sg13g2_fill_2 FILLER_5_1891 ();
 sg13g2_fill_1 FILLER_5_1893 ();
 sg13g2_fill_1 FILLER_5_1903 ();
 sg13g2_decap_8 FILLER_5_1914 ();
 sg13g2_decap_4 FILLER_5_1921 ();
 sg13g2_fill_2 FILLER_5_1986 ();
 sg13g2_fill_1 FILLER_5_1988 ();
 sg13g2_decap_8 FILLER_5_2019 ();
 sg13g2_fill_2 FILLER_5_2030 ();
 sg13g2_fill_1 FILLER_5_2063 ();
 sg13g2_fill_2 FILLER_5_2089 ();
 sg13g2_fill_2 FILLER_5_2134 ();
 sg13g2_decap_8 FILLER_5_2145 ();
 sg13g2_fill_1 FILLER_5_2161 ();
 sg13g2_fill_2 FILLER_5_2166 ();
 sg13g2_fill_1 FILLER_5_2172 ();
 sg13g2_decap_8 FILLER_5_2182 ();
 sg13g2_fill_2 FILLER_5_2189 ();
 sg13g2_decap_8 FILLER_5_2222 ();
 sg13g2_fill_2 FILLER_5_2229 ();
 sg13g2_fill_1 FILLER_5_2231 ();
 sg13g2_decap_4 FILLER_5_2236 ();
 sg13g2_fill_2 FILLER_5_2266 ();
 sg13g2_fill_1 FILLER_5_2268 ();
 sg13g2_fill_1 FILLER_5_2309 ();
 sg13g2_fill_1 FILLER_5_2345 ();
 sg13g2_decap_4 FILLER_5_2377 ();
 sg13g2_fill_2 FILLER_5_2381 ();
 sg13g2_fill_2 FILLER_5_2392 ();
 sg13g2_fill_1 FILLER_5_2394 ();
 sg13g2_decap_8 FILLER_5_2421 ();
 sg13g2_decap_4 FILLER_5_2428 ();
 sg13g2_fill_1 FILLER_5_2432 ();
 sg13g2_decap_4 FILLER_5_2437 ();
 sg13g2_decap_8 FILLER_5_2470 ();
 sg13g2_decap_8 FILLER_5_2503 ();
 sg13g2_decap_4 FILLER_5_2510 ();
 sg13g2_decap_8 FILLER_5_2545 ();
 sg13g2_decap_8 FILLER_5_2552 ();
 sg13g2_decap_8 FILLER_5_2559 ();
 sg13g2_fill_2 FILLER_5_2566 ();
 sg13g2_fill_1 FILLER_5_2568 ();
 sg13g2_fill_1 FILLER_5_2574 ();
 sg13g2_fill_1 FILLER_5_2583 ();
 sg13g2_decap_4 FILLER_5_2589 ();
 sg13g2_fill_2 FILLER_5_2593 ();
 sg13g2_fill_2 FILLER_5_2600 ();
 sg13g2_fill_1 FILLER_5_2644 ();
 sg13g2_fill_1 FILLER_5_2671 ();
 sg13g2_fill_2 FILLER_5_2698 ();
 sg13g2_fill_1 FILLER_5_2700 ();
 sg13g2_decap_4 FILLER_5_2749 ();
 sg13g2_fill_1 FILLER_5_2819 ();
 sg13g2_fill_1 FILLER_5_2824 ();
 sg13g2_fill_1 FILLER_5_2834 ();
 sg13g2_decap_4 FILLER_5_2861 ();
 sg13g2_fill_2 FILLER_5_2873 ();
 sg13g2_decap_4 FILLER_5_2953 ();
 sg13g2_fill_2 FILLER_5_2961 ();
 sg13g2_fill_1 FILLER_5_2963 ();
 sg13g2_fill_2 FILLER_5_2977 ();
 sg13g2_fill_2 FILLER_5_3010 ();
 sg13g2_fill_1 FILLER_5_3012 ();
 sg13g2_fill_2 FILLER_5_3022 ();
 sg13g2_fill_1 FILLER_5_3024 ();
 sg13g2_fill_1 FILLER_5_3051 ();
 sg13g2_fill_1 FILLER_5_3066 ();
 sg13g2_fill_2 FILLER_5_3093 ();
 sg13g2_fill_1 FILLER_5_3135 ();
 sg13g2_decap_8 FILLER_5_3145 ();
 sg13g2_fill_2 FILLER_5_3152 ();
 sg13g2_fill_2 FILLER_5_3168 ();
 sg13g2_fill_1 FILLER_5_3170 ();
 sg13g2_fill_2 FILLER_5_3180 ();
 sg13g2_fill_1 FILLER_5_3182 ();
 sg13g2_fill_2 FILLER_5_3223 ();
 sg13g2_fill_1 FILLER_5_3225 ();
 sg13g2_fill_2 FILLER_5_3236 ();
 sg13g2_fill_1 FILLER_5_3238 ();
 sg13g2_decap_8 FILLER_5_3265 ();
 sg13g2_decap_4 FILLER_5_3272 ();
 sg13g2_fill_1 FILLER_5_3281 ();
 sg13g2_decap_8 FILLER_5_3290 ();
 sg13g2_decap_4 FILLER_5_3297 ();
 sg13g2_fill_1 FILLER_5_3301 ();
 sg13g2_decap_8 FILLER_5_3328 ();
 sg13g2_fill_2 FILLER_5_3335 ();
 sg13g2_fill_2 FILLER_5_3369 ();
 sg13g2_fill_2 FILLER_5_3380 ();
 sg13g2_fill_1 FILLER_5_3382 ();
 sg13g2_decap_8 FILLER_5_3418 ();
 sg13g2_decap_4 FILLER_5_3425 ();
 sg13g2_fill_2 FILLER_5_3455 ();
 sg13g2_fill_1 FILLER_5_3457 ();
 sg13g2_decap_8 FILLER_5_3462 ();
 sg13g2_fill_1 FILLER_5_3469 ();
 sg13g2_fill_1 FILLER_5_3492 ();
 sg13g2_fill_1 FILLER_5_3506 ();
 sg13g2_fill_1 FILLER_5_3516 ();
 sg13g2_fill_2 FILLER_5_3526 ();
 sg13g2_fill_2 FILLER_5_3537 ();
 sg13g2_decap_8 FILLER_5_3544 ();
 sg13g2_decap_8 FILLER_5_3555 ();
 sg13g2_decap_8 FILLER_5_3562 ();
 sg13g2_decap_8 FILLER_5_3569 ();
 sg13g2_decap_4 FILLER_5_3576 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_fill_2 FILLER_6_15 ();
 sg13g2_fill_1 FILLER_6_17 ();
 sg13g2_fill_1 FILLER_6_61 ();
 sg13g2_fill_1 FILLER_6_70 ();
 sg13g2_decap_4 FILLER_6_81 ();
 sg13g2_fill_2 FILLER_6_100 ();
 sg13g2_fill_2 FILLER_6_111 ();
 sg13g2_fill_2 FILLER_6_140 ();
 sg13g2_decap_4 FILLER_6_158 ();
 sg13g2_fill_1 FILLER_6_162 ();
 sg13g2_fill_2 FILLER_6_178 ();
 sg13g2_fill_1 FILLER_6_180 ();
 sg13g2_decap_4 FILLER_6_230 ();
 sg13g2_fill_2 FILLER_6_234 ();
 sg13g2_fill_2 FILLER_6_320 ();
 sg13g2_fill_1 FILLER_6_388 ();
 sg13g2_decap_4 FILLER_6_406 ();
 sg13g2_fill_2 FILLER_6_436 ();
 sg13g2_fill_1 FILLER_6_447 ();
 sg13g2_fill_1 FILLER_6_468 ();
 sg13g2_decap_8 FILLER_6_478 ();
 sg13g2_fill_1 FILLER_6_485 ();
 sg13g2_fill_2 FILLER_6_490 ();
 sg13g2_fill_2 FILLER_6_509 ();
 sg13g2_decap_8 FILLER_6_524 ();
 sg13g2_decap_4 FILLER_6_531 ();
 sg13g2_fill_2 FILLER_6_535 ();
 sg13g2_decap_8 FILLER_6_550 ();
 sg13g2_decap_8 FILLER_6_557 ();
 sg13g2_fill_2 FILLER_6_564 ();
 sg13g2_fill_2 FILLER_6_571 ();
 sg13g2_fill_2 FILLER_6_577 ();
 sg13g2_fill_1 FILLER_6_579 ();
 sg13g2_decap_8 FILLER_6_611 ();
 sg13g2_fill_1 FILLER_6_623 ();
 sg13g2_decap_8 FILLER_6_632 ();
 sg13g2_decap_4 FILLER_6_639 ();
 sg13g2_fill_1 FILLER_6_643 ();
 sg13g2_fill_2 FILLER_6_648 ();
 sg13g2_fill_1 FILLER_6_654 ();
 sg13g2_fill_1 FILLER_6_664 ();
 sg13g2_decap_8 FILLER_6_691 ();
 sg13g2_decap_4 FILLER_6_698 ();
 sg13g2_fill_2 FILLER_6_702 ();
 sg13g2_fill_2 FILLER_6_715 ();
 sg13g2_decap_8 FILLER_6_729 ();
 sg13g2_fill_1 FILLER_6_736 ();
 sg13g2_decap_8 FILLER_6_762 ();
 sg13g2_decap_8 FILLER_6_769 ();
 sg13g2_decap_8 FILLER_6_776 ();
 sg13g2_fill_2 FILLER_6_783 ();
 sg13g2_fill_1 FILLER_6_785 ();
 sg13g2_decap_8 FILLER_6_796 ();
 sg13g2_decap_4 FILLER_6_803 ();
 sg13g2_fill_2 FILLER_6_807 ();
 sg13g2_fill_2 FILLER_6_817 ();
 sg13g2_fill_2 FILLER_6_824 ();
 sg13g2_fill_2 FILLER_6_836 ();
 sg13g2_fill_1 FILLER_6_838 ();
 sg13g2_fill_2 FILLER_6_864 ();
 sg13g2_decap_8 FILLER_6_886 ();
 sg13g2_fill_2 FILLER_6_893 ();
 sg13g2_fill_1 FILLER_6_895 ();
 sg13g2_decap_8 FILLER_6_904 ();
 sg13g2_decap_4 FILLER_6_911 ();
 sg13g2_decap_4 FILLER_6_932 ();
 sg13g2_fill_2 FILLER_6_944 ();
 sg13g2_fill_1 FILLER_6_951 ();
 sg13g2_fill_2 FILLER_6_982 ();
 sg13g2_fill_1 FILLER_6_984 ();
 sg13g2_decap_8 FILLER_6_994 ();
 sg13g2_fill_2 FILLER_6_1001 ();
 sg13g2_fill_1 FILLER_6_1003 ();
 sg13g2_fill_1 FILLER_6_1020 ();
 sg13g2_decap_8 FILLER_6_1047 ();
 sg13g2_fill_2 FILLER_6_1075 ();
 sg13g2_decap_8 FILLER_6_1082 ();
 sg13g2_decap_8 FILLER_6_1102 ();
 sg13g2_decap_8 FILLER_6_1109 ();
 sg13g2_decap_4 FILLER_6_1116 ();
 sg13g2_fill_2 FILLER_6_1120 ();
 sg13g2_fill_2 FILLER_6_1126 ();
 sg13g2_fill_2 FILLER_6_1146 ();
 sg13g2_fill_2 FILLER_6_1178 ();
 sg13g2_decap_8 FILLER_6_1230 ();
 sg13g2_decap_8 FILLER_6_1237 ();
 sg13g2_decap_4 FILLER_6_1244 ();
 sg13g2_fill_1 FILLER_6_1278 ();
 sg13g2_decap_4 FILLER_6_1318 ();
 sg13g2_fill_2 FILLER_6_1322 ();
 sg13g2_decap_4 FILLER_6_1328 ();
 sg13g2_fill_1 FILLER_6_1363 ();
 sg13g2_fill_1 FILLER_6_1369 ();
 sg13g2_decap_8 FILLER_6_1386 ();
 sg13g2_decap_8 FILLER_6_1393 ();
 sg13g2_fill_2 FILLER_6_1400 ();
 sg13g2_fill_1 FILLER_6_1402 ();
 sg13g2_decap_4 FILLER_6_1407 ();
 sg13g2_fill_2 FILLER_6_1426 ();
 sg13g2_decap_8 FILLER_6_1471 ();
 sg13g2_decap_4 FILLER_6_1478 ();
 sg13g2_fill_2 FILLER_6_1496 ();
 sg13g2_fill_1 FILLER_6_1529 ();
 sg13g2_fill_1 FILLER_6_1551 ();
 sg13g2_decap_4 FILLER_6_1569 ();
 sg13g2_fill_1 FILLER_6_1573 ();
 sg13g2_fill_2 FILLER_6_1587 ();
 sg13g2_fill_1 FILLER_6_1611 ();
 sg13g2_fill_1 FILLER_6_1647 ();
 sg13g2_decap_4 FILLER_6_1700 ();
 sg13g2_fill_2 FILLER_6_1704 ();
 sg13g2_decap_4 FILLER_6_1711 ();
 sg13g2_fill_2 FILLER_6_1715 ();
 sg13g2_decap_8 FILLER_6_1726 ();
 sg13g2_decap_8 FILLER_6_1733 ();
 sg13g2_fill_1 FILLER_6_1740 ();
 sg13g2_fill_1 FILLER_6_1745 ();
 sg13g2_fill_2 FILLER_6_1750 ();
 sg13g2_fill_1 FILLER_6_1761 ();
 sg13g2_fill_1 FILLER_6_1783 ();
 sg13g2_fill_2 FILLER_6_1810 ();
 sg13g2_decap_8 FILLER_6_1833 ();
 sg13g2_fill_2 FILLER_6_1840 ();
 sg13g2_fill_1 FILLER_6_1842 ();
 sg13g2_fill_2 FILLER_6_1899 ();
 sg13g2_decap_8 FILLER_6_1922 ();
 sg13g2_decap_4 FILLER_6_1929 ();
 sg13g2_fill_2 FILLER_6_1933 ();
 sg13g2_fill_2 FILLER_6_1947 ();
 sg13g2_decap_8 FILLER_6_1970 ();
 sg13g2_decap_8 FILLER_6_1977 ();
 sg13g2_fill_2 FILLER_6_1984 ();
 sg13g2_fill_1 FILLER_6_1999 ();
 sg13g2_decap_4 FILLER_6_2004 ();
 sg13g2_fill_2 FILLER_6_2008 ();
 sg13g2_fill_2 FILLER_6_2049 ();
 sg13g2_decap_8 FILLER_6_2073 ();
 sg13g2_fill_1 FILLER_6_2085 ();
 sg13g2_decap_4 FILLER_6_2090 ();
 sg13g2_fill_2 FILLER_6_2107 ();
 sg13g2_decap_8 FILLER_6_2119 ();
 sg13g2_fill_2 FILLER_6_2156 ();
 sg13g2_fill_1 FILLER_6_2158 ();
 sg13g2_decap_8 FILLER_6_2206 ();
 sg13g2_fill_2 FILLER_6_2213 ();
 sg13g2_fill_1 FILLER_6_2215 ();
 sg13g2_fill_1 FILLER_6_2281 ();
 sg13g2_decap_8 FILLER_6_2290 ();
 sg13g2_fill_2 FILLER_6_2297 ();
 sg13g2_fill_1 FILLER_6_2299 ();
 sg13g2_fill_2 FILLER_6_2320 ();
 sg13g2_fill_1 FILLER_6_2322 ();
 sg13g2_decap_4 FILLER_6_2341 ();
 sg13g2_fill_1 FILLER_6_2345 ();
 sg13g2_decap_8 FILLER_6_2356 ();
 sg13g2_decap_4 FILLER_6_2363 ();
 sg13g2_fill_2 FILLER_6_2367 ();
 sg13g2_fill_1 FILLER_6_2382 ();
 sg13g2_decap_4 FILLER_6_2396 ();
 sg13g2_fill_1 FILLER_6_2400 ();
 sg13g2_decap_8 FILLER_6_2436 ();
 sg13g2_fill_1 FILLER_6_2443 ();
 sg13g2_fill_2 FILLER_6_2457 ();
 sg13g2_fill_1 FILLER_6_2468 ();
 sg13g2_decap_4 FILLER_6_2526 ();
 sg13g2_decap_8 FILLER_6_2534 ();
 sg13g2_fill_1 FILLER_6_2541 ();
 sg13g2_fill_1 FILLER_6_2568 ();
 sg13g2_decap_8 FILLER_6_2620 ();
 sg13g2_decap_4 FILLER_6_2627 ();
 sg13g2_decap_4 FILLER_6_2636 ();
 sg13g2_fill_1 FILLER_6_2640 ();
 sg13g2_fill_1 FILLER_6_2646 ();
 sg13g2_fill_2 FILLER_6_2660 ();
 sg13g2_fill_1 FILLER_6_2662 ();
 sg13g2_decap_8 FILLER_6_2672 ();
 sg13g2_fill_2 FILLER_6_2679 ();
 sg13g2_fill_1 FILLER_6_2681 ();
 sg13g2_fill_2 FILLER_6_2686 ();
 sg13g2_decap_8 FILLER_6_2704 ();
 sg13g2_fill_2 FILLER_6_2711 ();
 sg13g2_fill_1 FILLER_6_2713 ();
 sg13g2_decap_4 FILLER_6_2752 ();
 sg13g2_fill_1 FILLER_6_2756 ();
 sg13g2_fill_2 FILLER_6_2770 ();
 sg13g2_fill_1 FILLER_6_2772 ();
 sg13g2_decap_4 FILLER_6_2786 ();
 sg13g2_decap_8 FILLER_6_2793 ();
 sg13g2_decap_4 FILLER_6_2800 ();
 sg13g2_decap_8 FILLER_6_2816 ();
 sg13g2_decap_4 FILLER_6_2828 ();
 sg13g2_decap_8 FILLER_6_2866 ();
 sg13g2_decap_8 FILLER_6_2873 ();
 sg13g2_fill_2 FILLER_6_2880 ();
 sg13g2_fill_1 FILLER_6_2882 ();
 sg13g2_decap_4 FILLER_6_2887 ();
 sg13g2_fill_1 FILLER_6_2891 ();
 sg13g2_decap_4 FILLER_6_2902 ();
 sg13g2_fill_1 FILLER_6_2906 ();
 sg13g2_fill_2 FILLER_6_2911 ();
 sg13g2_fill_1 FILLER_6_2917 ();
 sg13g2_fill_1 FILLER_6_2927 ();
 sg13g2_fill_2 FILLER_6_2951 ();
 sg13g2_fill_2 FILLER_6_2979 ();
 sg13g2_fill_2 FILLER_6_2999 ();
 sg13g2_decap_8 FILLER_6_3036 ();
 sg13g2_fill_1 FILLER_6_3043 ();
 sg13g2_decap_4 FILLER_6_3074 ();
 sg13g2_decap_8 FILLER_6_3091 ();
 sg13g2_decap_4 FILLER_6_3098 ();
 sg13g2_fill_1 FILLER_6_3107 ();
 sg13g2_fill_2 FILLER_6_3112 ();
 sg13g2_fill_1 FILLER_6_3114 ();
 sg13g2_fill_2 FILLER_6_3124 ();
 sg13g2_decap_4 FILLER_6_3152 ();
 sg13g2_fill_2 FILLER_6_3182 ();
 sg13g2_decap_4 FILLER_6_3189 ();
 sg13g2_fill_2 FILLER_6_3197 ();
 sg13g2_fill_2 FILLER_6_3212 ();
 sg13g2_decap_4 FILLER_6_3223 ();
 sg13g2_decap_4 FILLER_6_3257 ();
 sg13g2_fill_2 FILLER_6_3261 ();
 sg13g2_fill_1 FILLER_6_3268 ();
 sg13g2_fill_2 FILLER_6_3332 ();
 sg13g2_decap_4 FILLER_6_3360 ();
 sg13g2_fill_1 FILLER_6_3364 ();
 sg13g2_decap_8 FILLER_6_3373 ();
 sg13g2_fill_2 FILLER_6_3384 ();
 sg13g2_fill_1 FILLER_6_3386 ();
 sg13g2_fill_2 FILLER_6_3391 ();
 sg13g2_fill_1 FILLER_6_3402 ();
 sg13g2_fill_2 FILLER_6_3407 ();
 sg13g2_fill_2 FILLER_6_3426 ();
 sg13g2_fill_1 FILLER_6_3428 ();
 sg13g2_decap_8 FILLER_6_3452 ();
 sg13g2_decap_4 FILLER_6_3459 ();
 sg13g2_fill_1 FILLER_6_3463 ();
 sg13g2_decap_4 FILLER_6_3472 ();
 sg13g2_fill_1 FILLER_6_3476 ();
 sg13g2_decap_4 FILLER_6_3498 ();
 sg13g2_fill_2 FILLER_6_3510 ();
 sg13g2_fill_1 FILLER_6_3512 ();
 sg13g2_fill_2 FILLER_6_3539 ();
 sg13g2_decap_8 FILLER_6_3567 ();
 sg13g2_decap_4 FILLER_6_3574 ();
 sg13g2_fill_2 FILLER_6_3578 ();
 sg13g2_decap_8 FILLER_7_26 ();
 sg13g2_fill_1 FILLER_7_33 ();
 sg13g2_fill_2 FILLER_7_60 ();
 sg13g2_fill_1 FILLER_7_88 ();
 sg13g2_decap_4 FILLER_7_115 ();
 sg13g2_decap_4 FILLER_7_143 ();
 sg13g2_fill_2 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_165 ();
 sg13g2_decap_4 FILLER_7_172 ();
 sg13g2_fill_2 FILLER_7_176 ();
 sg13g2_fill_1 FILLER_7_191 ();
 sg13g2_fill_2 FILLER_7_228 ();
 sg13g2_fill_1 FILLER_7_230 ();
 sg13g2_decap_8 FILLER_7_257 ();
 sg13g2_fill_2 FILLER_7_264 ();
 sg13g2_fill_1 FILLER_7_266 ();
 sg13g2_decap_4 FILLER_7_281 ();
 sg13g2_fill_1 FILLER_7_285 ();
 sg13g2_decap_8 FILLER_7_346 ();
 sg13g2_decap_4 FILLER_7_353 ();
 sg13g2_fill_1 FILLER_7_396 ();
 sg13g2_decap_8 FILLER_7_410 ();
 sg13g2_decap_4 FILLER_7_443 ();
 sg13g2_decap_4 FILLER_7_473 ();
 sg13g2_fill_1 FILLER_7_477 ();
 sg13g2_decap_4 FILLER_7_483 ();
 sg13g2_fill_1 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_517 ();
 sg13g2_decap_8 FILLER_7_593 ();
 sg13g2_decap_8 FILLER_7_600 ();
 sg13g2_fill_2 FILLER_7_607 ();
 sg13g2_fill_1 FILLER_7_609 ();
 sg13g2_decap_4 FILLER_7_656 ();
 sg13g2_decap_4 FILLER_7_665 ();
 sg13g2_fill_1 FILLER_7_669 ();
 sg13g2_fill_1 FILLER_7_726 ();
 sg13g2_decap_4 FILLER_7_745 ();
 sg13g2_decap_4 FILLER_7_759 ();
 sg13g2_fill_2 FILLER_7_763 ();
 sg13g2_fill_2 FILLER_7_785 ();
 sg13g2_decap_4 FILLER_7_802 ();
 sg13g2_decap_4 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_862 ();
 sg13g2_fill_2 FILLER_7_869 ();
 sg13g2_fill_2 FILLER_7_879 ();
 sg13g2_fill_1 FILLER_7_881 ();
 sg13g2_decap_8 FILLER_7_886 ();
 sg13g2_fill_1 FILLER_7_898 ();
 sg13g2_decap_4 FILLER_7_925 ();
 sg13g2_fill_2 FILLER_7_929 ();
 sg13g2_fill_1 FILLER_7_957 ();
 sg13g2_fill_2 FILLER_7_967 ();
 sg13g2_fill_2 FILLER_7_979 ();
 sg13g2_fill_2 FILLER_7_994 ();
 sg13g2_fill_2 FILLER_7_1000 ();
 sg13g2_fill_1 FILLER_7_1002 ();
 sg13g2_fill_2 FILLER_7_1011 ();
 sg13g2_fill_1 FILLER_7_1013 ();
 sg13g2_fill_1 FILLER_7_1019 ();
 sg13g2_decap_4 FILLER_7_1025 ();
 sg13g2_decap_8 FILLER_7_1037 ();
 sg13g2_decap_4 FILLER_7_1044 ();
 sg13g2_fill_2 FILLER_7_1058 ();
 sg13g2_fill_1 FILLER_7_1060 ();
 sg13g2_decap_4 FILLER_7_1069 ();
 sg13g2_decap_4 FILLER_7_1081 ();
 sg13g2_fill_1 FILLER_7_1085 ();
 sg13g2_fill_1 FILLER_7_1100 ();
 sg13g2_fill_1 FILLER_7_1140 ();
 sg13g2_fill_2 FILLER_7_1194 ();
 sg13g2_fill_1 FILLER_7_1196 ();
 sg13g2_decap_8 FILLER_7_1226 ();
 sg13g2_fill_2 FILLER_7_1233 ();
 sg13g2_decap_8 FILLER_7_1248 ();
 sg13g2_decap_8 FILLER_7_1255 ();
 sg13g2_decap_4 FILLER_7_1276 ();
 sg13g2_fill_1 FILLER_7_1280 ();
 sg13g2_decap_8 FILLER_7_1300 ();
 sg13g2_fill_2 FILLER_7_1307 ();
 sg13g2_fill_1 FILLER_7_1309 ();
 sg13g2_decap_8 FILLER_7_1315 ();
 sg13g2_decap_8 FILLER_7_1329 ();
 sg13g2_fill_2 FILLER_7_1336 ();
 sg13g2_fill_2 FILLER_7_1345 ();
 sg13g2_fill_1 FILLER_7_1347 ();
 sg13g2_fill_2 FILLER_7_1352 ();
 sg13g2_fill_1 FILLER_7_1354 ();
 sg13g2_decap_8 FILLER_7_1370 ();
 sg13g2_fill_1 FILLER_7_1377 ();
 sg13g2_fill_2 FILLER_7_1428 ();
 sg13g2_fill_1 FILLER_7_1430 ();
 sg13g2_fill_2 FILLER_7_1448 ();
 sg13g2_fill_1 FILLER_7_1450 ();
 sg13g2_decap_4 FILLER_7_1468 ();
 sg13g2_fill_2 FILLER_7_1472 ();
 sg13g2_decap_4 FILLER_7_1498 ();
 sg13g2_fill_1 FILLER_7_1502 ();
 sg13g2_fill_2 FILLER_7_1522 ();
 sg13g2_fill_1 FILLER_7_1529 ();
 sg13g2_fill_2 FILLER_7_1535 ();
 sg13g2_decap_4 FILLER_7_1557 ();
 sg13g2_fill_2 FILLER_7_1561 ();
 sg13g2_fill_2 FILLER_7_1571 ();
 sg13g2_fill_2 FILLER_7_1578 ();
 sg13g2_fill_2 FILLER_7_1593 ();
 sg13g2_fill_1 FILLER_7_1595 ();
 sg13g2_decap_8 FILLER_7_1632 ();
 sg13g2_decap_4 FILLER_7_1639 ();
 sg13g2_fill_1 FILLER_7_1643 ();
 sg13g2_decap_4 FILLER_7_1649 ();
 sg13g2_fill_1 FILLER_7_1657 ();
 sg13g2_fill_1 FILLER_7_1702 ();
 sg13g2_decap_4 FILLER_7_1747 ();
 sg13g2_fill_2 FILLER_7_1751 ();
 sg13g2_fill_2 FILLER_7_1759 ();
 sg13g2_fill_1 FILLER_7_1761 ();
 sg13g2_fill_1 FILLER_7_1767 ();
 sg13g2_decap_8 FILLER_7_1779 ();
 sg13g2_fill_1 FILLER_7_1786 ();
 sg13g2_fill_2 FILLER_7_1790 ();
 sg13g2_fill_1 FILLER_7_1792 ();
 sg13g2_fill_2 FILLER_7_1802 ();
 sg13g2_fill_2 FILLER_7_1807 ();
 sg13g2_fill_1 FILLER_7_1809 ();
 sg13g2_decap_8 FILLER_7_1841 ();
 sg13g2_decap_4 FILLER_7_1852 ();
 sg13g2_fill_2 FILLER_7_1856 ();
 sg13g2_decap_8 FILLER_7_1871 ();
 sg13g2_decap_4 FILLER_7_1878 ();
 sg13g2_fill_1 FILLER_7_1882 ();
 sg13g2_decap_4 FILLER_7_1893 ();
 sg13g2_fill_2 FILLER_7_1902 ();
 sg13g2_fill_1 FILLER_7_1904 ();
 sg13g2_decap_8 FILLER_7_1911 ();
 sg13g2_fill_2 FILLER_7_1927 ();
 sg13g2_fill_1 FILLER_7_1933 ();
 sg13g2_fill_1 FILLER_7_1943 ();
 sg13g2_decap_8 FILLER_7_1967 ();
 sg13g2_fill_2 FILLER_7_1974 ();
 sg13g2_decap_8 FILLER_7_2001 ();
 sg13g2_decap_8 FILLER_7_2008 ();
 sg13g2_decap_4 FILLER_7_2025 ();
 sg13g2_fill_2 FILLER_7_2043 ();
 sg13g2_fill_2 FILLER_7_2071 ();
 sg13g2_fill_1 FILLER_7_2073 ();
 sg13g2_decap_4 FILLER_7_2100 ();
 sg13g2_fill_2 FILLER_7_2104 ();
 sg13g2_decap_8 FILLER_7_2127 ();
 sg13g2_fill_2 FILLER_7_2134 ();
 sg13g2_fill_1 FILLER_7_2136 ();
 sg13g2_decap_8 FILLER_7_2141 ();
 sg13g2_decap_8 FILLER_7_2148 ();
 sg13g2_decap_4 FILLER_7_2175 ();
 sg13g2_fill_1 FILLER_7_2187 ();
 sg13g2_fill_2 FILLER_7_2193 ();
 sg13g2_fill_1 FILLER_7_2195 ();
 sg13g2_decap_8 FILLER_7_2199 ();
 sg13g2_decap_8 FILLER_7_2211 ();
 sg13g2_fill_1 FILLER_7_2218 ();
 sg13g2_decap_4 FILLER_7_2233 ();
 sg13g2_fill_1 FILLER_7_2242 ();
 sg13g2_decap_8 FILLER_7_2246 ();
 sg13g2_decap_4 FILLER_7_2253 ();
 sg13g2_fill_1 FILLER_7_2257 ();
 sg13g2_fill_2 FILLER_7_2279 ();
 sg13g2_fill_1 FILLER_7_2281 ();
 sg13g2_fill_2 FILLER_7_2303 ();
 sg13g2_fill_1 FILLER_7_2305 ();
 sg13g2_fill_2 FILLER_7_2336 ();
 sg13g2_fill_1 FILLER_7_2338 ();
 sg13g2_decap_8 FILLER_7_2364 ();
 sg13g2_decap_4 FILLER_7_2401 ();
 sg13g2_fill_1 FILLER_7_2405 ();
 sg13g2_decap_4 FILLER_7_2410 ();
 sg13g2_fill_2 FILLER_7_2428 ();
 sg13g2_decap_8 FILLER_7_2451 ();
 sg13g2_fill_2 FILLER_7_2458 ();
 sg13g2_decap_8 FILLER_7_2484 ();
 sg13g2_fill_1 FILLER_7_2491 ();
 sg13g2_decap_4 FILLER_7_2496 ();
 sg13g2_fill_1 FILLER_7_2500 ();
 sg13g2_fill_1 FILLER_7_2523 ();
 sg13g2_decap_8 FILLER_7_2534 ();
 sg13g2_fill_2 FILLER_7_2541 ();
 sg13g2_fill_1 FILLER_7_2543 ();
 sg13g2_fill_2 FILLER_7_2557 ();
 sg13g2_fill_2 FILLER_7_2568 ();
 sg13g2_decap_8 FILLER_7_2578 ();
 sg13g2_decap_4 FILLER_7_2585 ();
 sg13g2_fill_2 FILLER_7_2589 ();
 sg13g2_decap_8 FILLER_7_2596 ();
 sg13g2_decap_4 FILLER_7_2603 ();
 sg13g2_fill_2 FILLER_7_2607 ();
 sg13g2_decap_4 FILLER_7_2619 ();
 sg13g2_fill_1 FILLER_7_2647 ();
 sg13g2_fill_2 FILLER_7_2709 ();
 sg13g2_decap_4 FILLER_7_2732 ();
 sg13g2_decap_8 FILLER_7_2771 ();
 sg13g2_fill_2 FILLER_7_2778 ();
 sg13g2_decap_4 FILLER_7_2807 ();
 sg13g2_fill_2 FILLER_7_2837 ();
 sg13g2_decap_8 FILLER_7_2865 ();
 sg13g2_fill_2 FILLER_7_2898 ();
 sg13g2_fill_1 FILLER_7_2900 ();
 sg13g2_decap_8 FILLER_7_2914 ();
 sg13g2_fill_2 FILLER_7_2921 ();
 sg13g2_decap_8 FILLER_7_2957 ();
 sg13g2_decap_8 FILLER_7_2964 ();
 sg13g2_decap_8 FILLER_7_2971 ();
 sg13g2_decap_8 FILLER_7_2978 ();
 sg13g2_decap_8 FILLER_7_3011 ();
 sg13g2_fill_2 FILLER_7_3018 ();
 sg13g2_fill_1 FILLER_7_3020 ();
 sg13g2_fill_2 FILLER_7_3029 ();
 sg13g2_decap_8 FILLER_7_3040 ();
 sg13g2_fill_2 FILLER_7_3052 ();
 sg13g2_fill_1 FILLER_7_3062 ();
 sg13g2_decap_4 FILLER_7_3075 ();
 sg13g2_fill_2 FILLER_7_3105 ();
 sg13g2_fill_1 FILLER_7_3107 ();
 sg13g2_fill_2 FILLER_7_3142 ();
 sg13g2_fill_1 FILLER_7_3144 ();
 sg13g2_fill_1 FILLER_7_3158 ();
 sg13g2_decap_4 FILLER_7_3163 ();
 sg13g2_fill_1 FILLER_7_3180 ();
 sg13g2_fill_2 FILLER_7_3207 ();
 sg13g2_fill_1 FILLER_7_3221 ();
 sg13g2_fill_1 FILLER_7_3227 ();
 sg13g2_fill_1 FILLER_7_3236 ();
 sg13g2_decap_8 FILLER_7_3272 ();
 sg13g2_fill_2 FILLER_7_3279 ();
 sg13g2_fill_1 FILLER_7_3281 ();
 sg13g2_fill_1 FILLER_7_3296 ();
 sg13g2_fill_2 FILLER_7_3305 ();
 sg13g2_decap_8 FILLER_7_3338 ();
 sg13g2_fill_2 FILLER_7_3353 ();
 sg13g2_decap_4 FILLER_7_3399 ();
 sg13g2_fill_2 FILLER_7_3408 ();
 sg13g2_fill_1 FILLER_7_3410 ();
 sg13g2_decap_8 FILLER_7_3427 ();
 sg13g2_fill_2 FILLER_7_3434 ();
 sg13g2_fill_2 FILLER_7_3476 ();
 sg13g2_fill_1 FILLER_7_3478 ();
 sg13g2_decap_8 FILLER_7_3489 ();
 sg13g2_decap_8 FILLER_7_3496 ();
 sg13g2_decap_4 FILLER_7_3503 ();
 sg13g2_fill_2 FILLER_7_3507 ();
 sg13g2_fill_1 FILLER_7_3522 ();
 sg13g2_fill_1 FILLER_7_3527 ();
 sg13g2_decap_8 FILLER_7_3533 ();
 sg13g2_fill_1 FILLER_7_3552 ();
 sg13g2_decap_4 FILLER_7_3575 ();
 sg13g2_fill_1 FILLER_7_3579 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_4 FILLER_8_7 ();
 sg13g2_decap_4 FILLER_8_15 ();
 sg13g2_decap_4 FILLER_8_38 ();
 sg13g2_fill_1 FILLER_8_42 ();
 sg13g2_fill_1 FILLER_8_53 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_fill_1 FILLER_8_70 ();
 sg13g2_fill_2 FILLER_8_80 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_fill_2 FILLER_8_98 ();
 sg13g2_fill_1 FILLER_8_100 ();
 sg13g2_fill_2 FILLER_8_111 ();
 sg13g2_fill_2 FILLER_8_127 ();
 sg13g2_fill_1 FILLER_8_129 ();
 sg13g2_decap_8 FILLER_8_142 ();
 sg13g2_decap_4 FILLER_8_149 ();
 sg13g2_fill_1 FILLER_8_157 ();
 sg13g2_fill_1 FILLER_8_204 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_fill_1 FILLER_8_238 ();
 sg13g2_fill_2 FILLER_8_244 ();
 sg13g2_fill_1 FILLER_8_246 ();
 sg13g2_fill_1 FILLER_8_251 ();
 sg13g2_decap_8 FILLER_8_256 ();
 sg13g2_fill_2 FILLER_8_263 ();
 sg13g2_fill_1 FILLER_8_265 ();
 sg13g2_decap_4 FILLER_8_292 ();
 sg13g2_fill_1 FILLER_8_296 ();
 sg13g2_decap_4 FILLER_8_316 ();
 sg13g2_fill_1 FILLER_8_320 ();
 sg13g2_fill_2 FILLER_8_387 ();
 sg13g2_fill_1 FILLER_8_389 ();
 sg13g2_decap_8 FILLER_8_425 ();
 sg13g2_fill_2 FILLER_8_432 ();
 sg13g2_decap_8 FILLER_8_442 ();
 sg13g2_decap_4 FILLER_8_449 ();
 sg13g2_decap_8 FILLER_8_457 ();
 sg13g2_decap_8 FILLER_8_464 ();
 sg13g2_decap_8 FILLER_8_471 ();
 sg13g2_decap_8 FILLER_8_486 ();
 sg13g2_fill_2 FILLER_8_493 ();
 sg13g2_fill_2 FILLER_8_515 ();
 sg13g2_fill_2 FILLER_8_527 ();
 sg13g2_fill_2 FILLER_8_543 ();
 sg13g2_fill_1 FILLER_8_545 ();
 sg13g2_decap_4 FILLER_8_559 ();
 sg13g2_fill_2 FILLER_8_563 ();
 sg13g2_fill_2 FILLER_8_601 ();
 sg13g2_fill_1 FILLER_8_603 ();
 sg13g2_decap_8 FILLER_8_626 ();
 sg13g2_fill_2 FILLER_8_633 ();
 sg13g2_fill_1 FILLER_8_635 ();
 sg13g2_decap_8 FILLER_8_662 ();
 sg13g2_decap_4 FILLER_8_669 ();
 sg13g2_fill_2 FILLER_8_678 ();
 sg13g2_fill_1 FILLER_8_684 ();
 sg13g2_fill_2 FILLER_8_689 ();
 sg13g2_decap_4 FILLER_8_700 ();
 sg13g2_fill_2 FILLER_8_704 ();
 sg13g2_fill_2 FILLER_8_711 ();
 sg13g2_fill_1 FILLER_8_774 ();
 sg13g2_decap_4 FILLER_8_796 ();
 sg13g2_fill_2 FILLER_8_818 ();
 sg13g2_fill_1 FILLER_8_820 ();
 sg13g2_fill_2 FILLER_8_829 ();
 sg13g2_fill_1 FILLER_8_831 ();
 sg13g2_fill_2 FILLER_8_840 ();
 sg13g2_fill_1 FILLER_8_842 ();
 sg13g2_fill_2 FILLER_8_861 ();
 sg13g2_fill_2 FILLER_8_897 ();
 sg13g2_fill_1 FILLER_8_899 ();
 sg13g2_fill_1 FILLER_8_909 ();
 sg13g2_fill_2 FILLER_8_918 ();
 sg13g2_decap_8 FILLER_8_934 ();
 sg13g2_fill_2 FILLER_8_941 ();
 sg13g2_decap_4 FILLER_8_952 ();
 sg13g2_fill_1 FILLER_8_965 ();
 sg13g2_fill_1 FILLER_8_999 ();
 sg13g2_fill_1 FILLER_8_1016 ();
 sg13g2_decap_8 FILLER_8_1043 ();
 sg13g2_fill_2 FILLER_8_1050 ();
 sg13g2_fill_1 FILLER_8_1052 ();
 sg13g2_fill_2 FILLER_8_1100 ();
 sg13g2_decap_8 FILLER_8_1105 ();
 sg13g2_decap_8 FILLER_8_1112 ();
 sg13g2_fill_2 FILLER_8_1123 ();
 sg13g2_decap_8 FILLER_8_1129 ();
 sg13g2_fill_1 FILLER_8_1146 ();
 sg13g2_decap_4 FILLER_8_1154 ();
 sg13g2_fill_2 FILLER_8_1158 ();
 sg13g2_decap_8 FILLER_8_1164 ();
 sg13g2_fill_2 FILLER_8_1202 ();
 sg13g2_fill_2 FILLER_8_1212 ();
 sg13g2_fill_1 FILLER_8_1214 ();
 sg13g2_decap_4 FILLER_8_1220 ();
 sg13g2_fill_1 FILLER_8_1240 ();
 sg13g2_decap_8 FILLER_8_1267 ();
 sg13g2_fill_2 FILLER_8_1285 ();
 sg13g2_fill_1 FILLER_8_1314 ();
 sg13g2_fill_2 FILLER_8_1336 ();
 sg13g2_fill_1 FILLER_8_1338 ();
 sg13g2_decap_4 FILLER_8_1356 ();
 sg13g2_decap_8 FILLER_8_1398 ();
 sg13g2_decap_8 FILLER_8_1405 ();
 sg13g2_decap_4 FILLER_8_1412 ();
 sg13g2_fill_1 FILLER_8_1416 ();
 sg13g2_fill_1 FILLER_8_1448 ();
 sg13g2_decap_4 FILLER_8_1479 ();
 sg13g2_fill_2 FILLER_8_1488 ();
 sg13g2_fill_1 FILLER_8_1490 ();
 sg13g2_decap_4 FILLER_8_1495 ();
 sg13g2_fill_1 FILLER_8_1499 ();
 sg13g2_fill_2 FILLER_8_1543 ();
 sg13g2_fill_2 FILLER_8_1550 ();
 sg13g2_fill_2 FILLER_8_1560 ();
 sg13g2_decap_4 FILLER_8_1575 ();
 sg13g2_decap_8 FILLER_8_1583 ();
 sg13g2_fill_1 FILLER_8_1590 ();
 sg13g2_decap_8 FILLER_8_1599 ();
 sg13g2_decap_8 FILLER_8_1606 ();
 sg13g2_decap_8 FILLER_8_1630 ();
 sg13g2_fill_2 FILLER_8_1637 ();
 sg13g2_fill_1 FILLER_8_1639 ();
 sg13g2_fill_1 FILLER_8_1713 ();
 sg13g2_decap_8 FILLER_8_1718 ();
 sg13g2_decap_4 FILLER_8_1725 ();
 sg13g2_decap_4 FILLER_8_1776 ();
 sg13g2_fill_2 FILLER_8_1780 ();
 sg13g2_fill_2 FILLER_8_1815 ();
 sg13g2_fill_2 FILLER_8_1822 ();
 sg13g2_fill_1 FILLER_8_1824 ();
 sg13g2_decap_8 FILLER_8_1846 ();
 sg13g2_fill_2 FILLER_8_1853 ();
 sg13g2_fill_2 FILLER_8_1860 ();
 sg13g2_fill_2 FILLER_8_1875 ();
 sg13g2_decap_8 FILLER_8_1890 ();
 sg13g2_fill_2 FILLER_8_1915 ();
 sg13g2_fill_1 FILLER_8_1917 ();
 sg13g2_fill_2 FILLER_8_1944 ();
 sg13g2_decap_4 FILLER_8_1964 ();
 sg13g2_fill_1 FILLER_8_1968 ();
 sg13g2_fill_1 FILLER_8_1974 ();
 sg13g2_fill_2 FILLER_8_1980 ();
 sg13g2_fill_1 FILLER_8_1987 ();
 sg13g2_decap_4 FILLER_8_1996 ();
 sg13g2_fill_2 FILLER_8_2029 ();
 sg13g2_decap_8 FILLER_8_2066 ();
 sg13g2_decap_8 FILLER_8_2073 ();
 sg13g2_decap_4 FILLER_8_2080 ();
 sg13g2_fill_1 FILLER_8_2084 ();
 sg13g2_decap_8 FILLER_8_2089 ();
 sg13g2_fill_2 FILLER_8_2096 ();
 sg13g2_fill_1 FILLER_8_2115 ();
 sg13g2_decap_8 FILLER_8_2127 ();
 sg13g2_fill_2 FILLER_8_2134 ();
 sg13g2_decap_8 FILLER_8_2150 ();
 sg13g2_decap_4 FILLER_8_2157 ();
 sg13g2_fill_2 FILLER_8_2161 ();
 sg13g2_fill_2 FILLER_8_2171 ();
 sg13g2_fill_1 FILLER_8_2173 ();
 sg13g2_decap_4 FILLER_8_2179 ();
 sg13g2_decap_8 FILLER_8_2188 ();
 sg13g2_decap_4 FILLER_8_2220 ();
 sg13g2_decap_8 FILLER_8_2253 ();
 sg13g2_decap_4 FILLER_8_2260 ();
 sg13g2_fill_2 FILLER_8_2264 ();
 sg13g2_decap_4 FILLER_8_2279 ();
 sg13g2_fill_2 FILLER_8_2283 ();
 sg13g2_fill_2 FILLER_8_2290 ();
 sg13g2_fill_1 FILLER_8_2292 ();
 sg13g2_fill_1 FILLER_8_2301 ();
 sg13g2_fill_1 FILLER_8_2311 ();
 sg13g2_decap_8 FILLER_8_2321 ();
 sg13g2_decap_8 FILLER_8_2336 ();
 sg13g2_fill_2 FILLER_8_2343 ();
 sg13g2_decap_8 FILLER_8_2356 ();
 sg13g2_decap_4 FILLER_8_2363 ();
 sg13g2_fill_2 FILLER_8_2380 ();
 sg13g2_fill_2 FILLER_8_2396 ();
 sg13g2_fill_1 FILLER_8_2398 ();
 sg13g2_fill_1 FILLER_8_2425 ();
 sg13g2_decap_8 FILLER_8_2447 ();
 sg13g2_decap_8 FILLER_8_2454 ();
 sg13g2_fill_1 FILLER_8_2485 ();
 sg13g2_fill_2 FILLER_8_2521 ();
 sg13g2_fill_1 FILLER_8_2523 ();
 sg13g2_fill_1 FILLER_8_2545 ();
 sg13g2_fill_2 FILLER_8_2550 ();
 sg13g2_decap_8 FILLER_8_2573 ();
 sg13g2_decap_8 FILLER_8_2580 ();
 sg13g2_fill_2 FILLER_8_2606 ();
 sg13g2_fill_1 FILLER_8_2608 ();
 sg13g2_decap_4 FILLER_8_2618 ();
 sg13g2_fill_2 FILLER_8_2622 ();
 sg13g2_decap_8 FILLER_8_2647 ();
 sg13g2_decap_8 FILLER_8_2654 ();
 sg13g2_decap_4 FILLER_8_2661 ();
 sg13g2_fill_1 FILLER_8_2665 ();
 sg13g2_decap_4 FILLER_8_2670 ();
 sg13g2_fill_1 FILLER_8_2674 ();
 sg13g2_decap_4 FILLER_8_2684 ();
 sg13g2_fill_1 FILLER_8_2688 ();
 sg13g2_fill_1 FILLER_8_2694 ();
 sg13g2_decap_8 FILLER_8_2700 ();
 sg13g2_decap_8 FILLER_8_2707 ();
 sg13g2_fill_1 FILLER_8_2714 ();
 sg13g2_decap_8 FILLER_8_2729 ();
 sg13g2_fill_2 FILLER_8_2736 ();
 sg13g2_fill_1 FILLER_8_2738 ();
 sg13g2_decap_4 FILLER_8_2767 ();
 sg13g2_fill_2 FILLER_8_2784 ();
 sg13g2_fill_1 FILLER_8_2786 ();
 sg13g2_fill_2 FILLER_8_2805 ();
 sg13g2_fill_1 FILLER_8_2807 ();
 sg13g2_decap_8 FILLER_8_2818 ();
 sg13g2_decap_4 FILLER_8_2825 ();
 sg13g2_fill_1 FILLER_8_2829 ();
 sg13g2_decap_4 FILLER_8_2834 ();
 sg13g2_fill_2 FILLER_8_2838 ();
 sg13g2_decap_8 FILLER_8_2875 ();
 sg13g2_decap_4 FILLER_8_2882 ();
 sg13g2_decap_4 FILLER_8_2925 ();
 sg13g2_fill_1 FILLER_8_2929 ();
 sg13g2_fill_1 FILLER_8_2938 ();
 sg13g2_decap_8 FILLER_8_2986 ();
 sg13g2_fill_1 FILLER_8_3001 ();
 sg13g2_decap_4 FILLER_8_3011 ();
 sg13g2_fill_1 FILLER_8_3015 ();
 sg13g2_decap_8 FILLER_8_3040 ();
 sg13g2_fill_2 FILLER_8_3047 ();
 sg13g2_fill_1 FILLER_8_3049 ();
 sg13g2_fill_2 FILLER_8_3076 ();
 sg13g2_fill_2 FILLER_8_3087 ();
 sg13g2_fill_2 FILLER_8_3147 ();
 sg13g2_fill_1 FILLER_8_3149 ();
 sg13g2_decap_8 FILLER_8_3176 ();
 sg13g2_fill_1 FILLER_8_3191 ();
 sg13g2_decap_8 FILLER_8_3222 ();
 sg13g2_fill_2 FILLER_8_3229 ();
 sg13g2_fill_1 FILLER_8_3252 ();
 sg13g2_decap_4 FILLER_8_3257 ();
 sg13g2_fill_1 FILLER_8_3261 ();
 sg13g2_fill_2 FILLER_8_3275 ();
 sg13g2_decap_4 FILLER_8_3282 ();
 sg13g2_fill_2 FILLER_8_3286 ();
 sg13g2_decap_4 FILLER_8_3293 ();
 sg13g2_decap_4 FILLER_8_3312 ();
 sg13g2_fill_1 FILLER_8_3321 ();
 sg13g2_decap_4 FILLER_8_3326 ();
 sg13g2_fill_1 FILLER_8_3330 ();
 sg13g2_fill_2 FILLER_8_3353 ();
 sg13g2_decap_8 FILLER_8_3380 ();
 sg13g2_decap_4 FILLER_8_3402 ();
 sg13g2_fill_1 FILLER_8_3406 ();
 sg13g2_fill_1 FILLER_8_3412 ();
 sg13g2_decap_4 FILLER_8_3431 ();
 sg13g2_decap_8 FILLER_8_3457 ();
 sg13g2_fill_1 FILLER_8_3464 ();
 sg13g2_decap_8 FILLER_8_3500 ();
 sg13g2_fill_2 FILLER_8_3538 ();
 sg13g2_fill_1 FILLER_8_3540 ();
 sg13g2_fill_2 FILLER_8_3577 ();
 sg13g2_fill_1 FILLER_8_3579 ();
 sg13g2_fill_2 FILLER_9_26 ();
 sg13g2_fill_1 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_52 ();
 sg13g2_decap_4 FILLER_9_59 ();
 sg13g2_fill_1 FILLER_9_67 ();
 sg13g2_fill_1 FILLER_9_78 ();
 sg13g2_decap_4 FILLER_9_100 ();
 sg13g2_fill_2 FILLER_9_130 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_4 FILLER_9_175 ();
 sg13g2_fill_1 FILLER_9_179 ();
 sg13g2_fill_2 FILLER_9_193 ();
 sg13g2_fill_1 FILLER_9_195 ();
 sg13g2_fill_1 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_fill_1 FILLER_9_294 ();
 sg13g2_decap_4 FILLER_9_305 ();
 sg13g2_fill_2 FILLER_9_309 ();
 sg13g2_decap_8 FILLER_9_338 ();
 sg13g2_decap_8 FILLER_9_345 ();
 sg13g2_fill_1 FILLER_9_382 ();
 sg13g2_fill_1 FILLER_9_392 ();
 sg13g2_fill_2 FILLER_9_402 ();
 sg13g2_fill_1 FILLER_9_409 ();
 sg13g2_fill_2 FILLER_9_414 ();
 sg13g2_fill_1 FILLER_9_416 ();
 sg13g2_fill_1 FILLER_9_451 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_fill_2 FILLER_9_469 ();
 sg13g2_fill_2 FILLER_9_497 ();
 sg13g2_decap_8 FILLER_9_507 ();
 sg13g2_fill_1 FILLER_9_514 ();
 sg13g2_decap_8 FILLER_9_519 ();
 sg13g2_decap_8 FILLER_9_526 ();
 sg13g2_fill_2 FILLER_9_533 ();
 sg13g2_fill_1 FILLER_9_535 ();
 sg13g2_fill_2 FILLER_9_541 ();
 sg13g2_fill_2 FILLER_9_547 ();
 sg13g2_fill_1 FILLER_9_549 ();
 sg13g2_decap_4 FILLER_9_572 ();
 sg13g2_fill_1 FILLER_9_576 ();
 sg13g2_decap_8 FILLER_9_590 ();
 sg13g2_fill_2 FILLER_9_597 ();
 sg13g2_fill_1 FILLER_9_599 ();
 sg13g2_decap_8 FILLER_9_626 ();
 sg13g2_fill_1 FILLER_9_633 ();
 sg13g2_fill_2 FILLER_9_643 ();
 sg13g2_fill_2 FILLER_9_650 ();
 sg13g2_fill_1 FILLER_9_666 ();
 sg13g2_decap_8 FILLER_9_671 ();
 sg13g2_fill_1 FILLER_9_678 ();
 sg13g2_decap_4 FILLER_9_687 ();
 sg13g2_fill_2 FILLER_9_691 ();
 sg13g2_decap_8 FILLER_9_706 ();
 sg13g2_decap_8 FILLER_9_713 ();
 sg13g2_fill_2 FILLER_9_720 ();
 sg13g2_fill_1 FILLER_9_722 ();
 sg13g2_fill_2 FILLER_9_731 ();
 sg13g2_fill_1 FILLER_9_733 ();
 sg13g2_fill_1 FILLER_9_739 ();
 sg13g2_fill_1 FILLER_9_757 ();
 sg13g2_fill_1 FILLER_9_772 ();
 sg13g2_fill_2 FILLER_9_794 ();
 sg13g2_fill_1 FILLER_9_796 ();
 sg13g2_decap_8 FILLER_9_802 ();
 sg13g2_decap_8 FILLER_9_873 ();
 sg13g2_decap_8 FILLER_9_880 ();
 sg13g2_decap_8 FILLER_9_887 ();
 sg13g2_fill_2 FILLER_9_908 ();
 sg13g2_decap_8 FILLER_9_962 ();
 sg13g2_decap_8 FILLER_9_991 ();
 sg13g2_decap_8 FILLER_9_998 ();
 sg13g2_decap_8 FILLER_9_1005 ();
 sg13g2_fill_2 FILLER_9_1012 ();
 sg13g2_fill_2 FILLER_9_1018 ();
 sg13g2_fill_1 FILLER_9_1020 ();
 sg13g2_fill_2 FILLER_9_1026 ();
 sg13g2_fill_1 FILLER_9_1028 ();
 sg13g2_fill_1 FILLER_9_1043 ();
 sg13g2_decap_8 FILLER_9_1052 ();
 sg13g2_fill_2 FILLER_9_1059 ();
 sg13g2_fill_1 FILLER_9_1080 ();
 sg13g2_decap_4 FILLER_9_1090 ();
 sg13g2_fill_1 FILLER_9_1094 ();
 sg13g2_fill_1 FILLER_9_1127 ();
 sg13g2_fill_1 FILLER_9_1141 ();
 sg13g2_fill_2 FILLER_9_1147 ();
 sg13g2_fill_2 FILLER_9_1167 ();
 sg13g2_decap_4 FILLER_9_1188 ();
 sg13g2_fill_2 FILLER_9_1192 ();
 sg13g2_decap_8 FILLER_9_1225 ();
 sg13g2_decap_8 FILLER_9_1232 ();
 sg13g2_fill_1 FILLER_9_1239 ();
 sg13g2_fill_2 FILLER_9_1249 ();
 sg13g2_fill_1 FILLER_9_1251 ();
 sg13g2_fill_1 FILLER_9_1256 ();
 sg13g2_decap_8 FILLER_9_1266 ();
 sg13g2_decap_4 FILLER_9_1278 ();
 sg13g2_fill_2 FILLER_9_1287 ();
 sg13g2_fill_1 FILLER_9_1289 ();
 sg13g2_decap_8 FILLER_9_1302 ();
 sg13g2_fill_2 FILLER_9_1309 ();
 sg13g2_fill_1 FILLER_9_1311 ();
 sg13g2_fill_2 FILLER_9_1326 ();
 sg13g2_fill_1 FILLER_9_1341 ();
 sg13g2_decap_8 FILLER_9_1349 ();
 sg13g2_decap_4 FILLER_9_1356 ();
 sg13g2_fill_2 FILLER_9_1360 ();
 sg13g2_decap_8 FILLER_9_1367 ();
 sg13g2_decap_4 FILLER_9_1374 ();
 sg13g2_fill_1 FILLER_9_1378 ();
 sg13g2_fill_1 FILLER_9_1383 ();
 sg13g2_fill_2 FILLER_9_1424 ();
 sg13g2_fill_1 FILLER_9_1426 ();
 sg13g2_decap_8 FILLER_9_1437 ();
 sg13g2_decap_8 FILLER_9_1444 ();
 sg13g2_fill_2 FILLER_9_1451 ();
 sg13g2_fill_1 FILLER_9_1453 ();
 sg13g2_fill_2 FILLER_9_1462 ();
 sg13g2_fill_2 FILLER_9_1524 ();
 sg13g2_fill_2 FILLER_9_1550 ();
 sg13g2_fill_2 FILLER_9_1560 ();
 sg13g2_fill_1 FILLER_9_1578 ();
 sg13g2_decap_8 FILLER_9_1622 ();
 sg13g2_decap_4 FILLER_9_1629 ();
 sg13g2_decap_8 FILLER_9_1641 ();
 sg13g2_fill_2 FILLER_9_1648 ();
 sg13g2_fill_1 FILLER_9_1650 ();
 sg13g2_decap_4 FILLER_9_1655 ();
 sg13g2_fill_1 FILLER_9_1659 ();
 sg13g2_fill_1 FILLER_9_1669 ();
 sg13g2_decap_4 FILLER_9_1681 ();
 sg13g2_decap_4 FILLER_9_1694 ();
 sg13g2_decap_8 FILLER_9_1711 ();
 sg13g2_decap_8 FILLER_9_1774 ();
 sg13g2_decap_4 FILLER_9_1781 ();
 sg13g2_fill_2 FILLER_9_1785 ();
 sg13g2_fill_2 FILLER_9_1798 ();
 sg13g2_fill_1 FILLER_9_1800 ();
 sg13g2_decap_4 FILLER_9_1811 ();
 sg13g2_fill_2 FILLER_9_1815 ();
 sg13g2_fill_2 FILLER_9_1848 ();
 sg13g2_decap_4 FILLER_9_1876 ();
 sg13g2_fill_2 FILLER_9_1880 ();
 sg13g2_decap_4 FILLER_9_1892 ();
 sg13g2_decap_8 FILLER_9_1901 ();
 sg13g2_fill_1 FILLER_9_1908 ();
 sg13g2_decap_8 FILLER_9_1914 ();
 sg13g2_decap_8 FILLER_9_1925 ();
 sg13g2_decap_4 FILLER_9_1932 ();
 sg13g2_fill_2 FILLER_9_1936 ();
 sg13g2_fill_1 FILLER_9_1946 ();
 sg13g2_decap_8 FILLER_9_1957 ();
 sg13g2_decap_4 FILLER_9_1964 ();
 sg13g2_fill_1 FILLER_9_1968 ();
 sg13g2_fill_2 FILLER_9_1973 ();
 sg13g2_decap_8 FILLER_9_1989 ();
 sg13g2_decap_4 FILLER_9_1996 ();
 sg13g2_decap_4 FILLER_9_2015 ();
 sg13g2_fill_2 FILLER_9_2019 ();
 sg13g2_decap_4 FILLER_9_2028 ();
 sg13g2_fill_2 FILLER_9_2032 ();
 sg13g2_fill_2 FILLER_9_2047 ();
 sg13g2_fill_1 FILLER_9_2049 ();
 sg13g2_decap_4 FILLER_9_2063 ();
 sg13g2_fill_1 FILLER_9_2067 ();
 sg13g2_decap_4 FILLER_9_2077 ();
 sg13g2_fill_2 FILLER_9_2081 ();
 sg13g2_decap_4 FILLER_9_2092 ();
 sg13g2_decap_4 FILLER_9_2101 ();
 sg13g2_fill_2 FILLER_9_2114 ();
 sg13g2_decap_4 FILLER_9_2129 ();
 sg13g2_fill_2 FILLER_9_2159 ();
 sg13g2_decap_4 FILLER_9_2173 ();
 sg13g2_fill_2 FILLER_9_2182 ();
 sg13g2_fill_2 FILLER_9_2192 ();
 sg13g2_decap_8 FILLER_9_2198 ();
 sg13g2_fill_2 FILLER_9_2205 ();
 sg13g2_fill_2 FILLER_9_2226 ();
 sg13g2_fill_1 FILLER_9_2228 ();
 sg13g2_decap_8 FILLER_9_2264 ();
 sg13g2_fill_2 FILLER_9_2271 ();
 sg13g2_decap_8 FILLER_9_2282 ();
 sg13g2_fill_1 FILLER_9_2295 ();
 sg13g2_fill_2 FILLER_9_2301 ();
 sg13g2_decap_8 FILLER_9_2313 ();
 sg13g2_fill_2 FILLER_9_2320 ();
 sg13g2_fill_1 FILLER_9_2322 ();
 sg13g2_fill_1 FILLER_9_2332 ();
 sg13g2_fill_1 FILLER_9_2337 ();
 sg13g2_decap_8 FILLER_9_2365 ();
 sg13g2_fill_2 FILLER_9_2372 ();
 sg13g2_fill_1 FILLER_9_2374 ();
 sg13g2_decap_8 FILLER_9_2401 ();
 sg13g2_fill_2 FILLER_9_2408 ();
 sg13g2_fill_1 FILLER_9_2423 ();
 sg13g2_fill_2 FILLER_9_2452 ();
 sg13g2_fill_1 FILLER_9_2454 ();
 sg13g2_decap_8 FILLER_9_2485 ();
 sg13g2_decap_8 FILLER_9_2492 ();
 sg13g2_fill_2 FILLER_9_2499 ();
 sg13g2_fill_1 FILLER_9_2501 ();
 sg13g2_decap_8 FILLER_9_2506 ();
 sg13g2_decap_4 FILLER_9_2513 ();
 sg13g2_decap_4 FILLER_9_2525 ();
 sg13g2_fill_1 FILLER_9_2529 ();
 sg13g2_fill_2 FILLER_9_2545 ();
 sg13g2_fill_2 FILLER_9_2558 ();
 sg13g2_fill_1 FILLER_9_2560 ();
 sg13g2_decap_4 FILLER_9_2569 ();
 sg13g2_decap_4 FILLER_9_2581 ();
 sg13g2_fill_1 FILLER_9_2585 ();
 sg13g2_fill_2 FILLER_9_2594 ();
 sg13g2_fill_1 FILLER_9_2596 ();
 sg13g2_decap_8 FILLER_9_2604 ();
 sg13g2_decap_4 FILLER_9_2611 ();
 sg13g2_fill_1 FILLER_9_2615 ();
 sg13g2_decap_8 FILLER_9_2641 ();
 sg13g2_fill_1 FILLER_9_2648 ();
 sg13g2_decap_8 FILLER_9_2684 ();
 sg13g2_decap_8 FILLER_9_2691 ();
 sg13g2_fill_2 FILLER_9_2698 ();
 sg13g2_fill_2 FILLER_9_2705 ();
 sg13g2_decap_8 FILLER_9_2711 ();
 sg13g2_fill_2 FILLER_9_2718 ();
 sg13g2_decap_8 FILLER_9_2741 ();
 sg13g2_decap_8 FILLER_9_2748 ();
 sg13g2_fill_1 FILLER_9_2755 ();
 sg13g2_decap_8 FILLER_9_2782 ();
 sg13g2_fill_1 FILLER_9_2789 ();
 sg13g2_fill_2 FILLER_9_2795 ();
 sg13g2_decap_4 FILLER_9_2802 ();
 sg13g2_fill_2 FILLER_9_2810 ();
 sg13g2_fill_1 FILLER_9_2812 ();
 sg13g2_decap_4 FILLER_9_2818 ();
 sg13g2_fill_1 FILLER_9_2822 ();
 sg13g2_decap_4 FILLER_9_2827 ();
 sg13g2_fill_2 FILLER_9_2848 ();
 sg13g2_fill_2 FILLER_9_2867 ();
 sg13g2_decap_4 FILLER_9_2882 ();
 sg13g2_decap_4 FILLER_9_2899 ();
 sg13g2_fill_1 FILLER_9_2907 ();
 sg13g2_decap_4 FILLER_9_2913 ();
 sg13g2_fill_1 FILLER_9_2917 ();
 sg13g2_decap_8 FILLER_9_2929 ();
 sg13g2_fill_2 FILLER_9_2941 ();
 sg13g2_fill_1 FILLER_9_2943 ();
 sg13g2_fill_1 FILLER_9_2975 ();
 sg13g2_fill_1 FILLER_9_2990 ();
 sg13g2_fill_2 FILLER_9_3020 ();
 sg13g2_fill_2 FILLER_9_3040 ();
 sg13g2_fill_1 FILLER_9_3042 ();
 sg13g2_fill_2 FILLER_9_3052 ();
 sg13g2_fill_1 FILLER_9_3064 ();
 sg13g2_decap_8 FILLER_9_3078 ();
 sg13g2_decap_4 FILLER_9_3085 ();
 sg13g2_decap_4 FILLER_9_3105 ();
 sg13g2_fill_1 FILLER_9_3109 ();
 sg13g2_decap_4 FILLER_9_3120 ();
 sg13g2_fill_1 FILLER_9_3154 ();
 sg13g2_decap_4 FILLER_9_3182 ();
 sg13g2_fill_1 FILLER_9_3186 ();
 sg13g2_fill_1 FILLER_9_3192 ();
 sg13g2_decap_4 FILLER_9_3197 ();
 sg13g2_fill_2 FILLER_9_3201 ();
 sg13g2_decap_8 FILLER_9_3216 ();
 sg13g2_decap_4 FILLER_9_3223 ();
 sg13g2_decap_4 FILLER_9_3258 ();
 sg13g2_fill_1 FILLER_9_3267 ();
 sg13g2_fill_2 FILLER_9_3272 ();
 sg13g2_fill_1 FILLER_9_3274 ();
 sg13g2_fill_2 FILLER_9_3286 ();
 sg13g2_fill_1 FILLER_9_3288 ();
 sg13g2_fill_2 FILLER_9_3294 ();
 sg13g2_fill_2 FILLER_9_3310 ();
 sg13g2_decap_8 FILLER_9_3404 ();
 sg13g2_decap_4 FILLER_9_3411 ();
 sg13g2_fill_1 FILLER_9_3415 ();
 sg13g2_fill_2 FILLER_9_3424 ();
 sg13g2_decap_8 FILLER_9_3452 ();
 sg13g2_fill_2 FILLER_9_3473 ();
 sg13g2_fill_2 FILLER_9_3481 ();
 sg13g2_fill_2 FILLER_9_3504 ();
 sg13g2_fill_1 FILLER_9_3506 ();
 sg13g2_decap_4 FILLER_9_3515 ();
 sg13g2_decap_8 FILLER_9_3523 ();
 sg13g2_fill_1 FILLER_9_3530 ();
 sg13g2_fill_2 FILLER_9_3536 ();
 sg13g2_fill_2 FILLER_9_3577 ();
 sg13g2_fill_1 FILLER_9_3579 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_4 FILLER_10_7 ();
 sg13g2_fill_2 FILLER_10_11 ();
 sg13g2_decap_4 FILLER_10_22 ();
 sg13g2_decap_8 FILLER_10_87 ();
 sg13g2_fill_2 FILLER_10_94 ();
 sg13g2_fill_1 FILLER_10_114 ();
 sg13g2_fill_2 FILLER_10_129 ();
 sg13g2_fill_1 FILLER_10_151 ();
 sg13g2_fill_2 FILLER_10_161 ();
 sg13g2_fill_1 FILLER_10_163 ();
 sg13g2_decap_8 FILLER_10_200 ();
 sg13g2_fill_1 FILLER_10_233 ();
 sg13g2_fill_2 FILLER_10_238 ();
 sg13g2_fill_1 FILLER_10_276 ();
 sg13g2_fill_1 FILLER_10_281 ();
 sg13g2_decap_4 FILLER_10_299 ();
 sg13g2_fill_1 FILLER_10_303 ();
 sg13g2_fill_2 FILLER_10_324 ();
 sg13g2_decap_4 FILLER_10_339 ();
 sg13g2_fill_1 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_348 ();
 sg13g2_fill_1 FILLER_10_355 ();
 sg13g2_fill_1 FILLER_10_361 ();
 sg13g2_fill_2 FILLER_10_470 ();
 sg13g2_fill_1 FILLER_10_472 ();
 sg13g2_fill_2 FILLER_10_495 ();
 sg13g2_fill_2 FILLER_10_518 ();
 sg13g2_fill_1 FILLER_10_520 ();
 sg13g2_fill_2 FILLER_10_530 ();
 sg13g2_fill_2 FILLER_10_550 ();
 sg13g2_fill_1 FILLER_10_552 ();
 sg13g2_fill_2 FILLER_10_571 ();
 sg13g2_fill_1 FILLER_10_573 ();
 sg13g2_decap_8 FILLER_10_583 ();
 sg13g2_fill_1 FILLER_10_590 ();
 sg13g2_fill_1 FILLER_10_600 ();
 sg13g2_fill_2 FILLER_10_609 ();
 sg13g2_fill_2 FILLER_10_615 ();
 sg13g2_fill_1 FILLER_10_617 ();
 sg13g2_decap_4 FILLER_10_623 ();
 sg13g2_fill_2 FILLER_10_653 ();
 sg13g2_fill_1 FILLER_10_655 ();
 sg13g2_fill_1 FILLER_10_735 ();
 sg13g2_fill_1 FILLER_10_762 ();
 sg13g2_decap_8 FILLER_10_798 ();
 sg13g2_decap_8 FILLER_10_805 ();
 sg13g2_fill_1 FILLER_10_812 ();
 sg13g2_decap_8 FILLER_10_843 ();
 sg13g2_fill_2 FILLER_10_850 ();
 sg13g2_fill_1 FILLER_10_852 ();
 sg13g2_fill_2 FILLER_10_861 ();
 sg13g2_fill_1 FILLER_10_863 ();
 sg13g2_decap_4 FILLER_10_873 ();
 sg13g2_fill_2 FILLER_10_908 ();
 sg13g2_fill_1 FILLER_10_910 ();
 sg13g2_fill_2 FILLER_10_919 ();
 sg13g2_fill_2 FILLER_10_924 ();
 sg13g2_fill_1 FILLER_10_926 ();
 sg13g2_decap_8 FILLER_10_935 ();
 sg13g2_decap_4 FILLER_10_942 ();
 sg13g2_fill_1 FILLER_10_946 ();
 sg13g2_fill_2 FILLER_10_951 ();
 sg13g2_fill_1 FILLER_10_953 ();
 sg13g2_fill_2 FILLER_10_989 ();
 sg13g2_fill_1 FILLER_10_991 ();
 sg13g2_decap_8 FILLER_10_1006 ();
 sg13g2_decap_8 FILLER_10_1013 ();
 sg13g2_decap_8 FILLER_10_1020 ();
 sg13g2_fill_1 FILLER_10_1027 ();
 sg13g2_decap_4 FILLER_10_1076 ();
 sg13g2_fill_2 FILLER_10_1080 ();
 sg13g2_decap_8 FILLER_10_1100 ();
 sg13g2_decap_8 FILLER_10_1107 ();
 sg13g2_fill_2 FILLER_10_1114 ();
 sg13g2_fill_1 FILLER_10_1116 ();
 sg13g2_fill_2 FILLER_10_1169 ();
 sg13g2_fill_2 FILLER_10_1198 ();
 sg13g2_decap_4 FILLER_10_1235 ();
 sg13g2_fill_2 FILLER_10_1239 ();
 sg13g2_fill_2 FILLER_10_1323 ();
 sg13g2_decap_8 FILLER_10_1360 ();
 sg13g2_fill_1 FILLER_10_1367 ();
 sg13g2_fill_1 FILLER_10_1373 ();
 sg13g2_decap_8 FILLER_10_1378 ();
 sg13g2_decap_4 FILLER_10_1385 ();
 sg13g2_decap_4 FILLER_10_1403 ();
 sg13g2_fill_2 FILLER_10_1450 ();
 sg13g2_decap_4 FILLER_10_1478 ();
 sg13g2_fill_2 FILLER_10_1487 ();
 sg13g2_decap_8 FILLER_10_1493 ();
 sg13g2_decap_8 FILLER_10_1500 ();
 sg13g2_decap_4 FILLER_10_1507 ();
 sg13g2_decap_8 FILLER_10_1555 ();
 sg13g2_fill_2 FILLER_10_1562 ();
 sg13g2_fill_1 FILLER_10_1564 ();
 sg13g2_decap_8 FILLER_10_1573 ();
 sg13g2_decap_8 FILLER_10_1580 ();
 sg13g2_fill_1 FILLER_10_1587 ();
 sg13g2_decap_8 FILLER_10_1601 ();
 sg13g2_fill_1 FILLER_10_1608 ();
 sg13g2_fill_1 FILLER_10_1644 ();
 sg13g2_decap_8 FILLER_10_1653 ();
 sg13g2_fill_2 FILLER_10_1660 ();
 sg13g2_fill_1 FILLER_10_1662 ();
 sg13g2_fill_2 FILLER_10_1668 ();
 sg13g2_fill_1 FILLER_10_1670 ();
 sg13g2_decap_4 FILLER_10_1675 ();
 sg13g2_fill_2 FILLER_10_1688 ();
 sg13g2_fill_1 FILLER_10_1690 ();
 sg13g2_decap_8 FILLER_10_1706 ();
 sg13g2_fill_1 FILLER_10_1760 ();
 sg13g2_fill_1 FILLER_10_1774 ();
 sg13g2_fill_1 FILLER_10_1783 ();
 sg13g2_decap_4 FILLER_10_1789 ();
 sg13g2_fill_1 FILLER_10_1793 ();
 sg13g2_decap_4 FILLER_10_1799 ();
 sg13g2_fill_1 FILLER_10_1813 ();
 sg13g2_decap_8 FILLER_10_1832 ();
 sg13g2_decap_4 FILLER_10_1839 ();
 sg13g2_fill_1 FILLER_10_1843 ();
 sg13g2_decap_4 FILLER_10_1849 ();
 sg13g2_fill_2 FILLER_10_1853 ();
 sg13g2_fill_1 FILLER_10_1867 ();
 sg13g2_fill_1 FILLER_10_1877 ();
 sg13g2_decap_8 FILLER_10_1891 ();
 sg13g2_fill_1 FILLER_10_1898 ();
 sg13g2_fill_2 FILLER_10_1907 ();
 sg13g2_fill_1 FILLER_10_1909 ();
 sg13g2_fill_2 FILLER_10_1991 ();
 sg13g2_fill_1 FILLER_10_1993 ();
 sg13g2_decap_8 FILLER_10_2012 ();
 sg13g2_decap_4 FILLER_10_2019 ();
 sg13g2_fill_2 FILLER_10_2023 ();
 sg13g2_decap_8 FILLER_10_2030 ();
 sg13g2_fill_1 FILLER_10_2037 ();
 sg13g2_decap_8 FILLER_10_2043 ();
 sg13g2_fill_2 FILLER_10_2050 ();
 sg13g2_decap_8 FILLER_10_2057 ();
 sg13g2_fill_2 FILLER_10_2064 ();
 sg13g2_fill_2 FILLER_10_2092 ();
 sg13g2_fill_1 FILLER_10_2150 ();
 sg13g2_fill_2 FILLER_10_2170 ();
 sg13g2_fill_1 FILLER_10_2172 ();
 sg13g2_fill_1 FILLER_10_2243 ();
 sg13g2_decap_8 FILLER_10_2253 ();
 sg13g2_decap_8 FILLER_10_2260 ();
 sg13g2_fill_2 FILLER_10_2267 ();
 sg13g2_fill_2 FILLER_10_2300 ();
 sg13g2_fill_1 FILLER_10_2302 ();
 sg13g2_fill_2 FILLER_10_2383 ();
 sg13g2_decap_8 FILLER_10_2393 ();
 sg13g2_decap_8 FILLER_10_2400 ();
 sg13g2_fill_1 FILLER_10_2407 ();
 sg13g2_decap_4 FILLER_10_2412 ();
 sg13g2_fill_2 FILLER_10_2416 ();
 sg13g2_decap_8 FILLER_10_2444 ();
 sg13g2_decap_4 FILLER_10_2451 ();
 sg13g2_fill_2 FILLER_10_2455 ();
 sg13g2_decap_8 FILLER_10_2483 ();
 sg13g2_decap_4 FILLER_10_2516 ();
 sg13g2_fill_2 FILLER_10_2550 ();
 sg13g2_fill_1 FILLER_10_2552 ();
 sg13g2_fill_1 FILLER_10_2563 ();
 sg13g2_decap_8 FILLER_10_2573 ();
 sg13g2_decap_4 FILLER_10_2580 ();
 sg13g2_fill_2 FILLER_10_2584 ();
 sg13g2_fill_1 FILLER_10_2594 ();
 sg13g2_decap_8 FILLER_10_2605 ();
 sg13g2_decap_8 FILLER_10_2612 ();
 sg13g2_fill_2 FILLER_10_2619 ();
 sg13g2_fill_1 FILLER_10_2621 ();
 sg13g2_fill_2 FILLER_10_2661 ();
 sg13g2_fill_1 FILLER_10_2663 ();
 sg13g2_fill_2 FILLER_10_2747 ();
 sg13g2_fill_1 FILLER_10_2749 ();
 sg13g2_fill_2 FILLER_10_2764 ();
 sg13g2_fill_1 FILLER_10_2766 ();
 sg13g2_decap_4 FILLER_10_2792 ();
 sg13g2_fill_1 FILLER_10_2796 ();
 sg13g2_fill_1 FILLER_10_2812 ();
 sg13g2_fill_2 FILLER_10_2823 ();
 sg13g2_fill_2 FILLER_10_2850 ();
 sg13g2_fill_2 FILLER_10_2883 ();
 sg13g2_fill_1 FILLER_10_2885 ();
 sg13g2_decap_4 FILLER_10_2904 ();
 sg13g2_fill_1 FILLER_10_2908 ();
 sg13g2_fill_1 FILLER_10_2930 ();
 sg13g2_decap_4 FILLER_10_2940 ();
 sg13g2_fill_2 FILLER_10_2953 ();
 sg13g2_fill_1 FILLER_10_2955 ();
 sg13g2_fill_1 FILLER_10_2969 ();
 sg13g2_fill_2 FILLER_10_2978 ();
 sg13g2_decap_8 FILLER_10_3006 ();
 sg13g2_decap_4 FILLER_10_3013 ();
 sg13g2_fill_2 FILLER_10_3017 ();
 sg13g2_fill_1 FILLER_10_3023 ();
 sg13g2_fill_2 FILLER_10_3029 ();
 sg13g2_fill_1 FILLER_10_3031 ();
 sg13g2_decap_8 FILLER_10_3042 ();
 sg13g2_fill_1 FILLER_10_3049 ();
 sg13g2_fill_2 FILLER_10_3064 ();
 sg13g2_decap_4 FILLER_10_3080 ();
 sg13g2_fill_1 FILLER_10_3084 ();
 sg13g2_fill_1 FILLER_10_3098 ();
 sg13g2_fill_1 FILLER_10_3129 ();
 sg13g2_decap_8 FILLER_10_3141 ();
 sg13g2_fill_1 FILLER_10_3148 ();
 sg13g2_fill_2 FILLER_10_3159 ();
 sg13g2_decap_4 FILLER_10_3178 ();
 sg13g2_fill_1 FILLER_10_3182 ();
 sg13g2_decap_8 FILLER_10_3209 ();
 sg13g2_fill_1 FILLER_10_3216 ();
 sg13g2_fill_1 FILLER_10_3221 ();
 sg13g2_fill_2 FILLER_10_3240 ();
 sg13g2_fill_1 FILLER_10_3242 ();
 sg13g2_fill_1 FILLER_10_3252 ();
 sg13g2_fill_2 FILLER_10_3280 ();
 sg13g2_decap_8 FILLER_10_3308 ();
 sg13g2_decap_8 FILLER_10_3315 ();
 sg13g2_decap_4 FILLER_10_3322 ();
 sg13g2_decap_4 FILLER_10_3335 ();
 sg13g2_fill_1 FILLER_10_3339 ();
 sg13g2_decap_4 FILLER_10_3349 ();
 sg13g2_fill_2 FILLER_10_3353 ();
 sg13g2_fill_2 FILLER_10_3377 ();
 sg13g2_fill_1 FILLER_10_3379 ();
 sg13g2_decap_4 FILLER_10_3389 ();
 sg13g2_fill_1 FILLER_10_3393 ();
 sg13g2_fill_2 FILLER_10_3413 ();
 sg13g2_decap_8 FILLER_10_3451 ();
 sg13g2_decap_8 FILLER_10_3458 ();
 sg13g2_decap_4 FILLER_10_3465 ();
 sg13g2_fill_2 FILLER_10_3474 ();
 sg13g2_fill_1 FILLER_10_3476 ();
 sg13g2_fill_2 FILLER_10_3508 ();
 sg13g2_fill_1 FILLER_10_3510 ();
 sg13g2_fill_2 FILLER_10_3515 ();
 sg13g2_fill_2 FILLER_10_3521 ();
 sg13g2_fill_2 FILLER_10_3542 ();
 sg13g2_fill_1 FILLER_10_3544 ();
 sg13g2_fill_1 FILLER_11_0 ();
 sg13g2_decap_4 FILLER_11_37 ();
 sg13g2_fill_2 FILLER_11_41 ();
 sg13g2_decap_8 FILLER_11_53 ();
 sg13g2_fill_2 FILLER_11_60 ();
 sg13g2_fill_1 FILLER_11_62 ();
 sg13g2_fill_1 FILLER_11_72 ();
 sg13g2_decap_4 FILLER_11_99 ();
 sg13g2_fill_2 FILLER_11_103 ();
 sg13g2_decap_8 FILLER_11_131 ();
 sg13g2_decap_4 FILLER_11_164 ();
 sg13g2_fill_2 FILLER_11_168 ();
 sg13g2_decap_4 FILLER_11_200 ();
 sg13g2_fill_1 FILLER_11_204 ();
 sg13g2_decap_4 FILLER_11_209 ();
 sg13g2_fill_1 FILLER_11_217 ();
 sg13g2_fill_2 FILLER_11_231 ();
 sg13g2_fill_1 FILLER_11_282 ();
 sg13g2_fill_2 FILLER_11_295 ();
 sg13g2_decap_8 FILLER_11_359 ();
 sg13g2_decap_8 FILLER_11_366 ();
 sg13g2_decap_4 FILLER_11_391 ();
 sg13g2_fill_1 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_413 ();
 sg13g2_fill_2 FILLER_11_429 ();
 sg13g2_fill_1 FILLER_11_431 ();
 sg13g2_fill_2 FILLER_11_441 ();
 sg13g2_fill_1 FILLER_11_443 ();
 sg13g2_fill_2 FILLER_11_453 ();
 sg13g2_fill_1 FILLER_11_469 ();
 sg13g2_fill_1 FILLER_11_507 ();
 sg13g2_decap_8 FILLER_11_518 ();
 sg13g2_decap_4 FILLER_11_525 ();
 sg13g2_fill_2 FILLER_11_529 ();
 sg13g2_fill_1 FILLER_11_535 ();
 sg13g2_fill_2 FILLER_11_636 ();
 sg13g2_decap_8 FILLER_11_671 ();
 sg13g2_decap_4 FILLER_11_678 ();
 sg13g2_fill_2 FILLER_11_682 ();
 sg13g2_decap_4 FILLER_11_689 ();
 sg13g2_fill_1 FILLER_11_698 ();
 sg13g2_decap_8 FILLER_11_703 ();
 sg13g2_fill_1 FILLER_11_710 ();
 sg13g2_decap_8 FILLER_11_741 ();
 sg13g2_decap_8 FILLER_11_748 ();
 sg13g2_fill_2 FILLER_11_760 ();
 sg13g2_decap_4 FILLER_11_766 ();
 sg13g2_fill_1 FILLER_11_770 ();
 sg13g2_fill_2 FILLER_11_781 ();
 sg13g2_fill_1 FILLER_11_783 ();
 sg13g2_fill_1 FILLER_11_802 ();
 sg13g2_fill_2 FILLER_11_811 ();
 sg13g2_fill_1 FILLER_11_813 ();
 sg13g2_fill_1 FILLER_11_832 ();
 sg13g2_fill_2 FILLER_11_842 ();
 sg13g2_fill_1 FILLER_11_847 ();
 sg13g2_fill_2 FILLER_11_866 ();
 sg13g2_decap_8 FILLER_11_883 ();
 sg13g2_decap_4 FILLER_11_920 ();
 sg13g2_fill_2 FILLER_11_924 ();
 sg13g2_decap_8 FILLER_11_955 ();
 sg13g2_fill_2 FILLER_11_962 ();
 sg13g2_fill_1 FILLER_11_964 ();
 sg13g2_fill_2 FILLER_11_969 ();
 sg13g2_fill_1 FILLER_11_971 ();
 sg13g2_fill_2 FILLER_11_981 ();
 sg13g2_fill_1 FILLER_11_988 ();
 sg13g2_fill_1 FILLER_11_1036 ();
 sg13g2_decap_8 FILLER_11_1042 ();
 sg13g2_fill_1 FILLER_11_1049 ();
 sg13g2_decap_8 FILLER_11_1110 ();
 sg13g2_decap_8 FILLER_11_1117 ();
 sg13g2_decap_8 FILLER_11_1124 ();
 sg13g2_decap_8 FILLER_11_1131 ();
 sg13g2_decap_8 FILLER_11_1138 ();
 sg13g2_decap_8 FILLER_11_1145 ();
 sg13g2_fill_2 FILLER_11_1160 ();
 sg13g2_fill_2 FILLER_11_1166 ();
 sg13g2_fill_1 FILLER_11_1216 ();
 sg13g2_decap_8 FILLER_11_1252 ();
 sg13g2_decap_8 FILLER_11_1259 ();
 sg13g2_fill_2 FILLER_11_1266 ();
 sg13g2_fill_2 FILLER_11_1272 ();
 sg13g2_fill_1 FILLER_11_1274 ();
 sg13g2_fill_1 FILLER_11_1298 ();
 sg13g2_fill_2 FILLER_11_1311 ();
 sg13g2_fill_1 FILLER_11_1313 ();
 sg13g2_fill_1 FILLER_11_1320 ();
 sg13g2_fill_2 FILLER_11_1361 ();
 sg13g2_fill_2 FILLER_11_1408 ();
 sg13g2_fill_1 FILLER_11_1410 ();
 sg13g2_fill_1 FILLER_11_1421 ();
 sg13g2_decap_8 FILLER_11_1432 ();
 sg13g2_decap_4 FILLER_11_1439 ();
 sg13g2_fill_1 FILLER_11_1443 ();
 sg13g2_fill_2 FILLER_11_1458 ();
 sg13g2_decap_8 FILLER_11_1493 ();
 sg13g2_fill_2 FILLER_11_1500 ();
 sg13g2_fill_1 FILLER_11_1502 ();
 sg13g2_fill_2 FILLER_11_1507 ();
 sg13g2_fill_1 FILLER_11_1509 ();
 sg13g2_decap_4 FILLER_11_1515 ();
 sg13g2_fill_1 FILLER_11_1524 ();
 sg13g2_decap_8 FILLER_11_1529 ();
 sg13g2_fill_1 FILLER_11_1536 ();
 sg13g2_decap_8 FILLER_11_1546 ();
 sg13g2_fill_2 FILLER_11_1553 ();
 sg13g2_fill_1 FILLER_11_1555 ();
 sg13g2_fill_1 FILLER_11_1569 ();
 sg13g2_fill_2 FILLER_11_1578 ();
 sg13g2_decap_4 FILLER_11_1614 ();
 sg13g2_fill_1 FILLER_11_1618 ();
 sg13g2_fill_2 FILLER_11_1640 ();
 sg13g2_decap_4 FILLER_11_1650 ();
 sg13g2_decap_8 FILLER_11_1712 ();
 sg13g2_decap_4 FILLER_11_1737 ();
 sg13g2_decap_4 FILLER_11_1750 ();
 sg13g2_fill_2 FILLER_11_1754 ();
 sg13g2_fill_1 FILLER_11_1782 ();
 sg13g2_decap_4 FILLER_11_1787 ();
 sg13g2_fill_1 FILLER_11_1791 ();
 sg13g2_fill_2 FILLER_11_1842 ();
 sg13g2_fill_1 FILLER_11_1844 ();
 sg13g2_decap_4 FILLER_11_1871 ();
 sg13g2_fill_2 FILLER_11_1875 ();
 sg13g2_fill_1 FILLER_11_1897 ();
 sg13g2_decap_4 FILLER_11_1908 ();
 sg13g2_fill_1 FILLER_11_1916 ();
 sg13g2_fill_2 FILLER_11_1957 ();
 sg13g2_fill_2 FILLER_11_1967 ();
 sg13g2_fill_1 FILLER_11_1969 ();
 sg13g2_fill_1 FILLER_11_1975 ();
 sg13g2_decap_8 FILLER_11_1980 ();
 sg13g2_decap_8 FILLER_11_1987 ();
 sg13g2_fill_2 FILLER_11_1994 ();
 sg13g2_fill_1 FILLER_11_2017 ();
 sg13g2_fill_2 FILLER_11_2048 ();
 sg13g2_decap_8 FILLER_11_2080 ();
 sg13g2_decap_8 FILLER_11_2087 ();
 sg13g2_decap_4 FILLER_11_2094 ();
 sg13g2_fill_2 FILLER_11_2102 ();
 sg13g2_decap_4 FILLER_11_2117 ();
 sg13g2_fill_2 FILLER_11_2134 ();
 sg13g2_fill_1 FILLER_11_2136 ();
 sg13g2_fill_1 FILLER_11_2146 ();
 sg13g2_decap_8 FILLER_11_2179 ();
 sg13g2_decap_8 FILLER_11_2196 ();
 sg13g2_decap_4 FILLER_11_2203 ();
 sg13g2_fill_2 FILLER_11_2207 ();
 sg13g2_fill_2 FILLER_11_2218 ();
 sg13g2_fill_1 FILLER_11_2220 ();
 sg13g2_fill_1 FILLER_11_2234 ();
 sg13g2_decap_4 FILLER_11_2272 ();
 sg13g2_fill_1 FILLER_11_2276 ();
 sg13g2_fill_2 FILLER_11_2294 ();
 sg13g2_fill_1 FILLER_11_2296 ();
 sg13g2_fill_1 FILLER_11_2319 ();
 sg13g2_fill_2 FILLER_11_2325 ();
 sg13g2_fill_1 FILLER_11_2327 ();
 sg13g2_decap_8 FILLER_11_2332 ();
 sg13g2_decap_4 FILLER_11_2339 ();
 sg13g2_fill_2 FILLER_11_2347 ();
 sg13g2_fill_2 FILLER_11_2369 ();
 sg13g2_decap_4 FILLER_11_2392 ();
 sg13g2_fill_1 FILLER_11_2396 ();
 sg13g2_decap_8 FILLER_11_2452 ();
 sg13g2_fill_1 FILLER_11_2459 ();
 sg13g2_decap_8 FILLER_11_2472 ();
 sg13g2_decap_8 FILLER_11_2479 ();
 sg13g2_decap_4 FILLER_11_2486 ();
 sg13g2_fill_1 FILLER_11_2499 ();
 sg13g2_fill_2 FILLER_11_2504 ();
 sg13g2_fill_1 FILLER_11_2515 ();
 sg13g2_fill_1 FILLER_11_2547 ();
 sg13g2_fill_1 FILLER_11_2557 ();
 sg13g2_fill_1 FILLER_11_2584 ();
 sg13g2_fill_1 FILLER_11_2619 ();
 sg13g2_fill_1 FILLER_11_2625 ();
 sg13g2_decap_4 FILLER_11_2639 ();
 sg13g2_fill_2 FILLER_11_2643 ();
 sg13g2_decap_4 FILLER_11_2649 ();
 sg13g2_fill_2 FILLER_11_2653 ();
 sg13g2_decap_4 FILLER_11_2668 ();
 sg13g2_fill_1 FILLER_11_2672 ();
 sg13g2_decap_8 FILLER_11_2694 ();
 sg13g2_decap_8 FILLER_11_2705 ();
 sg13g2_decap_8 FILLER_11_2712 ();
 sg13g2_fill_2 FILLER_11_2726 ();
 sg13g2_decap_8 FILLER_11_2741 ();
 sg13g2_fill_1 FILLER_11_2748 ();
 sg13g2_fill_1 FILLER_11_2801 ();
 sg13g2_fill_2 FILLER_11_2827 ();
 sg13g2_fill_1 FILLER_11_2834 ();
 sg13g2_decap_4 FILLER_11_2865 ();
 sg13g2_fill_1 FILLER_11_2869 ();
 sg13g2_decap_8 FILLER_11_2879 ();
 sg13g2_fill_2 FILLER_11_2886 ();
 sg13g2_fill_1 FILLER_11_2888 ();
 sg13g2_decap_8 FILLER_11_2902 ();
 sg13g2_decap_4 FILLER_11_2909 ();
 sg13g2_fill_1 FILLER_11_2913 ();
 sg13g2_fill_2 FILLER_11_2919 ();
 sg13g2_fill_2 FILLER_11_2926 ();
 sg13g2_fill_2 FILLER_11_2938 ();
 sg13g2_decap_8 FILLER_11_2971 ();
 sg13g2_fill_1 FILLER_11_2978 ();
 sg13g2_decap_4 FILLER_11_2983 ();
 sg13g2_fill_2 FILLER_11_2987 ();
 sg13g2_decap_4 FILLER_11_3002 ();
 sg13g2_decap_4 FILLER_11_3014 ();
 sg13g2_decap_4 FILLER_11_3036 ();
 sg13g2_fill_2 FILLER_11_3040 ();
 sg13g2_fill_1 FILLER_11_3054 ();
 sg13g2_fill_2 FILLER_11_3064 ();
 sg13g2_fill_2 FILLER_11_3075 ();
 sg13g2_decap_8 FILLER_11_3081 ();
 sg13g2_decap_8 FILLER_11_3088 ();
 sg13g2_decap_8 FILLER_11_3141 ();
 sg13g2_fill_2 FILLER_11_3148 ();
 sg13g2_fill_1 FILLER_11_3154 ();
 sg13g2_fill_1 FILLER_11_3163 ();
 sg13g2_fill_1 FILLER_11_3177 ();
 sg13g2_decap_8 FILLER_11_3182 ();
 sg13g2_decap_4 FILLER_11_3189 ();
 sg13g2_decap_4 FILLER_11_3197 ();
 sg13g2_fill_1 FILLER_11_3201 ();
 sg13g2_fill_2 FILLER_11_3211 ();
 sg13g2_fill_2 FILLER_11_3258 ();
 sg13g2_fill_2 FILLER_11_3279 ();
 sg13g2_fill_1 FILLER_11_3281 ();
 sg13g2_decap_4 FILLER_11_3299 ();
 sg13g2_fill_1 FILLER_11_3337 ();
 sg13g2_fill_2 FILLER_11_3364 ();
 sg13g2_decap_8 FILLER_11_3404 ();
 sg13g2_fill_2 FILLER_11_3411 ();
 sg13g2_fill_1 FILLER_11_3413 ();
 sg13g2_fill_1 FILLER_11_3418 ();
 sg13g2_fill_2 FILLER_11_3424 ();
 sg13g2_decap_4 FILLER_11_3462 ();
 sg13g2_fill_2 FILLER_11_3466 ();
 sg13g2_decap_4 FILLER_11_3499 ();
 sg13g2_fill_2 FILLER_11_3534 ();
 sg13g2_fill_1 FILLER_11_3536 ();
 sg13g2_decap_4 FILLER_11_3576 ();
 sg13g2_fill_1 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_97 ();
 sg13g2_decap_8 FILLER_12_104 ();
 sg13g2_decap_4 FILLER_12_111 ();
 sg13g2_fill_1 FILLER_12_115 ();
 sg13g2_decap_8 FILLER_12_124 ();
 sg13g2_fill_2 FILLER_12_131 ();
 sg13g2_fill_1 FILLER_12_160 ();
 sg13g2_fill_1 FILLER_12_175 ();
 sg13g2_decap_4 FILLER_12_226 ();
 sg13g2_fill_2 FILLER_12_284 ();
 sg13g2_fill_1 FILLER_12_286 ();
 sg13g2_fill_1 FILLER_12_296 ();
 sg13g2_decap_4 FILLER_12_316 ();
 sg13g2_fill_1 FILLER_12_320 ();
 sg13g2_decap_4 FILLER_12_340 ();
 sg13g2_fill_1 FILLER_12_344 ();
 sg13g2_decap_8 FILLER_12_358 ();
 sg13g2_decap_8 FILLER_12_365 ();
 sg13g2_decap_4 FILLER_12_412 ();
 sg13g2_fill_2 FILLER_12_416 ();
 sg13g2_fill_2 FILLER_12_444 ();
 sg13g2_fill_1 FILLER_12_446 ();
 sg13g2_fill_1 FILLER_12_461 ();
 sg13g2_fill_1 FILLER_12_493 ();
 sg13g2_fill_1 FILLER_12_521 ();
 sg13g2_fill_2 FILLER_12_532 ();
 sg13g2_decap_4 FILLER_12_580 ();
 sg13g2_fill_2 FILLER_12_584 ();
 sg13g2_decap_8 FILLER_12_590 ();
 sg13g2_decap_8 FILLER_12_597 ();
 sg13g2_decap_8 FILLER_12_604 ();
 sg13g2_fill_1 FILLER_12_611 ();
 sg13g2_fill_2 FILLER_12_616 ();
 sg13g2_fill_2 FILLER_12_636 ();
 sg13g2_fill_1 FILLER_12_638 ();
 sg13g2_fill_2 FILLER_12_721 ();
 sg13g2_decap_4 FILLER_12_728 ();
 sg13g2_fill_2 FILLER_12_732 ();
 sg13g2_decap_4 FILLER_12_742 ();
 sg13g2_fill_1 FILLER_12_809 ();
 sg13g2_fill_2 FILLER_12_823 ();
 sg13g2_fill_1 FILLER_12_825 ();
 sg13g2_fill_2 FILLER_12_841 ();
 sg13g2_fill_1 FILLER_12_843 ();
 sg13g2_fill_1 FILLER_12_854 ();
 sg13g2_decap_4 FILLER_12_886 ();
 sg13g2_decap_8 FILLER_12_926 ();
 sg13g2_decap_8 FILLER_12_933 ();
 sg13g2_decap_4 FILLER_12_948 ();
 sg13g2_fill_2 FILLER_12_952 ();
 sg13g2_decap_8 FILLER_12_989 ();
 sg13g2_fill_2 FILLER_12_996 ();
 sg13g2_fill_2 FILLER_12_1016 ();
 sg13g2_decap_4 FILLER_12_1039 ();
 sg13g2_decap_8 FILLER_12_1047 ();
 sg13g2_fill_1 FILLER_12_1054 ();
 sg13g2_fill_2 FILLER_12_1064 ();
 sg13g2_decap_4 FILLER_12_1083 ();
 sg13g2_fill_1 FILLER_12_1087 ();
 sg13g2_fill_2 FILLER_12_1092 ();
 sg13g2_fill_1 FILLER_12_1094 ();
 sg13g2_fill_1 FILLER_12_1099 ();
 sg13g2_fill_2 FILLER_12_1109 ();
 sg13g2_fill_2 FILLER_12_1128 ();
 sg13g2_fill_2 FILLER_12_1138 ();
 sg13g2_fill_1 FILLER_12_1145 ();
 sg13g2_fill_2 FILLER_12_1191 ();
 sg13g2_fill_1 FILLER_12_1210 ();
 sg13g2_decap_4 FILLER_12_1227 ();
 sg13g2_fill_2 FILLER_12_1231 ();
 sg13g2_fill_2 FILLER_12_1241 ();
 sg13g2_decap_8 FILLER_12_1251 ();
 sg13g2_decap_4 FILLER_12_1266 ();
 sg13g2_decap_4 FILLER_12_1278 ();
 sg13g2_fill_1 FILLER_12_1282 ();
 sg13g2_fill_2 FILLER_12_1291 ();
 sg13g2_fill_1 FILLER_12_1293 ();
 sg13g2_decap_4 FILLER_12_1302 ();
 sg13g2_fill_1 FILLER_12_1306 ();
 sg13g2_decap_8 FILLER_12_1354 ();
 sg13g2_fill_1 FILLER_12_1361 ();
 sg13g2_decap_4 FILLER_12_1379 ();
 sg13g2_fill_1 FILLER_12_1392 ();
 sg13g2_decap_4 FILLER_12_1414 ();
 sg13g2_decap_4 FILLER_12_1437 ();
 sg13g2_fill_2 FILLER_12_1441 ();
 sg13g2_fill_2 FILLER_12_1469 ();
 sg13g2_fill_1 FILLER_12_1471 ();
 sg13g2_fill_2 FILLER_12_1498 ();
 sg13g2_fill_1 FILLER_12_1500 ();
 sg13g2_decap_4 FILLER_12_1524 ();
 sg13g2_fill_1 FILLER_12_1528 ();
 sg13g2_decap_4 FILLER_12_1548 ();
 sg13g2_fill_2 FILLER_12_1552 ();
 sg13g2_decap_8 FILLER_12_1567 ();
 sg13g2_decap_8 FILLER_12_1574 ();
 sg13g2_decap_4 FILLER_12_1581 ();
 sg13g2_fill_1 FILLER_12_1585 ();
 sg13g2_fill_2 FILLER_12_1592 ();
 sg13g2_fill_1 FILLER_12_1594 ();
 sg13g2_decap_8 FILLER_12_1603 ();
 sg13g2_decap_4 FILLER_12_1610 ();
 sg13g2_decap_8 FILLER_12_1626 ();
 sg13g2_fill_2 FILLER_12_1633 ();
 sg13g2_fill_2 FILLER_12_1640 ();
 sg13g2_decap_4 FILLER_12_1660 ();
 sg13g2_fill_2 FILLER_12_1668 ();
 sg13g2_fill_1 FILLER_12_1670 ();
 sg13g2_decap_4 FILLER_12_1675 ();
 sg13g2_fill_2 FILLER_12_1679 ();
 sg13g2_decap_8 FILLER_12_1693 ();
 sg13g2_decap_8 FILLER_12_1700 ();
 sg13g2_decap_4 FILLER_12_1707 ();
 sg13g2_fill_1 FILLER_12_1711 ();
 sg13g2_decap_8 FILLER_12_1754 ();
 sg13g2_decap_8 FILLER_12_1761 ();
 sg13g2_decap_8 FILLER_12_1768 ();
 sg13g2_fill_2 FILLER_12_1775 ();
 sg13g2_fill_1 FILLER_12_1777 ();
 sg13g2_decap_4 FILLER_12_1786 ();
 sg13g2_fill_1 FILLER_12_1790 ();
 sg13g2_decap_8 FILLER_12_1801 ();
 sg13g2_decap_8 FILLER_12_1808 ();
 sg13g2_fill_1 FILLER_12_1828 ();
 sg13g2_decap_8 FILLER_12_1837 ();
 sg13g2_fill_2 FILLER_12_1844 ();
 sg13g2_fill_1 FILLER_12_1850 ();
 sg13g2_fill_2 FILLER_12_1856 ();
 sg13g2_decap_4 FILLER_12_1880 ();
 sg13g2_fill_2 FILLER_12_1884 ();
 sg13g2_fill_2 FILLER_12_1890 ();
 sg13g2_fill_1 FILLER_12_1892 ();
 sg13g2_fill_1 FILLER_12_1898 ();
 sg13g2_fill_1 FILLER_12_1944 ();
 sg13g2_fill_2 FILLER_12_1958 ();
 sg13g2_fill_2 FILLER_12_1968 ();
 sg13g2_fill_1 FILLER_12_1970 ();
 sg13g2_decap_4 FILLER_12_1997 ();
 sg13g2_fill_1 FILLER_12_2001 ();
 sg13g2_fill_2 FILLER_12_2005 ();
 sg13g2_decap_4 FILLER_12_2015 ();
 sg13g2_fill_2 FILLER_12_2019 ();
 sg13g2_decap_4 FILLER_12_2038 ();
 sg13g2_fill_1 FILLER_12_2042 ();
 sg13g2_decap_4 FILLER_12_2048 ();
 sg13g2_fill_2 FILLER_12_2052 ();
 sg13g2_fill_2 FILLER_12_2058 ();
 sg13g2_fill_1 FILLER_12_2060 ();
 sg13g2_fill_2 FILLER_12_2074 ();
 sg13g2_decap_4 FILLER_12_2087 ();
 sg13g2_fill_1 FILLER_12_2091 ();
 sg13g2_fill_2 FILLER_12_2111 ();
 sg13g2_fill_1 FILLER_12_2113 ();
 sg13g2_decap_8 FILLER_12_2119 ();
 sg13g2_decap_4 FILLER_12_2126 ();
 sg13g2_fill_2 FILLER_12_2156 ();
 sg13g2_fill_1 FILLER_12_2158 ();
 sg13g2_fill_2 FILLER_12_2163 ();
 sg13g2_fill_1 FILLER_12_2165 ();
 sg13g2_decap_8 FILLER_12_2174 ();
 sg13g2_decap_4 FILLER_12_2181 ();
 sg13g2_fill_2 FILLER_12_2185 ();
 sg13g2_fill_2 FILLER_12_2197 ();
 sg13g2_fill_1 FILLER_12_2199 ();
 sg13g2_fill_2 FILLER_12_2229 ();
 sg13g2_fill_1 FILLER_12_2231 ();
 sg13g2_fill_2 FILLER_12_2258 ();
 sg13g2_fill_1 FILLER_12_2260 ();
 sg13g2_decap_4 FILLER_12_2312 ();
 sg13g2_fill_1 FILLER_12_2316 ();
 sg13g2_decap_4 FILLER_12_2356 ();
 sg13g2_fill_1 FILLER_12_2360 ();
 sg13g2_decap_4 FILLER_12_2369 ();
 sg13g2_fill_2 FILLER_12_2373 ();
 sg13g2_fill_2 FILLER_12_2380 ();
 sg13g2_fill_1 FILLER_12_2382 ();
 sg13g2_fill_2 FILLER_12_2413 ();
 sg13g2_fill_2 FILLER_12_2429 ();
 sg13g2_fill_1 FILLER_12_2431 ();
 sg13g2_fill_2 FILLER_12_2447 ();
 sg13g2_fill_2 FILLER_12_2454 ();
 sg13g2_fill_1 FILLER_12_2456 ();
 sg13g2_fill_2 FILLER_12_2465 ();
 sg13g2_fill_1 FILLER_12_2467 ();
 sg13g2_decap_4 FILLER_12_2476 ();
 sg13g2_fill_1 FILLER_12_2480 ();
 sg13g2_decap_8 FILLER_12_2507 ();
 sg13g2_fill_1 FILLER_12_2514 ();
 sg13g2_decap_8 FILLER_12_2519 ();
 sg13g2_fill_1 FILLER_12_2526 ();
 sg13g2_fill_2 FILLER_12_2553 ();
 sg13g2_decap_4 FILLER_12_2568 ();
 sg13g2_fill_2 FILLER_12_2576 ();
 sg13g2_fill_1 FILLER_12_2578 ();
 sg13g2_fill_2 FILLER_12_2592 ();
 sg13g2_decap_8 FILLER_12_2611 ();
 sg13g2_decap_8 FILLER_12_2618 ();
 sg13g2_decap_8 FILLER_12_2625 ();
 sg13g2_decap_4 FILLER_12_2632 ();
 sg13g2_fill_1 FILLER_12_2636 ();
 sg13g2_fill_2 FILLER_12_2672 ();
 sg13g2_decap_8 FILLER_12_2741 ();
 sg13g2_decap_4 FILLER_12_2748 ();
 sg13g2_fill_1 FILLER_12_2752 ();
 sg13g2_fill_2 FILLER_12_2783 ();
 sg13g2_decap_4 FILLER_12_2811 ();
 sg13g2_fill_1 FILLER_12_2815 ();
 sg13g2_decap_4 FILLER_12_2821 ();
 sg13g2_fill_1 FILLER_12_2825 ();
 sg13g2_fill_2 FILLER_12_2892 ();
 sg13g2_fill_1 FILLER_12_2894 ();
 sg13g2_decap_8 FILLER_12_2903 ();
 sg13g2_decap_4 FILLER_12_2910 ();
 sg13g2_fill_1 FILLER_12_2914 ();
 sg13g2_fill_1 FILLER_12_2930 ();
 sg13g2_decap_8 FILLER_12_2941 ();
 sg13g2_fill_2 FILLER_12_2948 ();
 sg13g2_fill_1 FILLER_12_2950 ();
 sg13g2_decap_8 FILLER_12_2959 ();
 sg13g2_fill_2 FILLER_12_2966 ();
 sg13g2_fill_2 FILLER_12_2972 ();
 sg13g2_fill_1 FILLER_12_2974 ();
 sg13g2_fill_1 FILLER_12_2979 ();
 sg13g2_fill_2 FILLER_12_2997 ();
 sg13g2_fill_1 FILLER_12_2999 ();
 sg13g2_decap_8 FILLER_12_3017 ();
 sg13g2_decap_4 FILLER_12_3024 ();
 sg13g2_fill_2 FILLER_12_3038 ();
 sg13g2_fill_1 FILLER_12_3040 ();
 sg13g2_fill_2 FILLER_12_3057 ();
 sg13g2_fill_1 FILLER_12_3059 ();
 sg13g2_decap_4 FILLER_12_3091 ();
 sg13g2_fill_2 FILLER_12_3095 ();
 sg13g2_fill_2 FILLER_12_3102 ();
 sg13g2_fill_1 FILLER_12_3104 ();
 sg13g2_fill_2 FILLER_12_3114 ();
 sg13g2_fill_2 FILLER_12_3201 ();
 sg13g2_fill_1 FILLER_12_3203 ();
 sg13g2_decap_8 FILLER_12_3218 ();
 sg13g2_fill_1 FILLER_12_3225 ();
 sg13g2_fill_1 FILLER_12_3263 ();
 sg13g2_decap_8 FILLER_12_3295 ();
 sg13g2_decap_4 FILLER_12_3302 ();
 sg13g2_decap_8 FILLER_12_3314 ();
 sg13g2_decap_4 FILLER_12_3325 ();
 sg13g2_fill_1 FILLER_12_3329 ();
 sg13g2_fill_2 FILLER_12_3343 ();
 sg13g2_decap_8 FILLER_12_3354 ();
 sg13g2_decap_4 FILLER_12_3361 ();
 sg13g2_fill_2 FILLER_12_3365 ();
 sg13g2_decap_8 FILLER_12_3375 ();
 sg13g2_decap_8 FILLER_12_3382 ();
 sg13g2_fill_1 FILLER_12_3389 ();
 sg13g2_decap_4 FILLER_12_3408 ();
 sg13g2_fill_1 FILLER_12_3412 ();
 sg13g2_fill_2 FILLER_12_3439 ();
 sg13g2_decap_4 FILLER_12_3469 ();
 sg13g2_decap_4 FILLER_12_3483 ();
 sg13g2_fill_2 FILLER_12_3487 ();
 sg13g2_decap_8 FILLER_12_3497 ();
 sg13g2_fill_1 FILLER_12_3504 ();
 sg13g2_fill_2 FILLER_12_3510 ();
 sg13g2_fill_2 FILLER_12_3517 ();
 sg13g2_fill_2 FILLER_12_3533 ();
 sg13g2_fill_1 FILLER_12_3535 ();
 sg13g2_fill_1 FILLER_12_3553 ();
 sg13g2_decap_4 FILLER_13_36 ();
 sg13g2_fill_1 FILLER_13_58 ();
 sg13g2_decap_4 FILLER_13_63 ();
 sg13g2_fill_1 FILLER_13_67 ();
 sg13g2_fill_1 FILLER_13_108 ();
 sg13g2_fill_2 FILLER_13_155 ();
 sg13g2_fill_1 FILLER_13_157 ();
 sg13g2_fill_2 FILLER_13_222 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_4 FILLER_13_245 ();
 sg13g2_fill_2 FILLER_13_249 ();
 sg13g2_fill_1 FILLER_13_265 ();
 sg13g2_fill_1 FILLER_13_285 ();
 sg13g2_fill_2 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_390 ();
 sg13g2_decap_8 FILLER_13_409 ();
 sg13g2_fill_1 FILLER_13_416 ();
 sg13g2_fill_2 FILLER_13_480 ();
 sg13g2_decap_8 FILLER_13_494 ();
 sg13g2_decap_4 FILLER_13_501 ();
 sg13g2_decap_8 FILLER_13_513 ();
 sg13g2_decap_8 FILLER_13_525 ();
 sg13g2_decap_4 FILLER_13_532 ();
 sg13g2_fill_1 FILLER_13_536 ();
 sg13g2_decap_8 FILLER_13_541 ();
 sg13g2_decap_8 FILLER_13_556 ();
 sg13g2_fill_2 FILLER_13_563 ();
 sg13g2_decap_8 FILLER_13_569 ();
 sg13g2_fill_2 FILLER_13_576 ();
 sg13g2_fill_1 FILLER_13_578 ();
 sg13g2_fill_2 FILLER_13_584 ();
 sg13g2_decap_4 FILLER_13_612 ();
 sg13g2_fill_1 FILLER_13_616 ();
 sg13g2_fill_2 FILLER_13_661 ();
 sg13g2_fill_1 FILLER_13_668 ();
 sg13g2_fill_2 FILLER_13_683 ();
 sg13g2_fill_1 FILLER_13_685 ();
 sg13g2_fill_1 FILLER_13_690 ();
 sg13g2_fill_1 FILLER_13_696 ();
 sg13g2_decap_8 FILLER_13_705 ();
 sg13g2_decap_8 FILLER_13_712 ();
 sg13g2_decap_4 FILLER_13_719 ();
 sg13g2_fill_2 FILLER_13_767 ();
 sg13g2_fill_1 FILLER_13_769 ();
 sg13g2_decap_8 FILLER_13_779 ();
 sg13g2_decap_4 FILLER_13_786 ();
 sg13g2_fill_1 FILLER_13_799 ();
 sg13g2_decap_8 FILLER_13_804 ();
 sg13g2_fill_1 FILLER_13_820 ();
 sg13g2_decap_8 FILLER_13_830 ();
 sg13g2_fill_1 FILLER_13_837 ();
 sg13g2_fill_2 FILLER_13_841 ();
 sg13g2_decap_8 FILLER_13_847 ();
 sg13g2_fill_2 FILLER_13_854 ();
 sg13g2_fill_1 FILLER_13_874 ();
 sg13g2_fill_1 FILLER_13_883 ();
 sg13g2_decap_8 FILLER_13_897 ();
 sg13g2_fill_2 FILLER_13_904 ();
 sg13g2_decap_4 FILLER_13_910 ();
 sg13g2_fill_2 FILLER_13_914 ();
 sg13g2_decap_4 FILLER_13_931 ();
 sg13g2_fill_1 FILLER_13_935 ();
 sg13g2_fill_2 FILLER_13_941 ();
 sg13g2_fill_1 FILLER_13_943 ();
 sg13g2_fill_2 FILLER_13_952 ();
 sg13g2_fill_1 FILLER_13_954 ();
 sg13g2_decap_8 FILLER_13_963 ();
 sg13g2_decap_4 FILLER_13_970 ();
 sg13g2_fill_2 FILLER_13_978 ();
 sg13g2_fill_1 FILLER_13_980 ();
 sg13g2_decap_8 FILLER_13_986 ();
 sg13g2_decap_4 FILLER_13_1004 ();
 sg13g2_fill_1 FILLER_13_1008 ();
 sg13g2_fill_2 FILLER_13_1018 ();
 sg13g2_fill_2 FILLER_13_1029 ();
 sg13g2_fill_1 FILLER_13_1031 ();
 sg13g2_fill_1 FILLER_13_1066 ();
 sg13g2_decap_8 FILLER_13_1088 ();
 sg13g2_fill_1 FILLER_13_1095 ();
 sg13g2_fill_2 FILLER_13_1101 ();
 sg13g2_fill_1 FILLER_13_1103 ();
 sg13g2_fill_2 FILLER_13_1134 ();
 sg13g2_decap_8 FILLER_13_1141 ();
 sg13g2_decap_8 FILLER_13_1148 ();
 sg13g2_fill_2 FILLER_13_1164 ();
 sg13g2_fill_1 FILLER_13_1171 ();
 sg13g2_decap_8 FILLER_13_1180 ();
 sg13g2_decap_4 FILLER_13_1187 ();
 sg13g2_decap_8 FILLER_13_1195 ();
 sg13g2_decap_4 FILLER_13_1202 ();
 sg13g2_fill_2 FILLER_13_1214 ();
 sg13g2_fill_1 FILLER_13_1220 ();
 sg13g2_decap_4 FILLER_13_1233 ();
 sg13g2_decap_4 FILLER_13_1241 ();
 sg13g2_fill_1 FILLER_13_1245 ();
 sg13g2_fill_2 FILLER_13_1256 ();
 sg13g2_fill_1 FILLER_13_1298 ();
 sg13g2_decap_8 FILLER_13_1303 ();
 sg13g2_decap_4 FILLER_13_1310 ();
 sg13g2_fill_1 FILLER_13_1314 ();
 sg13g2_fill_1 FILLER_13_1328 ();
 sg13g2_fill_2 FILLER_13_1358 ();
 sg13g2_fill_1 FILLER_13_1360 ();
 sg13g2_fill_2 FILLER_13_1366 ();
 sg13g2_fill_1 FILLER_13_1368 ();
 sg13g2_decap_4 FILLER_13_1382 ();
 sg13g2_fill_2 FILLER_13_1386 ();
 sg13g2_decap_4 FILLER_13_1406 ();
 sg13g2_fill_1 FILLER_13_1410 ();
 sg13g2_decap_8 FILLER_13_1415 ();
 sg13g2_fill_2 FILLER_13_1422 ();
 sg13g2_fill_1 FILLER_13_1424 ();
 sg13g2_fill_2 FILLER_13_1434 ();
 sg13g2_fill_1 FILLER_13_1436 ();
 sg13g2_decap_4 FILLER_13_1450 ();
 sg13g2_decap_4 FILLER_13_1458 ();
 sg13g2_fill_1 FILLER_13_1462 ();
 sg13g2_decap_8 FILLER_13_1472 ();
 sg13g2_decap_4 FILLER_13_1483 ();
 sg13g2_fill_2 FILLER_13_1487 ();
 sg13g2_fill_2 FILLER_13_1497 ();
 sg13g2_fill_1 FILLER_13_1499 ();
 sg13g2_decap_8 FILLER_13_1521 ();
 sg13g2_decap_8 FILLER_13_1528 ();
 sg13g2_decap_8 FILLER_13_1535 ();
 sg13g2_fill_1 FILLER_13_1556 ();
 sg13g2_decap_8 FILLER_13_1562 ();
 sg13g2_decap_4 FILLER_13_1569 ();
 sg13g2_fill_1 FILLER_13_1573 ();
 sg13g2_decap_8 FILLER_13_1579 ();
 sg13g2_fill_1 FILLER_13_1599 ();
 sg13g2_fill_1 FILLER_13_1610 ();
 sg13g2_decap_4 FILLER_13_1624 ();
 sg13g2_fill_1 FILLER_13_1633 ();
 sg13g2_fill_2 FILLER_13_1648 ();
 sg13g2_fill_2 FILLER_13_1659 ();
 sg13g2_fill_1 FILLER_13_1661 ();
 sg13g2_fill_2 FILLER_13_1671 ();
 sg13g2_fill_1 FILLER_13_1673 ();
 sg13g2_fill_1 FILLER_13_1719 ();
 sg13g2_decap_8 FILLER_13_1728 ();
 sg13g2_fill_2 FILLER_13_1735 ();
 sg13g2_fill_1 FILLER_13_1737 ();
 sg13g2_decap_8 FILLER_13_1742 ();
 sg13g2_decap_4 FILLER_13_1749 ();
 sg13g2_fill_1 FILLER_13_1753 ();
 sg13g2_decap_8 FILLER_13_1806 ();
 sg13g2_decap_4 FILLER_13_1844 ();
 sg13g2_fill_1 FILLER_13_1861 ();
 sg13g2_decap_8 FILLER_13_1871 ();
 sg13g2_decap_4 FILLER_13_1878 ();
 sg13g2_fill_1 FILLER_13_1908 ();
 sg13g2_fill_2 FILLER_13_1923 ();
 sg13g2_fill_1 FILLER_13_1925 ();
 sg13g2_decap_4 FILLER_13_1929 ();
 sg13g2_fill_1 FILLER_13_1960 ();
 sg13g2_fill_2 FILLER_13_1990 ();
 sg13g2_decap_4 FILLER_13_2000 ();
 sg13g2_decap_8 FILLER_13_2017 ();
 sg13g2_fill_2 FILLER_13_2024 ();
 sg13g2_fill_1 FILLER_13_2026 ();
 sg13g2_fill_1 FILLER_13_2035 ();
 sg13g2_decap_4 FILLER_13_2045 ();
 sg13g2_fill_2 FILLER_13_2063 ();
 sg13g2_fill_1 FILLER_13_2124 ();
 sg13g2_fill_1 FILLER_13_2151 ();
 sg13g2_fill_2 FILLER_13_2161 ();
 sg13g2_fill_1 FILLER_13_2163 ();
 sg13g2_decap_8 FILLER_13_2174 ();
 sg13g2_decap_4 FILLER_13_2181 ();
 sg13g2_fill_1 FILLER_13_2185 ();
 sg13g2_decap_8 FILLER_13_2194 ();
 sg13g2_decap_8 FILLER_13_2201 ();
 sg13g2_fill_1 FILLER_13_2216 ();
 sg13g2_decap_4 FILLER_13_2230 ();
 sg13g2_fill_1 FILLER_13_2234 ();
 sg13g2_decap_8 FILLER_13_2272 ();
 sg13g2_decap_8 FILLER_13_2287 ();
 sg13g2_decap_4 FILLER_13_2303 ();
 sg13g2_fill_1 FILLER_13_2307 ();
 sg13g2_decap_8 FILLER_13_2316 ();
 sg13g2_decap_8 FILLER_13_2323 ();
 sg13g2_decap_4 FILLER_13_2330 ();
 sg13g2_fill_2 FILLER_13_2373 ();
 sg13g2_fill_1 FILLER_13_2375 ();
 sg13g2_decap_4 FILLER_13_2387 ();
 sg13g2_fill_1 FILLER_13_2391 ();
 sg13g2_fill_2 FILLER_13_2438 ();
 sg13g2_decap_4 FILLER_13_2444 ();
 sg13g2_fill_1 FILLER_13_2478 ();
 sg13g2_fill_2 FILLER_13_2488 ();
 sg13g2_fill_1 FILLER_13_2490 ();
 sg13g2_decap_8 FILLER_13_2531 ();
 sg13g2_fill_2 FILLER_13_2538 ();
 sg13g2_fill_1 FILLER_13_2540 ();
 sg13g2_decap_4 FILLER_13_2554 ();
 sg13g2_fill_1 FILLER_13_2558 ();
 sg13g2_decap_4 FILLER_13_2577 ();
 sg13g2_fill_1 FILLER_13_2581 ();
 sg13g2_fill_2 FILLER_13_2592 ();
 sg13g2_fill_1 FILLER_13_2594 ();
 sg13g2_decap_4 FILLER_13_2631 ();
 sg13g2_decap_8 FILLER_13_2640 ();
 sg13g2_decap_4 FILLER_13_2647 ();
 sg13g2_fill_1 FILLER_13_2651 ();
 sg13g2_fill_2 FILLER_13_2660 ();
 sg13g2_fill_1 FILLER_13_2662 ();
 sg13g2_decap_8 FILLER_13_2671 ();
 sg13g2_decap_8 FILLER_13_2678 ();
 sg13g2_decap_4 FILLER_13_2685 ();
 sg13g2_fill_2 FILLER_13_2689 ();
 sg13g2_fill_1 FILLER_13_2696 ();
 sg13g2_fill_1 FILLER_13_2705 ();
 sg13g2_fill_1 FILLER_13_2732 ();
 sg13g2_fill_1 FILLER_13_2754 ();
 sg13g2_fill_1 FILLER_13_2786 ();
 sg13g2_fill_1 FILLER_13_2797 ();
 sg13g2_decap_4 FILLER_13_2803 ();
 sg13g2_decap_4 FILLER_13_2816 ();
 sg13g2_fill_1 FILLER_13_2820 ();
 sg13g2_decap_4 FILLER_13_2833 ();
 sg13g2_fill_2 FILLER_13_2847 ();
 sg13g2_decap_8 FILLER_13_2858 ();
 sg13g2_decap_4 FILLER_13_2865 ();
 sg13g2_fill_1 FILLER_13_2869 ();
 sg13g2_decap_4 FILLER_13_2874 ();
 sg13g2_fill_2 FILLER_13_2878 ();
 sg13g2_decap_8 FILLER_13_2884 ();
 sg13g2_decap_8 FILLER_13_2891 ();
 sg13g2_decap_4 FILLER_13_2898 ();
 sg13g2_fill_1 FILLER_13_2902 ();
 sg13g2_fill_1 FILLER_13_2926 ();
 sg13g2_fill_2 FILLER_13_2958 ();
 sg13g2_fill_2 FILLER_13_2991 ();
 sg13g2_fill_1 FILLER_13_2998 ();
 sg13g2_decap_8 FILLER_13_3063 ();
 sg13g2_decap_4 FILLER_13_3083 ();
 sg13g2_fill_1 FILLER_13_3087 ();
 sg13g2_decap_8 FILLER_13_3092 ();
 sg13g2_fill_2 FILLER_13_3099 ();
 sg13g2_fill_1 FILLER_13_3141 ();
 sg13g2_fill_2 FILLER_13_3147 ();
 sg13g2_fill_1 FILLER_13_3149 ();
 sg13g2_fill_1 FILLER_13_3158 ();
 sg13g2_decap_8 FILLER_13_3172 ();
 sg13g2_decap_8 FILLER_13_3179 ();
 sg13g2_fill_1 FILLER_13_3186 ();
 sg13g2_fill_1 FILLER_13_3229 ();
 sg13g2_fill_2 FILLER_13_3239 ();
 sg13g2_fill_1 FILLER_13_3241 ();
 sg13g2_decap_8 FILLER_13_3269 ();
 sg13g2_decap_4 FILLER_13_3276 ();
 sg13g2_fill_1 FILLER_13_3280 ();
 sg13g2_decap_8 FILLER_13_3290 ();
 sg13g2_decap_8 FILLER_13_3297 ();
 sg13g2_fill_1 FILLER_13_3304 ();
 sg13g2_decap_8 FILLER_13_3321 ();
 sg13g2_fill_2 FILLER_13_3328 ();
 sg13g2_fill_1 FILLER_13_3330 ();
 sg13g2_fill_1 FILLER_13_3335 ();
 sg13g2_fill_2 FILLER_13_3344 ();
 sg13g2_decap_4 FILLER_13_3350 ();
 sg13g2_fill_1 FILLER_13_3354 ();
 sg13g2_decap_8 FILLER_13_3381 ();
 sg13g2_decap_4 FILLER_13_3388 ();
 sg13g2_decap_8 FILLER_13_3410 ();
 sg13g2_fill_1 FILLER_13_3417 ();
 sg13g2_decap_8 FILLER_13_3435 ();
 sg13g2_fill_2 FILLER_13_3442 ();
 sg13g2_fill_2 FILLER_13_3502 ();
 sg13g2_fill_1 FILLER_13_3504 ();
 sg13g2_decap_4 FILLER_13_3561 ();
 sg13g2_fill_2 FILLER_13_3578 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_92 ();
 sg13g2_fill_2 FILLER_14_97 ();
 sg13g2_fill_1 FILLER_14_99 ();
 sg13g2_fill_1 FILLER_14_122 ();
 sg13g2_fill_1 FILLER_14_128 ();
 sg13g2_fill_2 FILLER_14_138 ();
 sg13g2_decap_4 FILLER_14_145 ();
 sg13g2_fill_1 FILLER_14_149 ();
 sg13g2_decap_8 FILLER_14_249 ();
 sg13g2_decap_8 FILLER_14_282 ();
 sg13g2_fill_2 FILLER_14_289 ();
 sg13g2_fill_1 FILLER_14_319 ();
 sg13g2_fill_2 FILLER_14_347 ();
 sg13g2_fill_1 FILLER_14_349 ();
 sg13g2_decap_8 FILLER_14_354 ();
 sg13g2_decap_8 FILLER_14_361 ();
 sg13g2_fill_2 FILLER_14_382 ();
 sg13g2_fill_1 FILLER_14_384 ();
 sg13g2_fill_2 FILLER_14_408 ();
 sg13g2_fill_1 FILLER_14_410 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_fill_1 FILLER_14_427 ();
 sg13g2_decap_8 FILLER_14_436 ();
 sg13g2_decap_4 FILLER_14_443 ();
 sg13g2_fill_1 FILLER_14_447 ();
 sg13g2_decap_8 FILLER_14_469 ();
 sg13g2_fill_2 FILLER_14_476 ();
 sg13g2_decap_8 FILLER_14_518 ();
 sg13g2_fill_1 FILLER_14_525 ();
 sg13g2_fill_2 FILLER_14_538 ();
 sg13g2_fill_1 FILLER_14_540 ();
 sg13g2_decap_4 FILLER_14_544 ();
 sg13g2_fill_2 FILLER_14_548 ();
 sg13g2_fill_2 FILLER_14_562 ();
 sg13g2_fill_1 FILLER_14_564 ();
 sg13g2_decap_4 FILLER_14_578 ();
 sg13g2_fill_1 FILLER_14_582 ();
 sg13g2_fill_2 FILLER_14_591 ();
 sg13g2_fill_1 FILLER_14_593 ();
 sg13g2_decap_8 FILLER_14_618 ();
 sg13g2_fill_2 FILLER_14_638 ();
 sg13g2_fill_1 FILLER_14_640 ();
 sg13g2_decap_4 FILLER_14_679 ();
 sg13g2_fill_1 FILLER_14_683 ();
 sg13g2_fill_2 FILLER_14_702 ();
 sg13g2_fill_1 FILLER_14_708 ();
 sg13g2_fill_2 FILLER_14_714 ();
 sg13g2_decap_8 FILLER_14_724 ();
 sg13g2_decap_4 FILLER_14_731 ();
 sg13g2_decap_8 FILLER_14_761 ();
 sg13g2_fill_1 FILLER_14_768 ();
 sg13g2_decap_4 FILLER_14_773 ();
 sg13g2_fill_1 FILLER_14_777 ();
 sg13g2_fill_2 FILLER_14_787 ();
 sg13g2_fill_1 FILLER_14_854 ();
 sg13g2_decap_4 FILLER_14_899 ();
 sg13g2_fill_2 FILLER_14_903 ();
 sg13g2_fill_2 FILLER_14_915 ();
 sg13g2_fill_2 FILLER_14_934 ();
 sg13g2_fill_1 FILLER_14_936 ();
 sg13g2_decap_4 FILLER_14_950 ();
 sg13g2_fill_2 FILLER_14_965 ();
 sg13g2_decap_8 FILLER_14_981 ();
 sg13g2_fill_2 FILLER_14_988 ();
 sg13g2_fill_1 FILLER_14_990 ();
 sg13g2_decap_4 FILLER_14_1033 ();
 sg13g2_fill_1 FILLER_14_1037 ();
 sg13g2_fill_2 FILLER_14_1047 ();
 sg13g2_fill_2 FILLER_14_1058 ();
 sg13g2_fill_1 FILLER_14_1060 ();
 sg13g2_decap_8 FILLER_14_1101 ();
 sg13g2_decap_4 FILLER_14_1108 ();
 sg13g2_decap_8 FILLER_14_1155 ();
 sg13g2_decap_4 FILLER_14_1162 ();
 sg13g2_fill_1 FILLER_14_1166 ();
 sg13g2_fill_2 FILLER_14_1198 ();
 sg13g2_decap_4 FILLER_14_1236 ();
 sg13g2_fill_2 FILLER_14_1250 ();
 sg13g2_fill_1 FILLER_14_1256 ();
 sg13g2_decap_8 FILLER_14_1276 ();
 sg13g2_decap_8 FILLER_14_1314 ();
 sg13g2_decap_4 FILLER_14_1321 ();
 sg13g2_decap_4 FILLER_14_1351 ();
 sg13g2_fill_1 FILLER_14_1355 ();
 sg13g2_fill_2 FILLER_14_1382 ();
 sg13g2_fill_1 FILLER_14_1384 ();
 sg13g2_fill_1 FILLER_14_1425 ();
 sg13g2_decap_8 FILLER_14_1452 ();
 sg13g2_fill_1 FILLER_14_1459 ();
 sg13g2_decap_8 FILLER_14_1495 ();
 sg13g2_decap_8 FILLER_14_1502 ();
 sg13g2_fill_2 FILLER_14_1519 ();
 sg13g2_fill_1 FILLER_14_1521 ();
 sg13g2_fill_2 FILLER_14_1535 ();
 sg13g2_fill_1 FILLER_14_1537 ();
 sg13g2_fill_2 FILLER_14_1554 ();
 sg13g2_fill_1 FILLER_14_1556 ();
 sg13g2_decap_4 FILLER_14_1588 ();
 sg13g2_fill_1 FILLER_14_1592 ();
 sg13g2_decap_8 FILLER_14_1628 ();
 sg13g2_decap_4 FILLER_14_1684 ();
 sg13g2_fill_2 FILLER_14_1688 ();
 sg13g2_decap_8 FILLER_14_1694 ();
 sg13g2_decap_8 FILLER_14_1701 ();
 sg13g2_fill_2 FILLER_14_1708 ();
 sg13g2_fill_2 FILLER_14_1723 ();
 sg13g2_fill_1 FILLER_14_1725 ();
 sg13g2_decap_8 FILLER_14_1757 ();
 sg13g2_fill_1 FILLER_14_1764 ();
 sg13g2_decap_8 FILLER_14_1773 ();
 sg13g2_decap_8 FILLER_14_1785 ();
 sg13g2_fill_1 FILLER_14_1792 ();
 sg13g2_decap_8 FILLER_14_1805 ();
 sg13g2_decap_4 FILLER_14_1812 ();
 sg13g2_decap_8 FILLER_14_1821 ();
 sg13g2_fill_1 FILLER_14_1828 ();
 sg13g2_decap_8 FILLER_14_1833 ();
 sg13g2_fill_2 FILLER_14_1840 ();
 sg13g2_fill_1 FILLER_14_1842 ();
 sg13g2_decap_4 FILLER_14_1874 ();
 sg13g2_fill_2 FILLER_14_1906 ();
 sg13g2_fill_1 FILLER_14_1922 ();
 sg13g2_decap_4 FILLER_14_1935 ();
 sg13g2_fill_2 FILLER_14_1947 ();
 sg13g2_fill_2 FILLER_14_1974 ();
 sg13g2_fill_1 FILLER_14_1976 ();
 sg13g2_decap_4 FILLER_14_1991 ();
 sg13g2_fill_2 FILLER_14_2000 ();
 sg13g2_fill_1 FILLER_14_2006 ();
 sg13g2_fill_2 FILLER_14_2011 ();
 sg13g2_decap_4 FILLER_14_2070 ();
 sg13g2_fill_2 FILLER_14_2074 ();
 sg13g2_fill_1 FILLER_14_2079 ();
 sg13g2_decap_8 FILLER_14_2101 ();
 sg13g2_fill_1 FILLER_14_2113 ();
 sg13g2_fill_2 FILLER_14_2122 ();
 sg13g2_decap_8 FILLER_14_2137 ();
 sg13g2_fill_1 FILLER_14_2148 ();
 sg13g2_decap_8 FILLER_14_2176 ();
 sg13g2_decap_4 FILLER_14_2209 ();
 sg13g2_fill_2 FILLER_14_2222 ();
 sg13g2_fill_1 FILLER_14_2224 ();
 sg13g2_decap_8 FILLER_14_2233 ();
 sg13g2_fill_2 FILLER_14_2240 ();
 sg13g2_fill_1 FILLER_14_2242 ();
 sg13g2_decap_8 FILLER_14_2247 ();
 sg13g2_fill_1 FILLER_14_2259 ();
 sg13g2_fill_2 FILLER_14_2268 ();
 sg13g2_decap_8 FILLER_14_2278 ();
 sg13g2_fill_2 FILLER_14_2285 ();
 sg13g2_fill_1 FILLER_14_2287 ();
 sg13g2_fill_2 FILLER_14_2293 ();
 sg13g2_fill_1 FILLER_14_2295 ();
 sg13g2_decap_8 FILLER_14_2300 ();
 sg13g2_decap_8 FILLER_14_2307 ();
 sg13g2_fill_1 FILLER_14_2314 ();
 sg13g2_fill_1 FILLER_14_2345 ();
 sg13g2_fill_2 FILLER_14_2351 ();
 sg13g2_fill_1 FILLER_14_2353 ();
 sg13g2_fill_2 FILLER_14_2368 ();
 sg13g2_fill_1 FILLER_14_2370 ();
 sg13g2_decap_8 FILLER_14_2392 ();
 sg13g2_fill_2 FILLER_14_2399 ();
 sg13g2_decap_8 FILLER_14_2411 ();
 sg13g2_decap_4 FILLER_14_2418 ();
 sg13g2_fill_1 FILLER_14_2422 ();
 sg13g2_fill_1 FILLER_14_2427 ();
 sg13g2_decap_4 FILLER_14_2433 ();
 sg13g2_fill_1 FILLER_14_2437 ();
 sg13g2_decap_8 FILLER_14_2442 ();
 sg13g2_decap_8 FILLER_14_2449 ();
 sg13g2_fill_2 FILLER_14_2456 ();
 sg13g2_fill_1 FILLER_14_2458 ();
 sg13g2_decap_8 FILLER_14_2475 ();
 sg13g2_decap_8 FILLER_14_2482 ();
 sg13g2_fill_2 FILLER_14_2489 ();
 sg13g2_fill_2 FILLER_14_2500 ();
 sg13g2_fill_1 FILLER_14_2502 ();
 sg13g2_fill_2 FILLER_14_2516 ();
 sg13g2_decap_8 FILLER_14_2531 ();
 sg13g2_decap_8 FILLER_14_2551 ();
 sg13g2_fill_1 FILLER_14_2603 ();
 sg13g2_fill_1 FILLER_14_2639 ();
 sg13g2_decap_4 FILLER_14_2666 ();
 sg13g2_fill_2 FILLER_14_2723 ();
 sg13g2_decap_4 FILLER_14_2742 ();
 sg13g2_fill_1 FILLER_14_2754 ();
 sg13g2_decap_8 FILLER_14_2763 ();
 sg13g2_decap_4 FILLER_14_2770 ();
 sg13g2_fill_2 FILLER_14_2774 ();
 sg13g2_fill_2 FILLER_14_2789 ();
 sg13g2_decap_8 FILLER_14_2800 ();
 sg13g2_fill_2 FILLER_14_2812 ();
 sg13g2_decap_8 FILLER_14_2822 ();
 sg13g2_fill_2 FILLER_14_2829 ();
 sg13g2_fill_1 FILLER_14_2831 ();
 sg13g2_fill_1 FILLER_14_2837 ();
 sg13g2_decap_4 FILLER_14_2864 ();
 sg13g2_fill_1 FILLER_14_2868 ();
 sg13g2_decap_8 FILLER_14_2903 ();
 sg13g2_fill_1 FILLER_14_2910 ();
 sg13g2_decap_8 FILLER_14_2916 ();
 sg13g2_fill_1 FILLER_14_2932 ();
 sg13g2_fill_1 FILLER_14_2942 ();
 sg13g2_decap_4 FILLER_14_2947 ();
 sg13g2_fill_2 FILLER_14_2951 ();
 sg13g2_decap_8 FILLER_14_2961 ();
 sg13g2_fill_2 FILLER_14_2968 ();
 sg13g2_fill_1 FILLER_14_2970 ();
 sg13g2_decap_4 FILLER_14_2975 ();
 sg13g2_fill_1 FILLER_14_2979 ();
 sg13g2_decap_4 FILLER_14_2993 ();
 sg13g2_fill_1 FILLER_14_2997 ();
 sg13g2_decap_8 FILLER_14_3015 ();
 sg13g2_fill_1 FILLER_14_3036 ();
 sg13g2_fill_2 FILLER_14_3048 ();
 sg13g2_decap_4 FILLER_14_3107 ();
 sg13g2_fill_1 FILLER_14_3111 ();
 sg13g2_decap_8 FILLER_14_3116 ();
 sg13g2_decap_8 FILLER_14_3123 ();
 sg13g2_fill_2 FILLER_14_3130 ();
 sg13g2_fill_1 FILLER_14_3132 ();
 sg13g2_decap_8 FILLER_14_3138 ();
 sg13g2_fill_2 FILLER_14_3155 ();
 sg13g2_fill_2 FILLER_14_3197 ();
 sg13g2_fill_1 FILLER_14_3234 ();
 sg13g2_decap_4 FILLER_14_3270 ();
 sg13g2_fill_1 FILLER_14_3274 ();
 sg13g2_decap_8 FILLER_14_3309 ();
 sg13g2_decap_4 FILLER_14_3316 ();
 sg13g2_fill_1 FILLER_14_3364 ();
 sg13g2_decap_8 FILLER_14_3387 ();
 sg13g2_fill_2 FILLER_14_3394 ();
 sg13g2_decap_4 FILLER_14_3417 ();
 sg13g2_fill_1 FILLER_14_3421 ();
 sg13g2_decap_4 FILLER_14_3444 ();
 sg13g2_fill_2 FILLER_14_3448 ();
 sg13g2_fill_1 FILLER_14_3454 ();
 sg13g2_decap_4 FILLER_14_3459 ();
 sg13g2_fill_1 FILLER_14_3463 ();
 sg13g2_decap_8 FILLER_14_3477 ();
 sg13g2_decap_4 FILLER_14_3484 ();
 sg13g2_fill_2 FILLER_14_3488 ();
 sg13g2_decap_8 FILLER_14_3498 ();
 sg13g2_fill_2 FILLER_14_3505 ();
 sg13g2_fill_1 FILLER_14_3507 ();
 sg13g2_fill_2 FILLER_14_3513 ();
 sg13g2_fill_1 FILLER_14_3515 ();
 sg13g2_fill_2 FILLER_14_3520 ();
 sg13g2_fill_1 FILLER_14_3522 ();
 sg13g2_decap_8 FILLER_14_3527 ();
 sg13g2_fill_2 FILLER_14_3534 ();
 sg13g2_fill_1 FILLER_14_3536 ();
 sg13g2_decap_4 FILLER_14_3550 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_fill_2 FILLER_15_56 ();
 sg13g2_decap_4 FILLER_15_85 ();
 sg13g2_fill_2 FILLER_15_118 ();
 sg13g2_fill_1 FILLER_15_120 ();
 sg13g2_fill_1 FILLER_15_129 ();
 sg13g2_decap_4 FILLER_15_134 ();
 sg13g2_fill_2 FILLER_15_138 ();
 sg13g2_decap_8 FILLER_15_145 ();
 sg13g2_decap_8 FILLER_15_152 ();
 sg13g2_fill_1 FILLER_15_159 ();
 sg13g2_fill_2 FILLER_15_187 ();
 sg13g2_fill_1 FILLER_15_203 ();
 sg13g2_fill_2 FILLER_15_226 ();
 sg13g2_fill_1 FILLER_15_228 ();
 sg13g2_decap_8 FILLER_15_248 ();
 sg13g2_fill_1 FILLER_15_255 ();
 sg13g2_fill_2 FILLER_15_265 ();
 sg13g2_fill_2 FILLER_15_291 ();
 sg13g2_fill_2 FILLER_15_307 ();
 sg13g2_fill_1 FILLER_15_324 ();
 sg13g2_decap_4 FILLER_15_416 ();
 sg13g2_decap_8 FILLER_15_446 ();
 sg13g2_fill_2 FILLER_15_453 ();
 sg13g2_decap_8 FILLER_15_465 ();
 sg13g2_fill_1 FILLER_15_472 ();
 sg13g2_fill_2 FILLER_15_478 ();
 sg13g2_fill_1 FILLER_15_484 ();
 sg13g2_fill_2 FILLER_15_498 ();
 sg13g2_decap_4 FILLER_15_513 ();
 sg13g2_fill_2 FILLER_15_517 ();
 sg13g2_decap_4 FILLER_15_588 ();
 sg13g2_decap_4 FILLER_15_612 ();
 sg13g2_fill_1 FILLER_15_616 ();
 sg13g2_fill_2 FILLER_15_625 ();
 sg13g2_fill_1 FILLER_15_627 ();
 sg13g2_fill_1 FILLER_15_637 ();
 sg13g2_decap_8 FILLER_15_642 ();
 sg13g2_decap_4 FILLER_15_649 ();
 sg13g2_fill_2 FILLER_15_671 ();
 sg13g2_decap_4 FILLER_15_725 ();
 sg13g2_fill_2 FILLER_15_734 ();
 sg13g2_fill_1 FILLER_15_736 ();
 sg13g2_fill_1 FILLER_15_742 ();
 sg13g2_fill_2 FILLER_15_803 ();
 sg13g2_fill_1 FILLER_15_805 ();
 sg13g2_fill_1 FILLER_15_810 ();
 sg13g2_fill_1 FILLER_15_815 ();
 sg13g2_fill_2 FILLER_15_826 ();
 sg13g2_fill_1 FILLER_15_828 ();
 sg13g2_decap_4 FILLER_15_850 ();
 sg13g2_fill_1 FILLER_15_854 ();
 sg13g2_decap_4 FILLER_15_890 ();
 sg13g2_fill_2 FILLER_15_920 ();
 sg13g2_fill_2 FILLER_15_930 ();
 sg13g2_fill_1 FILLER_15_932 ();
 sg13g2_decap_8 FILLER_15_956 ();
 sg13g2_fill_2 FILLER_15_963 ();
 sg13g2_fill_2 FILLER_15_1017 ();
 sg13g2_fill_1 FILLER_15_1019 ();
 sg13g2_fill_1 FILLER_15_1071 ();
 sg13g2_decap_4 FILLER_15_1078 ();
 sg13g2_fill_2 FILLER_15_1091 ();
 sg13g2_fill_1 FILLER_15_1099 ();
 sg13g2_decap_4 FILLER_15_1105 ();
 sg13g2_fill_1 FILLER_15_1109 ();
 sg13g2_decap_8 FILLER_15_1114 ();
 sg13g2_fill_2 FILLER_15_1121 ();
 sg13g2_decap_8 FILLER_15_1141 ();
 sg13g2_fill_2 FILLER_15_1148 ();
 sg13g2_decap_4 FILLER_15_1155 ();
 sg13g2_fill_1 FILLER_15_1159 ();
 sg13g2_fill_2 FILLER_15_1186 ();
 sg13g2_fill_1 FILLER_15_1188 ();
 sg13g2_fill_1 FILLER_15_1207 ();
 sg13g2_fill_1 FILLER_15_1223 ();
 sg13g2_decap_4 FILLER_15_1229 ();
 sg13g2_fill_1 FILLER_15_1233 ();
 sg13g2_fill_1 FILLER_15_1245 ();
 sg13g2_fill_2 FILLER_15_1264 ();
 sg13g2_fill_1 FILLER_15_1274 ();
 sg13g2_decap_8 FILLER_15_1279 ();
 sg13g2_fill_2 FILLER_15_1286 ();
 sg13g2_fill_1 FILLER_15_1288 ();
 sg13g2_fill_2 FILLER_15_1298 ();
 sg13g2_fill_1 FILLER_15_1335 ();
 sg13g2_decap_8 FILLER_15_1340 ();
 sg13g2_decap_8 FILLER_15_1347 ();
 sg13g2_decap_8 FILLER_15_1354 ();
 sg13g2_fill_1 FILLER_15_1386 ();
 sg13g2_fill_2 FILLER_15_1395 ();
 sg13g2_fill_1 FILLER_15_1397 ();
 sg13g2_decap_4 FILLER_15_1432 ();
 sg13g2_fill_2 FILLER_15_1436 ();
 sg13g2_fill_2 FILLER_15_1443 ();
 sg13g2_fill_2 FILLER_15_1450 ();
 sg13g2_decap_4 FILLER_15_1456 ();
 sg13g2_fill_1 FILLER_15_1460 ();
 sg13g2_decap_4 FILLER_15_1466 ();
 sg13g2_fill_1 FILLER_15_1470 ();
 sg13g2_decap_8 FILLER_15_1475 ();
 sg13g2_fill_2 FILLER_15_1482 ();
 sg13g2_fill_1 FILLER_15_1484 ();
 sg13g2_fill_2 FILLER_15_1493 ();
 sg13g2_fill_2 FILLER_15_1503 ();
 sg13g2_fill_1 FILLER_15_1505 ();
 sg13g2_decap_8 FILLER_15_1537 ();
 sg13g2_decap_4 FILLER_15_1544 ();
 sg13g2_fill_1 FILLER_15_1548 ();
 sg13g2_fill_2 FILLER_15_1553 ();
 sg13g2_fill_1 FILLER_15_1555 ();
 sg13g2_decap_8 FILLER_15_1561 ();
 sg13g2_decap_4 FILLER_15_1568 ();
 sg13g2_fill_1 FILLER_15_1572 ();
 sg13g2_fill_2 FILLER_15_1582 ();
 sg13g2_fill_1 FILLER_15_1584 ();
 sg13g2_fill_2 FILLER_15_1599 ();
 sg13g2_fill_1 FILLER_15_1601 ();
 sg13g2_decap_8 FILLER_15_1612 ();
 sg13g2_decap_4 FILLER_15_1619 ();
 sg13g2_fill_2 FILLER_15_1640 ();
 sg13g2_fill_1 FILLER_15_1646 ();
 sg13g2_fill_2 FILLER_15_1656 ();
 sg13g2_decap_4 FILLER_15_1663 ();
 sg13g2_decap_8 FILLER_15_1677 ();
 sg13g2_decap_8 FILLER_15_1684 ();
 sg13g2_decap_4 FILLER_15_1691 ();
 sg13g2_fill_2 FILLER_15_1695 ();
 sg13g2_decap_8 FILLER_15_1726 ();
 sg13g2_fill_1 FILLER_15_1733 ();
 sg13g2_fill_2 FILLER_15_1739 ();
 sg13g2_fill_1 FILLER_15_1749 ();
 sg13g2_decap_4 FILLER_15_1785 ();
 sg13g2_fill_2 FILLER_15_1789 ();
 sg13g2_fill_2 FILLER_15_1806 ();
 sg13g2_fill_1 FILLER_15_1808 ();
 sg13g2_fill_1 FILLER_15_1844 ();
 sg13g2_decap_8 FILLER_15_1849 ();
 sg13g2_fill_2 FILLER_15_1856 ();
 sg13g2_fill_2 FILLER_15_1876 ();
 sg13g2_fill_1 FILLER_15_1878 ();
 sg13g2_fill_2 FILLER_15_1883 ();
 sg13g2_decap_4 FILLER_15_1908 ();
 sg13g2_decap_8 FILLER_15_1917 ();
 sg13g2_fill_2 FILLER_15_1924 ();
 sg13g2_decap_4 FILLER_15_1933 ();
 sg13g2_fill_1 FILLER_15_1937 ();
 sg13g2_fill_2 FILLER_15_1945 ();
 sg13g2_fill_2 FILLER_15_1978 ();
 sg13g2_fill_1 FILLER_15_1980 ();
 sg13g2_fill_2 FILLER_15_2029 ();
 sg13g2_decap_4 FILLER_15_2039 ();
 sg13g2_decap_4 FILLER_15_2047 ();
 sg13g2_fill_2 FILLER_15_2051 ();
 sg13g2_decap_4 FILLER_15_2063 ();
 sg13g2_fill_2 FILLER_15_2075 ();
 sg13g2_fill_1 FILLER_15_2077 ();
 sg13g2_decap_4 FILLER_15_2099 ();
 sg13g2_decap_8 FILLER_15_2169 ();
 sg13g2_fill_1 FILLER_15_2176 ();
 sg13g2_fill_1 FILLER_15_2181 ();
 sg13g2_decap_4 FILLER_15_2223 ();
 sg13g2_decap_4 FILLER_15_2245 ();
 sg13g2_fill_2 FILLER_15_2249 ();
 sg13g2_decap_8 FILLER_15_2277 ();
 sg13g2_fill_1 FILLER_15_2284 ();
 sg13g2_fill_2 FILLER_15_2311 ();
 sg13g2_fill_1 FILLER_15_2313 ();
 sg13g2_fill_1 FILLER_15_2325 ();
 sg13g2_decap_8 FILLER_15_2330 ();
 sg13g2_fill_1 FILLER_15_2337 ();
 sg13g2_fill_2 FILLER_15_2396 ();
 sg13g2_fill_2 FILLER_15_2412 ();
 sg13g2_fill_1 FILLER_15_2414 ();
 sg13g2_decap_8 FILLER_15_2419 ();
 sg13g2_fill_1 FILLER_15_2426 ();
 sg13g2_fill_2 FILLER_15_2462 ();
 sg13g2_fill_1 FILLER_15_2464 ();
 sg13g2_decap_4 FILLER_15_2473 ();
 sg13g2_fill_2 FILLER_15_2529 ();
 sg13g2_fill_1 FILLER_15_2531 ();
 sg13g2_decap_8 FILLER_15_2548 ();
 sg13g2_fill_2 FILLER_15_2555 ();
 sg13g2_fill_1 FILLER_15_2557 ();
 sg13g2_fill_2 FILLER_15_2574 ();
 sg13g2_fill_1 FILLER_15_2576 ();
 sg13g2_fill_2 FILLER_15_2591 ();
 sg13g2_fill_2 FILLER_15_2630 ();
 sg13g2_fill_1 FILLER_15_2632 ();
 sg13g2_decap_4 FILLER_15_2641 ();
 sg13g2_fill_2 FILLER_15_2645 ();
 sg13g2_decap_8 FILLER_15_2665 ();
 sg13g2_decap_8 FILLER_15_2672 ();
 sg13g2_fill_2 FILLER_15_2679 ();
 sg13g2_decap_8 FILLER_15_2685 ();
 sg13g2_decap_8 FILLER_15_2692 ();
 sg13g2_decap_8 FILLER_15_2699 ();
 sg13g2_fill_1 FILLER_15_2706 ();
 sg13g2_fill_2 FILLER_15_2711 ();
 sg13g2_fill_1 FILLER_15_2713 ();
 sg13g2_fill_1 FILLER_15_2719 ();
 sg13g2_decap_8 FILLER_15_2734 ();
 sg13g2_fill_2 FILLER_15_2741 ();
 sg13g2_fill_1 FILLER_15_2743 ();
 sg13g2_fill_1 FILLER_15_2748 ();
 sg13g2_fill_1 FILLER_15_2792 ();
 sg13g2_fill_2 FILLER_15_2847 ();
 sg13g2_decap_4 FILLER_15_2876 ();
 sg13g2_fill_2 FILLER_15_2880 ();
 sg13g2_decap_8 FILLER_15_2896 ();
 sg13g2_fill_1 FILLER_15_2903 ();
 sg13g2_fill_1 FILLER_15_2913 ();
 sg13g2_fill_2 FILLER_15_2919 ();
 sg13g2_fill_2 FILLER_15_2952 ();
 sg13g2_fill_2 FILLER_15_2962 ();
 sg13g2_fill_1 FILLER_15_2964 ();
 sg13g2_decap_8 FILLER_15_2996 ();
 sg13g2_fill_1 FILLER_15_3003 ();
 sg13g2_decap_4 FILLER_15_3012 ();
 sg13g2_decap_8 FILLER_15_3056 ();
 sg13g2_fill_2 FILLER_15_3063 ();
 sg13g2_fill_1 FILLER_15_3065 ();
 sg13g2_decap_8 FILLER_15_3070 ();
 sg13g2_decap_4 FILLER_15_3086 ();
 sg13g2_fill_1 FILLER_15_3094 ();
 sg13g2_fill_2 FILLER_15_3117 ();
 sg13g2_fill_1 FILLER_15_3119 ();
 sg13g2_decap_8 FILLER_15_3158 ();
 sg13g2_decap_8 FILLER_15_3165 ();
 sg13g2_fill_1 FILLER_15_3172 ();
 sg13g2_fill_1 FILLER_15_3177 ();
 sg13g2_fill_2 FILLER_15_3209 ();
 sg13g2_decap_8 FILLER_15_3251 ();
 sg13g2_fill_1 FILLER_15_3258 ();
 sg13g2_decap_8 FILLER_15_3269 ();
 sg13g2_decap_8 FILLER_15_3276 ();
 sg13g2_decap_4 FILLER_15_3287 ();
 sg13g2_fill_2 FILLER_15_3291 ();
 sg13g2_decap_8 FILLER_15_3306 ();
 sg13g2_fill_2 FILLER_15_3313 ();
 sg13g2_fill_2 FILLER_15_3331 ();
 sg13g2_decap_4 FILLER_15_3338 ();
 sg13g2_decap_8 FILLER_15_3346 ();
 sg13g2_decap_4 FILLER_15_3353 ();
 sg13g2_decap_8 FILLER_15_3388 ();
 sg13g2_decap_4 FILLER_15_3395 ();
 sg13g2_fill_2 FILLER_15_3413 ();
 sg13g2_fill_1 FILLER_15_3419 ();
 sg13g2_decap_4 FILLER_15_3451 ();
 sg13g2_fill_2 FILLER_15_3460 ();
 sg13g2_decap_8 FILLER_15_3466 ();
 sg13g2_fill_2 FILLER_15_3473 ();
 sg13g2_decap_8 FILLER_15_3494 ();
 sg13g2_fill_2 FILLER_15_3501 ();
 sg13g2_fill_2 FILLER_15_3521 ();
 sg13g2_fill_2 FILLER_15_3527 ();
 sg13g2_fill_1 FILLER_15_3529 ();
 sg13g2_decap_8 FILLER_15_3560 ();
 sg13g2_fill_2 FILLER_15_3567 ();
 sg13g2_fill_2 FILLER_15_3578 ();
 sg13g2_decap_4 FILLER_16_0 ();
 sg13g2_decap_4 FILLER_16_73 ();
 sg13g2_fill_2 FILLER_16_77 ();
 sg13g2_fill_2 FILLER_16_186 ();
 sg13g2_fill_1 FILLER_16_188 ();
 sg13g2_fill_2 FILLER_16_215 ();
 sg13g2_fill_2 FILLER_16_234 ();
 sg13g2_fill_1 FILLER_16_236 ();
 sg13g2_decap_4 FILLER_16_252 ();
 sg13g2_fill_1 FILLER_16_256 ();
 sg13g2_fill_1 FILLER_16_270 ();
 sg13g2_decap_8 FILLER_16_306 ();
 sg13g2_fill_1 FILLER_16_313 ();
 sg13g2_fill_2 FILLER_16_350 ();
 sg13g2_decap_4 FILLER_16_370 ();
 sg13g2_fill_2 FILLER_16_374 ();
 sg13g2_decap_8 FILLER_16_380 ();
 sg13g2_decap_4 FILLER_16_387 ();
 sg13g2_fill_1 FILLER_16_391 ();
 sg13g2_fill_1 FILLER_16_396 ();
 sg13g2_fill_1 FILLER_16_406 ();
 sg13g2_decap_8 FILLER_16_415 ();
 sg13g2_decap_4 FILLER_16_422 ();
 sg13g2_fill_2 FILLER_16_426 ();
 sg13g2_fill_1 FILLER_16_441 ();
 sg13g2_fill_2 FILLER_16_467 ();
 sg13g2_fill_1 FILLER_16_469 ();
 sg13g2_fill_2 FILLER_16_496 ();
 sg13g2_fill_1 FILLER_16_519 ();
 sg13g2_fill_1 FILLER_16_552 ();
 sg13g2_fill_1 FILLER_16_558 ();
 sg13g2_decap_4 FILLER_16_568 ();
 sg13g2_fill_1 FILLER_16_572 ();
 sg13g2_decap_4 FILLER_16_586 ();
 sg13g2_fill_1 FILLER_16_621 ();
 sg13g2_fill_2 FILLER_16_653 ();
 sg13g2_fill_1 FILLER_16_655 ();
 sg13g2_decap_8 FILLER_16_661 ();
 sg13g2_fill_1 FILLER_16_668 ();
 sg13g2_fill_2 FILLER_16_696 ();
 sg13g2_fill_2 FILLER_16_703 ();
 sg13g2_fill_1 FILLER_16_705 ();
 sg13g2_fill_1 FILLER_16_719 ();
 sg13g2_fill_1 FILLER_16_741 ();
 sg13g2_decap_4 FILLER_16_746 ();
 sg13g2_fill_2 FILLER_16_772 ();
 sg13g2_fill_1 FILLER_16_774 ();
 sg13g2_fill_1 FILLER_16_791 ();
 sg13g2_fill_1 FILLER_16_802 ();
 sg13g2_fill_2 FILLER_16_813 ();
 sg13g2_fill_1 FILLER_16_815 ();
 sg13g2_decap_8 FILLER_16_824 ();
 sg13g2_decap_8 FILLER_16_845 ();
 sg13g2_decap_8 FILLER_16_852 ();
 sg13g2_decap_4 FILLER_16_898 ();
 sg13g2_fill_2 FILLER_16_942 ();
 sg13g2_fill_1 FILLER_16_944 ();
 sg13g2_decap_8 FILLER_16_954 ();
 sg13g2_fill_1 FILLER_16_961 ();
 sg13g2_fill_2 FILLER_16_973 ();
 sg13g2_fill_1 FILLER_16_975 ();
 sg13g2_decap_8 FILLER_16_980 ();
 sg13g2_fill_2 FILLER_16_987 ();
 sg13g2_fill_2 FILLER_16_1020 ();
 sg13g2_fill_1 FILLER_16_1022 ();
 sg13g2_decap_8 FILLER_16_1028 ();
 sg13g2_fill_2 FILLER_16_1035 ();
 sg13g2_decap_4 FILLER_16_1041 ();
 sg13g2_decap_4 FILLER_16_1087 ();
 sg13g2_fill_2 FILLER_16_1125 ();
 sg13g2_fill_1 FILLER_16_1127 ();
 sg13g2_fill_1 FILLER_16_1133 ();
 sg13g2_decap_4 FILLER_16_1142 ();
 sg13g2_fill_1 FILLER_16_1182 ();
 sg13g2_fill_1 FILLER_16_1191 ();
 sg13g2_fill_2 FILLER_16_1233 ();
 sg13g2_fill_1 FILLER_16_1235 ();
 sg13g2_decap_8 FILLER_16_1241 ();
 sg13g2_decap_4 FILLER_16_1266 ();
 sg13g2_decap_4 FILLER_16_1301 ();
 sg13g2_fill_1 FILLER_16_1305 ();
 sg13g2_decap_4 FILLER_16_1310 ();
 sg13g2_fill_2 FILLER_16_1327 ();
 sg13g2_fill_1 FILLER_16_1329 ();
 sg13g2_decap_4 FILLER_16_1338 ();
 sg13g2_fill_1 FILLER_16_1350 ();
 sg13g2_fill_2 FILLER_16_1363 ();
 sg13g2_decap_8 FILLER_16_1391 ();
 sg13g2_fill_2 FILLER_16_1398 ();
 sg13g2_fill_1 FILLER_16_1420 ();
 sg13g2_decap_8 FILLER_16_1425 ();
 sg13g2_fill_2 FILLER_16_1432 ();
 sg13g2_fill_2 FILLER_16_1477 ();
 sg13g2_fill_2 FILLER_16_1519 ();
 sg13g2_fill_2 FILLER_16_1559 ();
 sg13g2_decap_4 FILLER_16_1627 ();
 sg13g2_decap_4 FILLER_16_1683 ();
 sg13g2_fill_2 FILLER_16_1687 ();
 sg13g2_decap_8 FILLER_16_1697 ();
 sg13g2_fill_2 FILLER_16_1704 ();
 sg13g2_fill_1 FILLER_16_1706 ();
 sg13g2_decap_4 FILLER_16_1715 ();
 sg13g2_fill_1 FILLER_16_1719 ();
 sg13g2_decap_8 FILLER_16_1728 ();
 sg13g2_decap_4 FILLER_16_1735 ();
 sg13g2_fill_1 FILLER_16_1739 ();
 sg13g2_fill_1 FILLER_16_1745 ();
 sg13g2_decap_8 FILLER_16_1754 ();
 sg13g2_fill_2 FILLER_16_1761 ();
 sg13g2_fill_1 FILLER_16_1763 ();
 sg13g2_fill_2 FILLER_16_1782 ();
 sg13g2_fill_2 FILLER_16_1814 ();
 sg13g2_fill_1 FILLER_16_1816 ();
 sg13g2_fill_1 FILLER_16_1989 ();
 sg13g2_decap_8 FILLER_16_2006 ();
 sg13g2_fill_2 FILLER_16_2021 ();
 sg13g2_decap_8 FILLER_16_2062 ();
 sg13g2_fill_2 FILLER_16_2069 ();
 sg13g2_fill_1 FILLER_16_2071 ();
 sg13g2_decap_8 FILLER_16_2080 ();
 sg13g2_decap_8 FILLER_16_2087 ();
 sg13g2_decap_4 FILLER_16_2094 ();
 sg13g2_fill_1 FILLER_16_2138 ();
 sg13g2_fill_1 FILLER_16_2152 ();
 sg13g2_fill_2 FILLER_16_2162 ();
 sg13g2_decap_8 FILLER_16_2195 ();
 sg13g2_fill_2 FILLER_16_2253 ();
 sg13g2_fill_2 FILLER_16_2303 ();
 sg13g2_decap_8 FILLER_16_2322 ();
 sg13g2_fill_2 FILLER_16_2334 ();
 sg13g2_decap_4 FILLER_16_2340 ();
 sg13g2_decap_4 FILLER_16_2348 ();
 sg13g2_fill_1 FILLER_16_2352 ();
 sg13g2_fill_1 FILLER_16_2381 ();
 sg13g2_decap_8 FILLER_16_2434 ();
 sg13g2_decap_8 FILLER_16_2441 ();
 sg13g2_fill_2 FILLER_16_2448 ();
 sg13g2_fill_1 FILLER_16_2481 ();
 sg13g2_fill_1 FILLER_16_2503 ();
 sg13g2_fill_2 FILLER_16_2508 ();
 sg13g2_decap_8 FILLER_16_2515 ();
 sg13g2_decap_4 FILLER_16_2522 ();
 sg13g2_fill_1 FILLER_16_2526 ();
 sg13g2_decap_8 FILLER_16_2542 ();
 sg13g2_fill_1 FILLER_16_2549 ();
 sg13g2_fill_2 FILLER_16_2568 ();
 sg13g2_fill_1 FILLER_16_2570 ();
 sg13g2_fill_2 FILLER_16_2597 ();
 sg13g2_fill_1 FILLER_16_2651 ();
 sg13g2_decap_8 FILLER_16_2665 ();
 sg13g2_fill_1 FILLER_16_2672 ();
 sg13g2_fill_1 FILLER_16_2711 ();
 sg13g2_fill_1 FILLER_16_2727 ();
 sg13g2_decap_4 FILLER_16_2769 ();
 sg13g2_fill_2 FILLER_16_2773 ();
 sg13g2_decap_4 FILLER_16_2781 ();
 sg13g2_decap_4 FILLER_16_2807 ();
 sg13g2_fill_1 FILLER_16_2811 ();
 sg13g2_fill_1 FILLER_16_2817 ();
 sg13g2_fill_2 FILLER_16_2826 ();
 sg13g2_decap_4 FILLER_16_2842 ();
 sg13g2_decap_8 FILLER_16_2850 ();
 sg13g2_decap_4 FILLER_16_2913 ();
 sg13g2_decap_8 FILLER_16_2939 ();
 sg13g2_decap_8 FILLER_16_2946 ();
 sg13g2_fill_1 FILLER_16_2953 ();
 sg13g2_fill_2 FILLER_16_2964 ();
 sg13g2_decap_8 FILLER_16_2977 ();
 sg13g2_decap_8 FILLER_16_2984 ();
 sg13g2_fill_1 FILLER_16_2991 ();
 sg13g2_fill_1 FILLER_16_3000 ();
 sg13g2_fill_2 FILLER_16_3006 ();
 sg13g2_decap_4 FILLER_16_3016 ();
 sg13g2_fill_2 FILLER_16_3020 ();
 sg13g2_fill_1 FILLER_16_3039 ();
 sg13g2_fill_1 FILLER_16_3057 ();
 sg13g2_decap_4 FILLER_16_3071 ();
 sg13g2_fill_2 FILLER_16_3080 ();
 sg13g2_decap_8 FILLER_16_3086 ();
 sg13g2_decap_4 FILLER_16_3093 ();
 sg13g2_fill_1 FILLER_16_3097 ();
 sg13g2_decap_4 FILLER_16_3133 ();
 sg13g2_fill_2 FILLER_16_3146 ();
 sg13g2_decap_4 FILLER_16_3152 ();
 sg13g2_fill_1 FILLER_16_3156 ();
 sg13g2_decap_8 FILLER_16_3175 ();
 sg13g2_fill_1 FILLER_16_3191 ();
 sg13g2_fill_1 FILLER_16_3210 ();
 sg13g2_decap_4 FILLER_16_3218 ();
 sg13g2_fill_2 FILLER_16_3222 ();
 sg13g2_fill_1 FILLER_16_3232 ();
 sg13g2_fill_2 FILLER_16_3251 ();
 sg13g2_fill_1 FILLER_16_3253 ();
 sg13g2_decap_8 FILLER_16_3286 ();
 sg13g2_fill_2 FILLER_16_3293 ();
 sg13g2_fill_1 FILLER_16_3295 ();
 sg13g2_fill_2 FILLER_16_3320 ();
 sg13g2_fill_1 FILLER_16_3353 ();
 sg13g2_fill_1 FILLER_16_3359 ();
 sg13g2_fill_2 FILLER_16_3372 ();
 sg13g2_fill_2 FILLER_16_3405 ();
 sg13g2_fill_2 FILLER_16_3411 ();
 sg13g2_decap_8 FILLER_16_3417 ();
 sg13g2_fill_2 FILLER_16_3424 ();
 sg13g2_fill_1 FILLER_16_3426 ();
 sg13g2_decap_8 FILLER_16_3440 ();
 sg13g2_decap_4 FILLER_16_3447 ();
 sg13g2_fill_2 FILLER_16_3477 ();
 sg13g2_decap_4 FILLER_16_3535 ();
 sg13g2_fill_1 FILLER_16_3539 ();
 sg13g2_decap_8 FILLER_16_3553 ();
 sg13g2_decap_4 FILLER_16_3560 ();
 sg13g2_fill_1 FILLER_16_3564 ();
 sg13g2_decap_8 FILLER_16_3569 ();
 sg13g2_decap_4 FILLER_16_3576 ();
 sg13g2_decap_4 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_40 ();
 sg13g2_fill_1 FILLER_17_73 ();
 sg13g2_fill_1 FILLER_17_106 ();
 sg13g2_decap_4 FILLER_17_151 ();
 sg13g2_fill_2 FILLER_17_155 ();
 sg13g2_fill_1 FILLER_17_243 ();
 sg13g2_decap_8 FILLER_17_275 ();
 sg13g2_fill_1 FILLER_17_309 ();
 sg13g2_decap_4 FILLER_17_323 ();
 sg13g2_fill_2 FILLER_17_341 ();
 sg13g2_decap_8 FILLER_17_369 ();
 sg13g2_decap_4 FILLER_17_376 ();
 sg13g2_fill_2 FILLER_17_380 ();
 sg13g2_decap_8 FILLER_17_436 ();
 sg13g2_fill_1 FILLER_17_443 ();
 sg13g2_decap_8 FILLER_17_473 ();
 sg13g2_fill_1 FILLER_17_480 ();
 sg13g2_decap_4 FILLER_17_485 ();
 sg13g2_fill_2 FILLER_17_489 ();
 sg13g2_decap_4 FILLER_17_497 ();
 sg13g2_fill_2 FILLER_17_501 ();
 sg13g2_decap_4 FILLER_17_508 ();
 sg13g2_fill_1 FILLER_17_512 ();
 sg13g2_fill_2 FILLER_17_528 ();
 sg13g2_fill_1 FILLER_17_530 ();
 sg13g2_decap_4 FILLER_17_540 ();
 sg13g2_decap_8 FILLER_17_570 ();
 sg13g2_fill_2 FILLER_17_577 ();
 sg13g2_decap_8 FILLER_17_592 ();
 sg13g2_fill_1 FILLER_17_599 ();
 sg13g2_decap_4 FILLER_17_604 ();
 sg13g2_decap_4 FILLER_17_621 ();
 sg13g2_fill_2 FILLER_17_639 ();
 sg13g2_fill_2 FILLER_17_649 ();
 sg13g2_fill_1 FILLER_17_659 ();
 sg13g2_fill_2 FILLER_17_695 ();
 sg13g2_fill_1 FILLER_17_697 ();
 sg13g2_fill_2 FILLER_17_741 ();
 sg13g2_fill_2 FILLER_17_778 ();
 sg13g2_decap_4 FILLER_17_785 ();
 sg13g2_fill_1 FILLER_17_789 ();
 sg13g2_fill_2 FILLER_17_795 ();
 sg13g2_fill_2 FILLER_17_802 ();
 sg13g2_decap_4 FILLER_17_822 ();
 sg13g2_fill_1 FILLER_17_826 ();
 sg13g2_fill_1 FILLER_17_843 ();
 sg13g2_fill_2 FILLER_17_860 ();
 sg13g2_fill_1 FILLER_17_888 ();
 sg13g2_fill_1 FILLER_17_920 ();
 sg13g2_fill_1 FILLER_17_936 ();
 sg13g2_decap_8 FILLER_17_963 ();
 sg13g2_decap_4 FILLER_17_970 ();
 sg13g2_decap_8 FILLER_17_982 ();
 sg13g2_decap_4 FILLER_17_989 ();
 sg13g2_decap_8 FILLER_17_998 ();
 sg13g2_decap_4 FILLER_17_1009 ();
 sg13g2_fill_2 FILLER_17_1013 ();
 sg13g2_decap_4 FILLER_17_1060 ();
 sg13g2_decap_8 FILLER_17_1078 ();
 sg13g2_decap_8 FILLER_17_1098 ();
 sg13g2_fill_2 FILLER_17_1105 ();
 sg13g2_fill_1 FILLER_17_1107 ();
 sg13g2_decap_4 FILLER_17_1112 ();
 sg13g2_fill_1 FILLER_17_1116 ();
 sg13g2_fill_1 FILLER_17_1131 ();
 sg13g2_decap_4 FILLER_17_1137 ();
 sg13g2_fill_1 FILLER_17_1150 ();
 sg13g2_decap_8 FILLER_17_1155 ();
 sg13g2_decap_4 FILLER_17_1162 ();
 sg13g2_fill_1 FILLER_17_1166 ();
 sg13g2_decap_4 FILLER_17_1175 ();
 sg13g2_fill_1 FILLER_17_1179 ();
 sg13g2_fill_1 FILLER_17_1207 ();
 sg13g2_decap_8 FILLER_17_1221 ();
 sg13g2_decap_4 FILLER_17_1228 ();
 sg13g2_decap_4 FILLER_17_1250 ();
 sg13g2_fill_1 FILLER_17_1259 ();
 sg13g2_fill_1 FILLER_17_1265 ();
 sg13g2_decap_8 FILLER_17_1274 ();
 sg13g2_fill_1 FILLER_17_1281 ();
 sg13g2_decap_4 FILLER_17_1325 ();
 sg13g2_fill_2 FILLER_17_1337 ();
 sg13g2_fill_2 FILLER_17_1365 ();
 sg13g2_fill_1 FILLER_17_1367 ();
 sg13g2_decap_4 FILLER_17_1395 ();
 sg13g2_fill_1 FILLER_17_1399 ();
 sg13g2_decap_8 FILLER_17_1426 ();
 sg13g2_decap_8 FILLER_17_1433 ();
 sg13g2_fill_2 FILLER_17_1457 ();
 sg13g2_fill_1 FILLER_17_1459 ();
 sg13g2_decap_4 FILLER_17_1490 ();
 sg13g2_fill_1 FILLER_17_1494 ();
 sg13g2_fill_2 FILLER_17_1499 ();
 sg13g2_fill_1 FILLER_17_1519 ();
 sg13g2_fill_2 FILLER_17_1549 ();
 sg13g2_decap_8 FILLER_17_1581 ();
 sg13g2_decap_8 FILLER_17_1588 ();
 sg13g2_fill_2 FILLER_17_1595 ();
 sg13g2_fill_1 FILLER_17_1636 ();
 sg13g2_decap_4 FILLER_17_1642 ();
 sg13g2_decap_4 FILLER_17_1654 ();
 sg13g2_decap_8 FILLER_17_1709 ();
 sg13g2_fill_2 FILLER_17_1737 ();
 sg13g2_fill_2 FILLER_17_1782 ();
 sg13g2_fill_1 FILLER_17_1784 ();
 sg13g2_decap_8 FILLER_17_1789 ();
 sg13g2_fill_2 FILLER_17_1812 ();
 sg13g2_fill_1 FILLER_17_1814 ();
 sg13g2_decap_4 FILLER_17_1841 ();
 sg13g2_fill_2 FILLER_17_1845 ();
 sg13g2_decap_4 FILLER_17_1860 ();
 sg13g2_fill_1 FILLER_17_1864 ();
 sg13g2_decap_8 FILLER_17_1874 ();
 sg13g2_decap_8 FILLER_17_1881 ();
 sg13g2_decap_4 FILLER_17_1888 ();
 sg13g2_fill_2 FILLER_17_1892 ();
 sg13g2_decap_4 FILLER_17_1898 ();
 sg13g2_fill_2 FILLER_17_1906 ();
 sg13g2_fill_1 FILLER_17_1908 ();
 sg13g2_decap_4 FILLER_17_1918 ();
 sg13g2_fill_2 FILLER_17_1922 ();
 sg13g2_decap_4 FILLER_17_1963 ();
 sg13g2_decap_8 FILLER_17_1984 ();
 sg13g2_decap_8 FILLER_17_1995 ();
 sg13g2_fill_2 FILLER_17_2002 ();
 sg13g2_fill_2 FILLER_17_2030 ();
 sg13g2_fill_1 FILLER_17_2080 ();
 sg13g2_decap_8 FILLER_17_2094 ();
 sg13g2_decap_8 FILLER_17_2101 ();
 sg13g2_fill_1 FILLER_17_2108 ();
 sg13g2_decap_8 FILLER_17_2113 ();
 sg13g2_fill_2 FILLER_17_2120 ();
 sg13g2_fill_1 FILLER_17_2148 ();
 sg13g2_fill_2 FILLER_17_2175 ();
 sg13g2_fill_2 FILLER_17_2190 ();
 sg13g2_fill_1 FILLER_17_2192 ();
 sg13g2_decap_8 FILLER_17_2197 ();
 sg13g2_fill_2 FILLER_17_2204 ();
 sg13g2_fill_1 FILLER_17_2206 ();
 sg13g2_decap_4 FILLER_17_2218 ();
 sg13g2_fill_2 FILLER_17_2222 ();
 sg13g2_decap_4 FILLER_17_2232 ();
 sg13g2_fill_2 FILLER_17_2236 ();
 sg13g2_decap_8 FILLER_17_2243 ();
 sg13g2_decap_8 FILLER_17_2250 ();
 sg13g2_decap_4 FILLER_17_2257 ();
 sg13g2_fill_1 FILLER_17_2261 ();
 sg13g2_fill_1 FILLER_17_2270 ();
 sg13g2_decap_4 FILLER_17_2280 ();
 sg13g2_decap_4 FILLER_17_2297 ();
 sg13g2_fill_1 FILLER_17_2301 ();
 sg13g2_decap_8 FILLER_17_2318 ();
 sg13g2_fill_2 FILLER_17_2351 ();
 sg13g2_fill_1 FILLER_17_2353 ();
 sg13g2_decap_8 FILLER_17_2385 ();
 sg13g2_decap_4 FILLER_17_2408 ();
 sg13g2_decap_8 FILLER_17_2441 ();
 sg13g2_decap_4 FILLER_17_2448 ();
 sg13g2_decap_4 FILLER_17_2478 ();
 sg13g2_fill_2 FILLER_17_2482 ();
 sg13g2_decap_8 FILLER_17_2519 ();
 sg13g2_fill_2 FILLER_17_2526 ();
 sg13g2_fill_2 FILLER_17_2536 ();
 sg13g2_fill_1 FILLER_17_2538 ();
 sg13g2_fill_2 FILLER_17_2565 ();
 sg13g2_fill_1 FILLER_17_2567 ();
 sg13g2_decap_4 FILLER_17_2573 ();
 sg13g2_decap_4 FILLER_17_2623 ();
 sg13g2_decap_4 FILLER_17_2631 ();
 sg13g2_fill_1 FILLER_17_2639 ();
 sg13g2_fill_1 FILLER_17_2649 ();
 sg13g2_fill_1 FILLER_17_2663 ();
 sg13g2_decap_8 FILLER_17_2668 ();
 sg13g2_decap_8 FILLER_17_2675 ();
 sg13g2_fill_2 FILLER_17_2682 ();
 sg13g2_fill_2 FILLER_17_2688 ();
 sg13g2_fill_1 FILLER_17_2690 ();
 sg13g2_fill_2 FILLER_17_2696 ();
 sg13g2_fill_2 FILLER_17_2707 ();
 sg13g2_decap_8 FILLER_17_2719 ();
 sg13g2_decap_8 FILLER_17_2731 ();
 sg13g2_decap_4 FILLER_17_2738 ();
 sg13g2_fill_2 FILLER_17_2750 ();
 sg13g2_fill_1 FILLER_17_2752 ();
 sg13g2_decap_4 FILLER_17_2757 ();
 sg13g2_fill_1 FILLER_17_2761 ();
 sg13g2_fill_2 FILLER_17_2783 ();
 sg13g2_decap_4 FILLER_17_2801 ();
 sg13g2_fill_2 FILLER_17_2805 ();
 sg13g2_fill_2 FILLER_17_2833 ();
 sg13g2_decap_4 FILLER_17_2865 ();
 sg13g2_fill_2 FILLER_17_2869 ();
 sg13g2_fill_2 FILLER_17_2884 ();
 sg13g2_decap_4 FILLER_17_2897 ();
 sg13g2_fill_2 FILLER_17_2901 ();
 sg13g2_fill_2 FILLER_17_2938 ();
 sg13g2_fill_2 FILLER_17_2964 ();
 sg13g2_fill_1 FILLER_17_2966 ();
 sg13g2_fill_2 FILLER_17_2999 ();
 sg13g2_fill_2 FILLER_17_3027 ();
 sg13g2_fill_1 FILLER_17_3029 ();
 sg13g2_fill_2 FILLER_17_3061 ();
 sg13g2_fill_1 FILLER_17_3063 ();
 sg13g2_decap_8 FILLER_17_3107 ();
 sg13g2_decap_4 FILLER_17_3119 ();
 sg13g2_fill_2 FILLER_17_3163 ();
 sg13g2_fill_1 FILLER_17_3165 ();
 sg13g2_fill_2 FILLER_17_3174 ();
 sg13g2_fill_1 FILLER_17_3176 ();
 sg13g2_decap_4 FILLER_17_3255 ();
 sg13g2_decap_4 FILLER_17_3264 ();
 sg13g2_fill_1 FILLER_17_3268 ();
 sg13g2_fill_1 FILLER_17_3277 ();
 sg13g2_decap_8 FILLER_17_3282 ();
 sg13g2_fill_1 FILLER_17_3319 ();
 sg13g2_fill_1 FILLER_17_3324 ();
 sg13g2_fill_2 FILLER_17_3337 ();
 sg13g2_fill_1 FILLER_17_3339 ();
 sg13g2_fill_2 FILLER_17_3354 ();
 sg13g2_decap_8 FILLER_17_3387 ();
 sg13g2_fill_1 FILLER_17_3394 ();
 sg13g2_fill_1 FILLER_17_3417 ();
 sg13g2_fill_2 FILLER_17_3423 ();
 sg13g2_decap_4 FILLER_17_3456 ();
 sg13g2_fill_1 FILLER_17_3460 ();
 sg13g2_decap_4 FILLER_17_3485 ();
 sg13g2_fill_1 FILLER_17_3489 ();
 sg13g2_decap_8 FILLER_17_3498 ();
 sg13g2_fill_2 FILLER_17_3505 ();
 sg13g2_fill_2 FILLER_17_3516 ();
 sg13g2_decap_8 FILLER_17_3562 ();
 sg13g2_decap_8 FILLER_17_3569 ();
 sg13g2_decap_4 FILLER_17_3576 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_2 ();
 sg13g2_decap_8 FILLER_18_39 ();
 sg13g2_decap_4 FILLER_18_46 ();
 sg13g2_fill_2 FILLER_18_50 ();
 sg13g2_fill_2 FILLER_18_78 ();
 sg13g2_fill_1 FILLER_18_96 ();
 sg13g2_fill_2 FILLER_18_151 ();
 sg13g2_fill_2 FILLER_18_193 ();
 sg13g2_fill_2 FILLER_18_217 ();
 sg13g2_fill_1 FILLER_18_232 ();
 sg13g2_fill_1 FILLER_18_242 ();
 sg13g2_fill_2 FILLER_18_287 ();
 sg13g2_fill_1 FILLER_18_289 ();
 sg13g2_fill_1 FILLER_18_326 ();
 sg13g2_decap_8 FILLER_18_337 ();
 sg13g2_decap_8 FILLER_18_400 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_18_440 ();
 sg13g2_fill_2 FILLER_18_447 ();
 sg13g2_fill_1 FILLER_18_453 ();
 sg13g2_decap_4 FILLER_18_459 ();
 sg13g2_decap_8 FILLER_18_473 ();
 sg13g2_fill_2 FILLER_18_480 ();
 sg13g2_fill_1 FILLER_18_490 ();
 sg13g2_decap_8 FILLER_18_512 ();
 sg13g2_decap_4 FILLER_18_519 ();
 sg13g2_fill_2 FILLER_18_536 ();
 sg13g2_fill_1 FILLER_18_538 ();
 sg13g2_decap_4 FILLER_18_544 ();
 sg13g2_fill_1 FILLER_18_548 ();
 sg13g2_fill_2 FILLER_18_553 ();
 sg13g2_decap_4 FILLER_18_563 ();
 sg13g2_fill_2 FILLER_18_567 ();
 sg13g2_decap_8 FILLER_18_573 ();
 sg13g2_decap_4 FILLER_18_580 ();
 sg13g2_fill_2 FILLER_18_584 ();
 sg13g2_fill_2 FILLER_18_649 ();
 sg13g2_fill_1 FILLER_18_651 ();
 sg13g2_decap_8 FILLER_18_662 ();
 sg13g2_decap_4 FILLER_18_669 ();
 sg13g2_fill_2 FILLER_18_673 ();
 sg13g2_fill_1 FILLER_18_693 ();
 sg13g2_fill_2 FILLER_18_699 ();
 sg13g2_fill_1 FILLER_18_701 ();
 sg13g2_fill_2 FILLER_18_706 ();
 sg13g2_decap_8 FILLER_18_712 ();
 sg13g2_decap_4 FILLER_18_719 ();
 sg13g2_fill_2 FILLER_18_723 ();
 sg13g2_decap_4 FILLER_18_729 ();
 sg13g2_fill_2 FILLER_18_733 ();
 sg13g2_decap_8 FILLER_18_749 ();
 sg13g2_decap_8 FILLER_18_766 ();
 sg13g2_fill_1 FILLER_18_773 ();
 sg13g2_decap_4 FILLER_18_778 ();
 sg13g2_fill_2 FILLER_18_782 ();
 sg13g2_fill_2 FILLER_18_797 ();
 sg13g2_fill_1 FILLER_18_799 ();
 sg13g2_fill_2 FILLER_18_829 ();
 sg13g2_fill_1 FILLER_18_831 ();
 sg13g2_decap_4 FILLER_18_837 ();
 sg13g2_fill_1 FILLER_18_841 ();
 sg13g2_decap_8 FILLER_18_847 ();
 sg13g2_decap_4 FILLER_18_854 ();
 sg13g2_fill_2 FILLER_18_858 ();
 sg13g2_fill_2 FILLER_18_870 ();
 sg13g2_fill_1 FILLER_18_880 ();
 sg13g2_fill_2 FILLER_18_898 ();
 sg13g2_fill_1 FILLER_18_900 ();
 sg13g2_decap_4 FILLER_18_914 ();
 sg13g2_fill_1 FILLER_18_918 ();
 sg13g2_fill_2 FILLER_18_932 ();
 sg13g2_fill_1 FILLER_18_969 ();
 sg13g2_fill_1 FILLER_18_979 ();
 sg13g2_fill_2 FILLER_18_984 ();
 sg13g2_fill_2 FILLER_18_1003 ();
 sg13g2_decap_8 FILLER_18_1031 ();
 sg13g2_fill_2 FILLER_18_1038 ();
 sg13g2_decap_4 FILLER_18_1052 ();
 sg13g2_fill_2 FILLER_18_1056 ();
 sg13g2_fill_1 FILLER_18_1119 ();
 sg13g2_fill_2 FILLER_18_1163 ();
 sg13g2_fill_2 FILLER_18_1196 ();
 sg13g2_fill_1 FILLER_18_1198 ();
 sg13g2_fill_2 FILLER_18_1225 ();
 sg13g2_fill_1 FILLER_18_1227 ();
 sg13g2_fill_1 FILLER_18_1254 ();
 sg13g2_fill_2 FILLER_18_1290 ();
 sg13g2_fill_1 FILLER_18_1292 ();
 sg13g2_fill_1 FILLER_18_1322 ();
 sg13g2_fill_1 FILLER_18_1350 ();
 sg13g2_fill_2 FILLER_18_1360 ();
 sg13g2_fill_1 FILLER_18_1362 ();
 sg13g2_fill_2 FILLER_18_1399 ();
 sg13g2_fill_1 FILLER_18_1401 ();
 sg13g2_fill_2 FILLER_18_1407 ();
 sg13g2_fill_1 FILLER_18_1409 ();
 sg13g2_decap_8 FILLER_18_1414 ();
 sg13g2_decap_8 FILLER_18_1421 ();
 sg13g2_fill_2 FILLER_18_1428 ();
 sg13g2_decap_8 FILLER_18_1456 ();
 sg13g2_fill_2 FILLER_18_1463 ();
 sg13g2_fill_1 FILLER_18_1470 ();
 sg13g2_decap_8 FILLER_18_1475 ();
 sg13g2_decap_4 FILLER_18_1482 ();
 sg13g2_fill_1 FILLER_18_1495 ();
 sg13g2_decap_8 FILLER_18_1522 ();
 sg13g2_decap_8 FILLER_18_1529 ();
 sg13g2_fill_2 FILLER_18_1536 ();
 sg13g2_fill_1 FILLER_18_1538 ();
 sg13g2_fill_2 FILLER_18_1565 ();
 sg13g2_fill_1 FILLER_18_1567 ();
 sg13g2_decap_8 FILLER_18_1612 ();
 sg13g2_decap_8 FILLER_18_1632 ();
 sg13g2_decap_4 FILLER_18_1639 ();
 sg13g2_decap_8 FILLER_18_1647 ();
 sg13g2_fill_2 FILLER_18_1685 ();
 sg13g2_fill_1 FILLER_18_1687 ();
 sg13g2_fill_1 FILLER_18_1709 ();
 sg13g2_decap_8 FILLER_18_1715 ();
 sg13g2_decap_8 FILLER_18_1735 ();
 sg13g2_decap_8 FILLER_18_1742 ();
 sg13g2_decap_4 FILLER_18_1749 ();
 sg13g2_fill_1 FILLER_18_1753 ();
 sg13g2_fill_2 FILLER_18_1762 ();
 sg13g2_fill_2 FILLER_18_1773 ();
 sg13g2_decap_4 FILLER_18_1837 ();
 sg13g2_fill_2 FILLER_18_1849 ();
 sg13g2_decap_4 FILLER_18_1877 ();
 sg13g2_fill_2 FILLER_18_1881 ();
 sg13g2_decap_8 FILLER_18_1908 ();
 sg13g2_fill_1 FILLER_18_1915 ();
 sg13g2_fill_1 FILLER_18_1937 ();
 sg13g2_fill_1 FILLER_18_1956 ();
 sg13g2_decap_4 FILLER_18_1979 ();
 sg13g2_fill_1 FILLER_18_1983 ();
 sg13g2_fill_1 FILLER_18_1988 ();
 sg13g2_decap_8 FILLER_18_2008 ();
 sg13g2_decap_8 FILLER_18_2015 ();
 sg13g2_decap_4 FILLER_18_2030 ();
 sg13g2_fill_1 FILLER_18_2034 ();
 sg13g2_fill_1 FILLER_18_2043 ();
 sg13g2_decap_8 FILLER_18_2056 ();
 sg13g2_decap_4 FILLER_18_2063 ();
 sg13g2_fill_1 FILLER_18_2122 ();
 sg13g2_decap_4 FILLER_18_2128 ();
 sg13g2_fill_1 FILLER_18_2132 ();
 sg13g2_decap_8 FILLER_18_2140 ();
 sg13g2_decap_8 FILLER_18_2147 ();
 sg13g2_decap_4 FILLER_18_2154 ();
 sg13g2_fill_2 FILLER_18_2170 ();
 sg13g2_fill_1 FILLER_18_2172 ();
 sg13g2_fill_1 FILLER_18_2222 ();
 sg13g2_decap_8 FILLER_18_2231 ();
 sg13g2_fill_2 FILLER_18_2238 ();
 sg13g2_fill_2 FILLER_18_2252 ();
 sg13g2_fill_1 FILLER_18_2254 ();
 sg13g2_fill_2 FILLER_18_2284 ();
 sg13g2_decap_4 FILLER_18_2299 ();
 sg13g2_fill_2 FILLER_18_2325 ();
 sg13g2_decap_4 FILLER_18_2339 ();
 sg13g2_fill_1 FILLER_18_2343 ();
 sg13g2_decap_4 FILLER_18_2361 ();
 sg13g2_fill_1 FILLER_18_2369 ();
 sg13g2_decap_4 FILLER_18_2374 ();
 sg13g2_decap_8 FILLER_18_2413 ();
 sg13g2_fill_2 FILLER_18_2447 ();
 sg13g2_fill_1 FILLER_18_2449 ();
 sg13g2_fill_2 FILLER_18_2468 ();
 sg13g2_decap_8 FILLER_18_2479 ();
 sg13g2_decap_4 FILLER_18_2486 ();
 sg13g2_fill_1 FILLER_18_2490 ();
 sg13g2_decap_4 FILLER_18_2509 ();
 sg13g2_fill_2 FILLER_18_2521 ();
 sg13g2_fill_1 FILLER_18_2523 ();
 sg13g2_decap_8 FILLER_18_2532 ();
 sg13g2_decap_4 FILLER_18_2539 ();
 sg13g2_fill_2 FILLER_18_2552 ();
 sg13g2_fill_1 FILLER_18_2558 ();
 sg13g2_fill_2 FILLER_18_2584 ();
 sg13g2_fill_2 FILLER_18_2621 ();
 sg13g2_fill_1 FILLER_18_2623 ();
 sg13g2_decap_4 FILLER_18_2642 ();
 sg13g2_fill_2 FILLER_18_2646 ();
 sg13g2_fill_1 FILLER_18_2679 ();
 sg13g2_decap_8 FILLER_18_2688 ();
 sg13g2_fill_1 FILLER_18_2695 ();
 sg13g2_decap_4 FILLER_18_2700 ();
 sg13g2_fill_1 FILLER_18_2704 ();
 sg13g2_decap_4 FILLER_18_2728 ();
 sg13g2_decap_8 FILLER_18_2758 ();
 sg13g2_decap_8 FILLER_18_2765 ();
 sg13g2_decap_4 FILLER_18_2772 ();
 sg13g2_decap_8 FILLER_18_2802 ();
 sg13g2_fill_1 FILLER_18_2809 ();
 sg13g2_fill_2 FILLER_18_2815 ();
 sg13g2_fill_1 FILLER_18_2817 ();
 sg13g2_decap_4 FILLER_18_2826 ();
 sg13g2_fill_2 FILLER_18_2840 ();
 sg13g2_fill_1 FILLER_18_2871 ();
 sg13g2_decap_8 FILLER_18_2876 ();
 sg13g2_fill_1 FILLER_18_2883 ();
 sg13g2_fill_1 FILLER_18_2888 ();
 sg13g2_decap_8 FILLER_18_2909 ();
 sg13g2_decap_4 FILLER_18_2916 ();
 sg13g2_fill_1 FILLER_18_2920 ();
 sg13g2_decap_8 FILLER_18_2934 ();
 sg13g2_decap_8 FILLER_18_2941 ();
 sg13g2_decap_4 FILLER_18_2948 ();
 sg13g2_fill_2 FILLER_18_2952 ();
 sg13g2_fill_2 FILLER_18_2962 ();
 sg13g2_fill_1 FILLER_18_2964 ();
 sg13g2_decap_4 FILLER_18_2970 ();
 sg13g2_decap_8 FILLER_18_2989 ();
 sg13g2_decap_8 FILLER_18_2996 ();
 sg13g2_fill_1 FILLER_18_3003 ();
 sg13g2_decap_4 FILLER_18_3008 ();
 sg13g2_decap_8 FILLER_18_3025 ();
 sg13g2_decap_4 FILLER_18_3032 ();
 sg13g2_fill_1 FILLER_18_3036 ();
 sg13g2_fill_2 FILLER_18_3044 ();
 sg13g2_decap_8 FILLER_18_3050 ();
 sg13g2_decap_4 FILLER_18_3057 ();
 sg13g2_fill_1 FILLER_18_3061 ();
 sg13g2_decap_8 FILLER_18_3070 ();
 sg13g2_decap_4 FILLER_18_3077 ();
 sg13g2_fill_1 FILLER_18_3081 ();
 sg13g2_decap_4 FILLER_18_3086 ();
 sg13g2_fill_2 FILLER_18_3090 ();
 sg13g2_decap_4 FILLER_18_3095 ();
 sg13g2_fill_2 FILLER_18_3099 ();
 sg13g2_fill_1 FILLER_18_3127 ();
 sg13g2_decap_4 FILLER_18_3149 ();
 sg13g2_decap_8 FILLER_18_3175 ();
 sg13g2_decap_4 FILLER_18_3182 ();
 sg13g2_fill_2 FILLER_18_3186 ();
 sg13g2_decap_4 FILLER_18_3192 ();
 sg13g2_fill_2 FILLER_18_3196 ();
 sg13g2_decap_8 FILLER_18_3211 ();
 sg13g2_decap_8 FILLER_18_3218 ();
 sg13g2_decap_8 FILLER_18_3225 ();
 sg13g2_decap_8 FILLER_18_3232 ();
 sg13g2_fill_1 FILLER_18_3239 ();
 sg13g2_decap_8 FILLER_18_3244 ();
 sg13g2_decap_4 FILLER_18_3251 ();
 sg13g2_fill_2 FILLER_18_3255 ();
 sg13g2_fill_2 FILLER_18_3302 ();
 sg13g2_fill_1 FILLER_18_3304 ();
 sg13g2_fill_2 FILLER_18_3318 ();
 sg13g2_decap_4 FILLER_18_3330 ();
 sg13g2_decap_8 FILLER_18_3389 ();
 sg13g2_fill_2 FILLER_18_3396 ();
 sg13g2_fill_1 FILLER_18_3398 ();
 sg13g2_fill_2 FILLER_18_3402 ();
 sg13g2_decap_8 FILLER_18_3433 ();
 sg13g2_fill_1 FILLER_18_3440 ();
 sg13g2_decap_8 FILLER_18_3445 ();
 sg13g2_decap_8 FILLER_18_3452 ();
 sg13g2_fill_1 FILLER_18_3459 ();
 sg13g2_fill_1 FILLER_18_3472 ();
 sg13g2_fill_2 FILLER_18_3499 ();
 sg13g2_decap_8 FILLER_18_3532 ();
 sg13g2_decap_4 FILLER_18_3539 ();
 sg13g2_fill_1 FILLER_18_3543 ();
 sg13g2_decap_8 FILLER_18_3557 ();
 sg13g2_decap_8 FILLER_18_3564 ();
 sg13g2_decap_8 FILLER_18_3571 ();
 sg13g2_fill_2 FILLER_18_3578 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_28 ();
 sg13g2_fill_1 FILLER_19_30 ();
 sg13g2_fill_2 FILLER_19_57 ();
 sg13g2_fill_1 FILLER_19_96 ();
 sg13g2_fill_2 FILLER_19_155 ();
 sg13g2_fill_1 FILLER_19_174 ();
 sg13g2_fill_2 FILLER_19_189 ();
 sg13g2_fill_1 FILLER_19_191 ();
 sg13g2_fill_1 FILLER_19_234 ();
 sg13g2_fill_2 FILLER_19_244 ();
 sg13g2_fill_2 FILLER_19_263 ();
 sg13g2_decap_8 FILLER_19_275 ();
 sg13g2_fill_2 FILLER_19_299 ();
 sg13g2_decap_4 FILLER_19_315 ();
 sg13g2_fill_1 FILLER_19_319 ();
 sg13g2_fill_1 FILLER_19_346 ();
 sg13g2_fill_1 FILLER_19_365 ();
 sg13g2_fill_2 FILLER_19_383 ();
 sg13g2_decap_4 FILLER_19_389 ();
 sg13g2_fill_2 FILLER_19_393 ();
 sg13g2_fill_1 FILLER_19_400 ();
 sg13g2_fill_2 FILLER_19_409 ();
 sg13g2_fill_2 FILLER_19_420 ();
 sg13g2_fill_2 FILLER_19_426 ();
 sg13g2_fill_2 FILLER_19_481 ();
 sg13g2_fill_1 FILLER_19_483 ();
 sg13g2_decap_8 FILLER_19_504 ();
 sg13g2_decap_8 FILLER_19_511 ();
 sg13g2_fill_2 FILLER_19_518 ();
 sg13g2_fill_1 FILLER_19_520 ();
 sg13g2_decap_4 FILLER_19_526 ();
 sg13g2_fill_1 FILLER_19_530 ();
 sg13g2_fill_2 FILLER_19_536 ();
 sg13g2_fill_1 FILLER_19_538 ();
 sg13g2_fill_2 FILLER_19_590 ();
 sg13g2_decap_8 FILLER_19_601 ();
 sg13g2_decap_8 FILLER_19_608 ();
 sg13g2_fill_1 FILLER_19_615 ();
 sg13g2_decap_4 FILLER_19_620 ();
 sg13g2_fill_1 FILLER_19_624 ();
 sg13g2_decap_8 FILLER_19_633 ();
 sg13g2_decap_8 FILLER_19_640 ();
 sg13g2_fill_1 FILLER_19_647 ();
 sg13g2_fill_2 FILLER_19_656 ();
 sg13g2_fill_1 FILLER_19_658 ();
 sg13g2_fill_1 FILLER_19_664 ();
 sg13g2_fill_2 FILLER_19_705 ();
 sg13g2_fill_1 FILLER_19_707 ();
 sg13g2_fill_1 FILLER_19_712 ();
 sg13g2_decap_4 FILLER_19_727 ();
 sg13g2_fill_1 FILLER_19_731 ();
 sg13g2_fill_1 FILLER_19_758 ();
 sg13g2_decap_8 FILLER_19_800 ();
 sg13g2_decap_4 FILLER_19_807 ();
 sg13g2_fill_1 FILLER_19_811 ();
 sg13g2_fill_2 FILLER_19_818 ();
 sg13g2_decap_8 FILLER_19_828 ();
 sg13g2_fill_1 FILLER_19_835 ();
 sg13g2_fill_2 FILLER_19_852 ();
 sg13g2_fill_2 FILLER_19_859 ();
 sg13g2_fill_1 FILLER_19_861 ();
 sg13g2_decap_4 FILLER_19_914 ();
 sg13g2_fill_2 FILLER_19_918 ();
 sg13g2_fill_2 FILLER_19_925 ();
 sg13g2_fill_2 FILLER_19_958 ();
 sg13g2_fill_2 FILLER_19_968 ();
 sg13g2_fill_2 FILLER_19_1005 ();
 sg13g2_fill_1 FILLER_19_1007 ();
 sg13g2_decap_4 FILLER_19_1031 ();
 sg13g2_decap_8 FILLER_19_1048 ();
 sg13g2_decap_8 FILLER_19_1055 ();
 sg13g2_decap_4 FILLER_19_1062 ();
 sg13g2_fill_1 FILLER_19_1075 ();
 sg13g2_fill_2 FILLER_19_1095 ();
 sg13g2_decap_8 FILLER_19_1136 ();
 sg13g2_decap_4 FILLER_19_1143 ();
 sg13g2_fill_1 FILLER_19_1147 ();
 sg13g2_fill_2 FILLER_19_1152 ();
 sg13g2_decap_8 FILLER_19_1159 ();
 sg13g2_fill_2 FILLER_19_1166 ();
 sg13g2_fill_1 FILLER_19_1168 ();
 sg13g2_decap_8 FILLER_19_1186 ();
 sg13g2_decap_8 FILLER_19_1193 ();
 sg13g2_decap_8 FILLER_19_1200 ();
 sg13g2_fill_2 FILLER_19_1207 ();
 sg13g2_decap_4 FILLER_19_1226 ();
 sg13g2_fill_2 FILLER_19_1235 ();
 sg13g2_fill_2 FILLER_19_1247 ();
 sg13g2_decap_4 FILLER_19_1271 ();
 sg13g2_fill_1 FILLER_19_1297 ();
 sg13g2_fill_1 FILLER_19_1302 ();
 sg13g2_fill_1 FILLER_19_1329 ();
 sg13g2_fill_2 FILLER_19_1335 ();
 sg13g2_fill_1 FILLER_19_1363 ();
 sg13g2_fill_2 FILLER_19_1453 ();
 sg13g2_fill_1 FILLER_19_1455 ();
 sg13g2_decap_4 FILLER_19_1460 ();
 sg13g2_decap_8 FILLER_19_1469 ();
 sg13g2_fill_1 FILLER_19_1476 ();
 sg13g2_decap_4 FILLER_19_1503 ();
 sg13g2_fill_2 FILLER_19_1507 ();
 sg13g2_decap_8 FILLER_19_1535 ();
 sg13g2_fill_1 FILLER_19_1542 ();
 sg13g2_fill_2 FILLER_19_1556 ();
 sg13g2_decap_4 FILLER_19_1563 ();
 sg13g2_fill_1 FILLER_19_1567 ();
 sg13g2_decap_4 FILLER_19_1577 ();
 sg13g2_fill_2 FILLER_19_1581 ();
 sg13g2_fill_2 FILLER_19_1592 ();
 sg13g2_fill_1 FILLER_19_1598 ();
 sg13g2_fill_2 FILLER_19_1665 ();
 sg13g2_fill_1 FILLER_19_1667 ();
 sg13g2_fill_2 FILLER_19_1676 ();
 sg13g2_fill_2 FILLER_19_1682 ();
 sg13g2_decap_4 FILLER_19_1715 ();
 sg13g2_decap_4 FILLER_19_1727 ();
 sg13g2_fill_2 FILLER_19_1731 ();
 sg13g2_fill_1 FILLER_19_1852 ();
 sg13g2_decap_8 FILLER_19_1873 ();
 sg13g2_decap_4 FILLER_19_1880 ();
 sg13g2_fill_1 FILLER_19_1884 ();
 sg13g2_fill_2 FILLER_19_1901 ();
 sg13g2_fill_1 FILLER_19_1903 ();
 sg13g2_decap_8 FILLER_19_1915 ();
 sg13g2_fill_1 FILLER_19_1922 ();
 sg13g2_decap_4 FILLER_19_1937 ();
 sg13g2_fill_1 FILLER_19_1988 ();
 sg13g2_decap_8 FILLER_19_1995 ();
 sg13g2_decap_8 FILLER_19_2002 ();
 sg13g2_fill_2 FILLER_19_2009 ();
 sg13g2_fill_2 FILLER_19_2029 ();
 sg13g2_fill_1 FILLER_19_2039 ();
 sg13g2_decap_8 FILLER_19_2071 ();
 sg13g2_fill_2 FILLER_19_2078 ();
 sg13g2_fill_1 FILLER_19_2080 ();
 sg13g2_fill_2 FILLER_19_2094 ();
 sg13g2_fill_1 FILLER_19_2100 ();
 sg13g2_fill_1 FILLER_19_2138 ();
 sg13g2_fill_1 FILLER_19_2157 ();
 sg13g2_decap_8 FILLER_19_2172 ();
 sg13g2_fill_2 FILLER_19_2187 ();
 sg13g2_fill_1 FILLER_19_2189 ();
 sg13g2_decap_4 FILLER_19_2194 ();
 sg13g2_fill_1 FILLER_19_2198 ();
 sg13g2_fill_2 FILLER_19_2226 ();
 sg13g2_fill_1 FILLER_19_2228 ();
 sg13g2_fill_2 FILLER_19_2282 ();
 sg13g2_decap_8 FILLER_19_2315 ();
 sg13g2_fill_2 FILLER_19_2322 ();
 sg13g2_fill_1 FILLER_19_2324 ();
 sg13g2_decap_8 FILLER_19_2373 ();
 sg13g2_fill_2 FILLER_19_2380 ();
 sg13g2_fill_1 FILLER_19_2382 ();
 sg13g2_decap_4 FILLER_19_2387 ();
 sg13g2_fill_2 FILLER_19_2391 ();
 sg13g2_fill_2 FILLER_19_2401 ();
 sg13g2_fill_1 FILLER_19_2403 ();
 sg13g2_decap_8 FILLER_19_2436 ();
 sg13g2_fill_2 FILLER_19_2443 ();
 sg13g2_fill_1 FILLER_19_2477 ();
 sg13g2_decap_4 FILLER_19_2505 ();
 sg13g2_fill_2 FILLER_19_2513 ();
 sg13g2_fill_2 FILLER_19_2524 ();
 sg13g2_decap_8 FILLER_19_2534 ();
 sg13g2_fill_2 FILLER_19_2541 ();
 sg13g2_decap_8 FILLER_19_2569 ();
 sg13g2_fill_2 FILLER_19_2584 ();
 sg13g2_decap_8 FILLER_19_2594 ();
 sg13g2_decap_8 FILLER_19_2601 ();
 sg13g2_decap_4 FILLER_19_2608 ();
 sg13g2_fill_2 FILLER_19_2620 ();
 sg13g2_fill_2 FILLER_19_2651 ();
 sg13g2_fill_1 FILLER_19_2653 ();
 sg13g2_decap_4 FILLER_19_2658 ();
 sg13g2_decap_4 FILLER_19_2676 ();
 sg13g2_decap_4 FILLER_19_2710 ();
 sg13g2_fill_1 FILLER_19_2714 ();
 sg13g2_fill_2 FILLER_19_2726 ();
 sg13g2_fill_2 FILLER_19_2771 ();
 sg13g2_decap_4 FILLER_19_2782 ();
 sg13g2_fill_1 FILLER_19_2786 ();
 sg13g2_fill_2 FILLER_19_2809 ();
 sg13g2_decap_4 FILLER_19_2831 ();
 sg13g2_fill_2 FILLER_19_2859 ();
 sg13g2_fill_1 FILLER_19_2861 ();
 sg13g2_fill_2 FILLER_19_2888 ();
 sg13g2_decap_8 FILLER_19_2916 ();
 sg13g2_decap_8 FILLER_19_2923 ();
 sg13g2_decap_8 FILLER_19_2943 ();
 sg13g2_fill_2 FILLER_19_2950 ();
 sg13g2_fill_1 FILLER_19_2952 ();
 sg13g2_decap_8 FILLER_19_2966 ();
 sg13g2_fill_2 FILLER_19_2981 ();
 sg13g2_decap_4 FILLER_19_2991 ();
 sg13g2_decap_4 FILLER_19_3026 ();
 sg13g2_decap_4 FILLER_19_3053 ();
 sg13g2_decap_4 FILLER_19_3080 ();
 sg13g2_fill_1 FILLER_19_3084 ();
 sg13g2_decap_4 FILLER_19_3109 ();
 sg13g2_fill_2 FILLER_19_3113 ();
 sg13g2_fill_2 FILLER_19_3124 ();
 sg13g2_fill_2 FILLER_19_3146 ();
 sg13g2_fill_2 FILLER_19_3184 ();
 sg13g2_fill_1 FILLER_19_3186 ();
 sg13g2_fill_2 FILLER_19_3201 ();
 sg13g2_fill_1 FILLER_19_3207 ();
 sg13g2_decap_8 FILLER_19_3222 ();
 sg13g2_fill_1 FILLER_19_3233 ();
 sg13g2_decap_8 FILLER_19_3247 ();
 sg13g2_fill_2 FILLER_19_3254 ();
 sg13g2_fill_2 FILLER_19_3264 ();
 sg13g2_fill_1 FILLER_19_3266 ();
 sg13g2_decap_8 FILLER_19_3276 ();
 sg13g2_fill_1 FILLER_19_3283 ();
 sg13g2_fill_2 FILLER_19_3297 ();
 sg13g2_decap_8 FILLER_19_3318 ();
 sg13g2_fill_1 FILLER_19_3325 ();
 sg13g2_fill_1 FILLER_19_3331 ();
 sg13g2_decap_8 FILLER_19_3337 ();
 sg13g2_decap_8 FILLER_19_3344 ();
 sg13g2_decap_4 FILLER_19_3351 ();
 sg13g2_fill_1 FILLER_19_3355 ();
 sg13g2_decap_4 FILLER_19_3368 ();
 sg13g2_fill_1 FILLER_19_3372 ();
 sg13g2_decap_8 FILLER_19_3403 ();
 sg13g2_decap_8 FILLER_19_3410 ();
 sg13g2_decap_4 FILLER_19_3417 ();
 sg13g2_fill_1 FILLER_19_3444 ();
 sg13g2_decap_8 FILLER_19_3471 ();
 sg13g2_decap_8 FILLER_19_3495 ();
 sg13g2_decap_4 FILLER_19_3502 ();
 sg13g2_fill_2 FILLER_19_3506 ();
 sg13g2_decap_4 FILLER_19_3525 ();
 sg13g2_decap_8 FILLER_19_3564 ();
 sg13g2_decap_8 FILLER_19_3571 ();
 sg13g2_fill_2 FILLER_19_3578 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_7 ();
 sg13g2_fill_1 FILLER_20_9 ();
 sg13g2_fill_2 FILLER_20_37 ();
 sg13g2_fill_2 FILLER_20_90 ();
 sg13g2_decap_8 FILLER_20_118 ();
 sg13g2_decap_8 FILLER_20_125 ();
 sg13g2_fill_2 FILLER_20_132 ();
 sg13g2_fill_1 FILLER_20_134 ();
 sg13g2_fill_1 FILLER_20_139 ();
 sg13g2_fill_1 FILLER_20_148 ();
 sg13g2_fill_2 FILLER_20_185 ();
 sg13g2_fill_1 FILLER_20_187 ();
 sg13g2_decap_4 FILLER_20_263 ();
 sg13g2_fill_1 FILLER_20_267 ();
 sg13g2_decap_4 FILLER_20_324 ();
 sg13g2_fill_1 FILLER_20_328 ();
 sg13g2_fill_1 FILLER_20_347 ();
 sg13g2_decap_4 FILLER_20_384 ();
 sg13g2_fill_2 FILLER_20_388 ();
 sg13g2_decap_4 FILLER_20_416 ();
 sg13g2_fill_2 FILLER_20_463 ();
 sg13g2_fill_1 FILLER_20_474 ();
 sg13g2_fill_1 FILLER_20_484 ();
 sg13g2_fill_1 FILLER_20_493 ();
 sg13g2_decap_4 FILLER_20_525 ();
 sg13g2_fill_1 FILLER_20_555 ();
 sg13g2_decap_8 FILLER_20_560 ();
 sg13g2_decap_4 FILLER_20_567 ();
 sg13g2_fill_2 FILLER_20_571 ();
 sg13g2_fill_1 FILLER_20_583 ();
 sg13g2_fill_2 FILLER_20_590 ();
 sg13g2_fill_1 FILLER_20_592 ();
 sg13g2_fill_1 FILLER_20_629 ();
 sg13g2_decap_8 FILLER_20_650 ();
 sg13g2_fill_2 FILLER_20_657 ();
 sg13g2_decap_8 FILLER_20_664 ();
 sg13g2_decap_4 FILLER_20_671 ();
 sg13g2_fill_1 FILLER_20_675 ();
 sg13g2_decap_8 FILLER_20_680 ();
 sg13g2_decap_8 FILLER_20_687 ();
 sg13g2_fill_2 FILLER_20_694 ();
 sg13g2_fill_1 FILLER_20_696 ();
 sg13g2_decap_8 FILLER_20_733 ();
 sg13g2_fill_1 FILLER_20_740 ();
 sg13g2_fill_2 FILLER_20_750 ();
 sg13g2_fill_2 FILLER_20_761 ();
 sg13g2_fill_1 FILLER_20_763 ();
 sg13g2_decap_4 FILLER_20_770 ();
 sg13g2_decap_8 FILLER_20_778 ();
 sg13g2_fill_1 FILLER_20_785 ();
 sg13g2_decap_8 FILLER_20_802 ();
 sg13g2_fill_2 FILLER_20_809 ();
 sg13g2_fill_1 FILLER_20_811 ();
 sg13g2_fill_2 FILLER_20_820 ();
 sg13g2_decap_8 FILLER_20_838 ();
 sg13g2_decap_8 FILLER_20_853 ();
 sg13g2_decap_8 FILLER_20_860 ();
 sg13g2_decap_4 FILLER_20_867 ();
 sg13g2_fill_2 FILLER_20_871 ();
 sg13g2_decap_8 FILLER_20_877 ();
 sg13g2_decap_8 FILLER_20_884 ();
 sg13g2_fill_2 FILLER_20_891 ();
 sg13g2_decap_8 FILLER_20_906 ();
 sg13g2_decap_8 FILLER_20_927 ();
 sg13g2_fill_1 FILLER_20_934 ();
 sg13g2_fill_2 FILLER_20_940 ();
 sg13g2_fill_1 FILLER_20_942 ();
 sg13g2_fill_1 FILLER_20_947 ();
 sg13g2_decap_8 FILLER_20_956 ();
 sg13g2_decap_4 FILLER_20_963 ();
 sg13g2_fill_1 FILLER_20_967 ();
 sg13g2_fill_2 FILLER_20_972 ();
 sg13g2_fill_1 FILLER_20_974 ();
 sg13g2_decap_8 FILLER_20_979 ();
 sg13g2_decap_4 FILLER_20_986 ();
 sg13g2_fill_2 FILLER_20_990 ();
 sg13g2_fill_1 FILLER_20_1023 ();
 sg13g2_decap_8 FILLER_20_1050 ();
 sg13g2_decap_8 FILLER_20_1057 ();
 sg13g2_fill_2 FILLER_20_1077 ();
 sg13g2_fill_2 FILLER_20_1097 ();
 sg13g2_decap_8 FILLER_20_1134 ();
 sg13g2_decap_4 FILLER_20_1141 ();
 sg13g2_decap_8 FILLER_20_1162 ();
 sg13g2_decap_8 FILLER_20_1169 ();
 sg13g2_decap_8 FILLER_20_1176 ();
 sg13g2_fill_2 FILLER_20_1183 ();
 sg13g2_decap_8 FILLER_20_1196 ();
 sg13g2_fill_1 FILLER_20_1203 ();
 sg13g2_fill_1 FILLER_20_1265 ();
 sg13g2_fill_2 FILLER_20_1297 ();
 sg13g2_fill_2 FILLER_20_1308 ();
 sg13g2_fill_2 FILLER_20_1328 ();
 sg13g2_fill_2 FILLER_20_1356 ();
 sg13g2_fill_1 FILLER_20_1358 ();
 sg13g2_fill_2 FILLER_20_1379 ();
 sg13g2_fill_1 FILLER_20_1381 ();
 sg13g2_fill_1 FILLER_20_1395 ();
 sg13g2_fill_2 FILLER_20_1471 ();
 sg13g2_fill_2 FILLER_20_1486 ();
 sg13g2_fill_2 FILLER_20_1492 ();
 sg13g2_fill_1 FILLER_20_1494 ();
 sg13g2_decap_8 FILLER_20_1500 ();
 sg13g2_fill_1 FILLER_20_1507 ();
 sg13g2_decap_4 FILLER_20_1513 ();
 sg13g2_decap_4 FILLER_20_1527 ();
 sg13g2_decap_4 FILLER_20_1535 ();
 sg13g2_fill_2 FILLER_20_1552 ();
 sg13g2_fill_1 FILLER_20_1554 ();
 sg13g2_fill_2 FILLER_20_1630 ();
 sg13g2_fill_1 FILLER_20_1632 ();
 sg13g2_fill_2 FILLER_20_1641 ();
 sg13g2_decap_4 FILLER_20_1664 ();
 sg13g2_fill_2 FILLER_20_1681 ();
 sg13g2_decap_8 FILLER_20_1692 ();
 sg13g2_fill_1 FILLER_20_1699 ();
 sg13g2_fill_2 FILLER_20_1708 ();
 sg13g2_decap_4 FILLER_20_1719 ();
 sg13g2_decap_4 FILLER_20_1736 ();
 sg13g2_fill_2 FILLER_20_1740 ();
 sg13g2_decap_4 FILLER_20_1747 ();
 sg13g2_fill_1 FILLER_20_1751 ();
 sg13g2_decap_8 FILLER_20_1760 ();
 sg13g2_decap_8 FILLER_20_1767 ();
 sg13g2_fill_2 FILLER_20_1774 ();
 sg13g2_decap_4 FILLER_20_1815 ();
 sg13g2_decap_8 FILLER_20_1823 ();
 sg13g2_fill_2 FILLER_20_1830 ();
 sg13g2_decap_4 FILLER_20_1845 ();
 sg13g2_fill_1 FILLER_20_1849 ();
 sg13g2_decap_4 FILLER_20_1873 ();
 sg13g2_decap_4 FILLER_20_1900 ();
 sg13g2_fill_1 FILLER_20_1919 ();
 sg13g2_decap_4 FILLER_20_1926 ();
 sg13g2_fill_2 FILLER_20_1930 ();
 sg13g2_decap_8 FILLER_20_1937 ();
 sg13g2_decap_8 FILLER_20_1951 ();
 sg13g2_decap_8 FILLER_20_1958 ();
 sg13g2_decap_8 FILLER_20_1965 ();
 sg13g2_fill_1 FILLER_20_1972 ();
 sg13g2_decap_8 FILLER_20_1977 ();
 sg13g2_decap_8 FILLER_20_1984 ();
 sg13g2_decap_4 FILLER_20_1991 ();
 sg13g2_fill_2 FILLER_20_1995 ();
 sg13g2_decap_4 FILLER_20_2020 ();
 sg13g2_fill_1 FILLER_20_2024 ();
 sg13g2_fill_2 FILLER_20_2046 ();
 sg13g2_fill_1 FILLER_20_2048 ();
 sg13g2_decap_8 FILLER_20_2066 ();
 sg13g2_fill_2 FILLER_20_2073 ();
 sg13g2_fill_1 FILLER_20_2075 ();
 sg13g2_fill_1 FILLER_20_2084 ();
 sg13g2_fill_2 FILLER_20_2111 ();
 sg13g2_fill_2 FILLER_20_2119 ();
 sg13g2_fill_1 FILLER_20_2166 ();
 sg13g2_fill_2 FILLER_20_2197 ();
 sg13g2_fill_1 FILLER_20_2199 ();
 sg13g2_decap_8 FILLER_20_2221 ();
 sg13g2_fill_1 FILLER_20_2236 ();
 sg13g2_fill_2 FILLER_20_2259 ();
 sg13g2_fill_2 FILLER_20_2266 ();
 sg13g2_fill_1 FILLER_20_2268 ();
 sg13g2_decap_8 FILLER_20_2274 ();
 sg13g2_decap_8 FILLER_20_2286 ();
 sg13g2_fill_2 FILLER_20_2293 ();
 sg13g2_decap_4 FILLER_20_2315 ();
 sg13g2_fill_2 FILLER_20_2319 ();
 sg13g2_decap_8 FILLER_20_2329 ();
 sg13g2_decap_8 FILLER_20_2336 ();
 sg13g2_fill_2 FILLER_20_2374 ();
 sg13g2_fill_1 FILLER_20_2389 ();
 sg13g2_fill_1 FILLER_20_2394 ();
 sg13g2_decap_4 FILLER_20_2404 ();
 sg13g2_decap_8 FILLER_20_2429 ();
 sg13g2_fill_2 FILLER_20_2436 ();
 sg13g2_fill_1 FILLER_20_2456 ();
 sg13g2_fill_1 FILLER_20_2475 ();
 sg13g2_decap_4 FILLER_20_2567 ();
 sg13g2_fill_2 FILLER_20_2571 ();
 sg13g2_decap_8 FILLER_20_2586 ();
 sg13g2_fill_2 FILLER_20_2593 ();
 sg13g2_fill_2 FILLER_20_2609 ();
 sg13g2_decap_4 FILLER_20_2625 ();
 sg13g2_fill_2 FILLER_20_2629 ();
 sg13g2_decap_8 FILLER_20_2641 ();
 sg13g2_fill_1 FILLER_20_2691 ();
 sg13g2_fill_2 FILLER_20_2701 ();
 sg13g2_fill_1 FILLER_20_2703 ();
 sg13g2_fill_1 FILLER_20_2709 ();
 sg13g2_decap_4 FILLER_20_2730 ();
 sg13g2_decap_8 FILLER_20_2765 ();
 sg13g2_decap_4 FILLER_20_2785 ();
 sg13g2_fill_1 FILLER_20_2789 ();
 sg13g2_decap_8 FILLER_20_2794 ();
 sg13g2_decap_8 FILLER_20_2801 ();
 sg13g2_decap_4 FILLER_20_2814 ();
 sg13g2_decap_8 FILLER_20_2828 ();
 sg13g2_decap_8 FILLER_20_2835 ();
 sg13g2_fill_2 FILLER_20_2842 ();
 sg13g2_fill_1 FILLER_20_2844 ();
 sg13g2_fill_1 FILLER_20_2853 ();
 sg13g2_decap_4 FILLER_20_2868 ();
 sg13g2_fill_1 FILLER_20_2876 ();
 sg13g2_decap_8 FILLER_20_2908 ();
 sg13g2_decap_8 FILLER_20_2915 ();
 sg13g2_decap_4 FILLER_20_2922 ();
 sg13g2_fill_1 FILLER_20_2926 ();
 sg13g2_decap_8 FILLER_20_2953 ();
 sg13g2_decap_4 FILLER_20_2960 ();
 sg13g2_fill_2 FILLER_20_2964 ();
 sg13g2_decap_4 FILLER_20_2971 ();
 sg13g2_decap_8 FILLER_20_3019 ();
 sg13g2_fill_1 FILLER_20_3026 ();
 sg13g2_decap_8 FILLER_20_3050 ();
 sg13g2_fill_2 FILLER_20_3057 ();
 sg13g2_fill_1 FILLER_20_3059 ();
 sg13g2_decap_4 FILLER_20_3100 ();
 sg13g2_fill_1 FILLER_20_3157 ();
 sg13g2_decap_4 FILLER_20_3179 ();
 sg13g2_fill_1 FILLER_20_3183 ();
 sg13g2_decap_4 FILLER_20_3248 ();
 sg13g2_decap_4 FILLER_20_3277 ();
 sg13g2_fill_2 FILLER_20_3301 ();
 sg13g2_fill_2 FILLER_20_3325 ();
 sg13g2_fill_1 FILLER_20_3327 ();
 sg13g2_fill_2 FILLER_20_3337 ();
 sg13g2_fill_1 FILLER_20_3339 ();
 sg13g2_decap_8 FILLER_20_3344 ();
 sg13g2_decap_4 FILLER_20_3351 ();
 sg13g2_fill_1 FILLER_20_3355 ();
 sg13g2_decap_4 FILLER_20_3361 ();
 sg13g2_fill_2 FILLER_20_3391 ();
 sg13g2_fill_2 FILLER_20_3428 ();
 sg13g2_decap_4 FILLER_20_3451 ();
 sg13g2_fill_1 FILLER_20_3455 ();
 sg13g2_decap_8 FILLER_20_3473 ();
 sg13g2_decap_8 FILLER_20_3480 ();
 sg13g2_fill_2 FILLER_20_3487 ();
 sg13g2_fill_1 FILLER_20_3489 ();
 sg13g2_fill_2 FILLER_20_3495 ();
 sg13g2_decap_4 FILLER_20_3523 ();
 sg13g2_fill_1 FILLER_20_3527 ();
 sg13g2_decap_8 FILLER_20_3533 ();
 sg13g2_decap_8 FILLER_20_3540 ();
 sg13g2_decap_8 FILLER_20_3560 ();
 sg13g2_decap_8 FILLER_20_3567 ();
 sg13g2_decap_4 FILLER_20_3574 ();
 sg13g2_fill_2 FILLER_20_3578 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_decap_4 FILLER_21_36 ();
 sg13g2_fill_1 FILLER_21_40 ();
 sg13g2_decap_8 FILLER_21_67 ();
 sg13g2_decap_4 FILLER_21_74 ();
 sg13g2_fill_2 FILLER_21_90 ();
 sg13g2_fill_1 FILLER_21_92 ();
 sg13g2_decap_4 FILLER_21_119 ();
 sg13g2_fill_1 FILLER_21_123 ();
 sg13g2_fill_2 FILLER_21_150 ();
 sg13g2_fill_2 FILLER_21_177 ();
 sg13g2_fill_2 FILLER_21_188 ();
 sg13g2_fill_1 FILLER_21_194 ();
 sg13g2_fill_1 FILLER_21_199 ();
 sg13g2_fill_2 FILLER_21_227 ();
 sg13g2_fill_1 FILLER_21_229 ();
 sg13g2_decap_8 FILLER_21_251 ();
 sg13g2_decap_4 FILLER_21_258 ();
 sg13g2_fill_2 FILLER_21_276 ();
 sg13g2_fill_1 FILLER_21_278 ();
 sg13g2_fill_2 FILLER_21_329 ();
 sg13g2_fill_1 FILLER_21_331 ();
 sg13g2_decap_4 FILLER_21_351 ();
 sg13g2_fill_2 FILLER_21_355 ();
 sg13g2_decap_4 FILLER_21_367 ();
 sg13g2_fill_1 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_398 ();
 sg13g2_fill_1 FILLER_21_405 ();
 sg13g2_decap_8 FILLER_21_411 ();
 sg13g2_fill_2 FILLER_21_418 ();
 sg13g2_fill_1 FILLER_21_420 ();
 sg13g2_fill_2 FILLER_21_425 ();
 sg13g2_decap_8 FILLER_21_436 ();
 sg13g2_fill_1 FILLER_21_443 ();
 sg13g2_fill_2 FILLER_21_492 ();
 sg13g2_decap_4 FILLER_21_506 ();
 sg13g2_fill_2 FILLER_21_528 ();
 sg13g2_decap_8 FILLER_21_538 ();
 sg13g2_decap_4 FILLER_21_545 ();
 sg13g2_decap_4 FILLER_21_554 ();
 sg13g2_decap_4 FILLER_21_583 ();
 sg13g2_fill_2 FILLER_21_587 ();
 sg13g2_decap_8 FILLER_21_599 ();
 sg13g2_decap_8 FILLER_21_606 ();
 sg13g2_decap_8 FILLER_21_613 ();
 sg13g2_decap_4 FILLER_21_620 ();
 sg13g2_fill_2 FILLER_21_624 ();
 sg13g2_decap_4 FILLER_21_652 ();
 sg13g2_fill_1 FILLER_21_656 ();
 sg13g2_decap_4 FILLER_21_671 ();
 sg13g2_fill_1 FILLER_21_675 ();
 sg13g2_fill_2 FILLER_21_681 ();
 sg13g2_fill_1 FILLER_21_683 ();
 sg13g2_decap_4 FILLER_21_692 ();
 sg13g2_decap_4 FILLER_21_717 ();
 sg13g2_decap_4 FILLER_21_725 ();
 sg13g2_fill_2 FILLER_21_729 ();
 sg13g2_fill_2 FILLER_21_737 ();
 sg13g2_fill_1 FILLER_21_739 ();
 sg13g2_decap_8 FILLER_21_749 ();
 sg13g2_fill_2 FILLER_21_805 ();
 sg13g2_fill_2 FILLER_21_835 ();
 sg13g2_fill_1 FILLER_21_837 ();
 sg13g2_fill_2 FILLER_21_854 ();
 sg13g2_decap_8 FILLER_21_880 ();
 sg13g2_fill_2 FILLER_21_887 ();
 sg13g2_fill_2 FILLER_21_914 ();
 sg13g2_fill_1 FILLER_21_924 ();
 sg13g2_fill_2 FILLER_21_938 ();
 sg13g2_fill_2 FILLER_21_1011 ();
 sg13g2_decap_8 FILLER_21_1022 ();
 sg13g2_decap_8 FILLER_21_1029 ();
 sg13g2_fill_2 FILLER_21_1045 ();
 sg13g2_decap_8 FILLER_21_1081 ();
 sg13g2_fill_1 FILLER_21_1088 ();
 sg13g2_fill_2 FILLER_21_1092 ();
 sg13g2_fill_1 FILLER_21_1094 ();
 sg13g2_decap_4 FILLER_21_1129 ();
 sg13g2_fill_1 FILLER_21_1169 ();
 sg13g2_fill_2 FILLER_21_1217 ();
 sg13g2_fill_1 FILLER_21_1229 ();
 sg13g2_fill_1 FILLER_21_1251 ();
 sg13g2_fill_1 FILLER_21_1279 ();
 sg13g2_fill_1 FILLER_21_1284 ();
 sg13g2_fill_2 FILLER_21_1294 ();
 sg13g2_fill_1 FILLER_21_1296 ();
 sg13g2_fill_2 FILLER_21_1336 ();
 sg13g2_decap_4 FILLER_21_1390 ();
 sg13g2_fill_2 FILLER_21_1420 ();
 sg13g2_fill_2 FILLER_21_1442 ();
 sg13g2_fill_1 FILLER_21_1444 ();
 sg13g2_fill_2 FILLER_21_1463 ();
 sg13g2_fill_1 FILLER_21_1465 ();
 sg13g2_decap_8 FILLER_21_1471 ();
 sg13g2_decap_8 FILLER_21_1478 ();
 sg13g2_decap_4 FILLER_21_1485 ();
 sg13g2_fill_1 FILLER_21_1489 ();
 sg13g2_fill_1 FILLER_21_1516 ();
 sg13g2_fill_2 FILLER_21_1546 ();
 sg13g2_fill_2 FILLER_21_1553 ();
 sg13g2_fill_1 FILLER_21_1555 ();
 sg13g2_fill_2 FILLER_21_1561 ();
 sg13g2_fill_2 FILLER_21_1577 ();
 sg13g2_decap_8 FILLER_21_1592 ();
 sg13g2_fill_2 FILLER_21_1599 ();
 sg13g2_fill_1 FILLER_21_1601 ();
 sg13g2_decap_4 FILLER_21_1624 ();
 sg13g2_fill_2 FILLER_21_1628 ();
 sg13g2_decap_4 FILLER_21_1661 ();
 sg13g2_fill_2 FILLER_21_1665 ();
 sg13g2_decap_8 FILLER_21_1693 ();
 sg13g2_fill_1 FILLER_21_1700 ();
 sg13g2_decap_4 FILLER_21_1714 ();
 sg13g2_decap_8 FILLER_21_1731 ();
 sg13g2_fill_2 FILLER_21_1738 ();
 sg13g2_fill_1 FILLER_21_1740 ();
 sg13g2_decap_8 FILLER_21_1776 ();
 sg13g2_fill_2 FILLER_21_1783 ();
 sg13g2_fill_1 FILLER_21_1785 ();
 sg13g2_decap_8 FILLER_21_1790 ();
 sg13g2_decap_4 FILLER_21_1810 ();
 sg13g2_decap_8 FILLER_21_1818 ();
 sg13g2_decap_8 FILLER_21_1825 ();
 sg13g2_fill_2 FILLER_21_1832 ();
 sg13g2_fill_1 FILLER_21_1834 ();
 sg13g2_decap_8 FILLER_21_1861 ();
 sg13g2_decap_4 FILLER_21_1875 ();
 sg13g2_fill_1 FILLER_21_1879 ();
 sg13g2_fill_1 FILLER_21_1885 ();
 sg13g2_decap_8 FILLER_21_1912 ();
 sg13g2_decap_4 FILLER_21_1939 ();
 sg13g2_decap_4 FILLER_21_1949 ();
 sg13g2_decap_4 FILLER_21_1966 ();
 sg13g2_fill_1 FILLER_21_1970 ();
 sg13g2_decap_8 FILLER_21_2001 ();
 sg13g2_decap_8 FILLER_21_2008 ();
 sg13g2_fill_2 FILLER_21_2015 ();
 sg13g2_decap_8 FILLER_21_2025 ();
 sg13g2_decap_8 FILLER_21_2045 ();
 sg13g2_decap_8 FILLER_21_2052 ();
 sg13g2_decap_8 FILLER_21_2072 ();
 sg13g2_decap_4 FILLER_21_2079 ();
 sg13g2_decap_8 FILLER_21_2091 ();
 sg13g2_decap_8 FILLER_21_2098 ();
 sg13g2_decap_4 FILLER_21_2105 ();
 sg13g2_fill_2 FILLER_21_2109 ();
 sg13g2_fill_2 FILLER_21_2128 ();
 sg13g2_decap_4 FILLER_21_2142 ();
 sg13g2_fill_2 FILLER_21_2150 ();
 sg13g2_fill_1 FILLER_21_2152 ();
 sg13g2_fill_2 FILLER_21_2158 ();
 sg13g2_fill_2 FILLER_21_2174 ();
 sg13g2_fill_1 FILLER_21_2176 ();
 sg13g2_fill_2 FILLER_21_2190 ();
 sg13g2_fill_1 FILLER_21_2192 ();
 sg13g2_fill_1 FILLER_21_2207 ();
 sg13g2_fill_1 FILLER_21_2221 ();
 sg13g2_fill_2 FILLER_21_2237 ();
 sg13g2_fill_1 FILLER_21_2239 ();
 sg13g2_fill_2 FILLER_21_2245 ();
 sg13g2_fill_1 FILLER_21_2247 ();
 sg13g2_decap_4 FILLER_21_2272 ();
 sg13g2_fill_2 FILLER_21_2276 ();
 sg13g2_fill_2 FILLER_21_2319 ();
 sg13g2_decap_4 FILLER_21_2353 ();
 sg13g2_fill_2 FILLER_21_2357 ();
 sg13g2_fill_2 FILLER_21_2367 ();
 sg13g2_fill_1 FILLER_21_2378 ();
 sg13g2_decap_8 FILLER_21_2405 ();
 sg13g2_fill_2 FILLER_21_2417 ();
 sg13g2_decap_4 FILLER_21_2424 ();
 sg13g2_fill_1 FILLER_21_2428 ();
 sg13g2_decap_8 FILLER_21_2438 ();
 sg13g2_decap_8 FILLER_21_2445 ();
 sg13g2_decap_4 FILLER_21_2452 ();
 sg13g2_fill_2 FILLER_21_2456 ();
 sg13g2_fill_1 FILLER_21_2472 ();
 sg13g2_decap_8 FILLER_21_2477 ();
 sg13g2_fill_1 FILLER_21_2484 ();
 sg13g2_decap_8 FILLER_21_2502 ();
 sg13g2_decap_8 FILLER_21_2509 ();
 sg13g2_decap_8 FILLER_21_2516 ();
 sg13g2_decap_8 FILLER_21_2523 ();
 sg13g2_decap_8 FILLER_21_2530 ();
 sg13g2_fill_1 FILLER_21_2537 ();
 sg13g2_fill_2 FILLER_21_2546 ();
 sg13g2_decap_8 FILLER_21_2562 ();
 sg13g2_fill_2 FILLER_21_2569 ();
 sg13g2_fill_1 FILLER_21_2571 ();
 sg13g2_fill_1 FILLER_21_2576 ();
 sg13g2_decap_8 FILLER_21_2582 ();
 sg13g2_fill_1 FILLER_21_2589 ();
 sg13g2_fill_2 FILLER_21_2598 ();
 sg13g2_fill_2 FILLER_21_2626 ();
 sg13g2_decap_8 FILLER_21_2654 ();
 sg13g2_fill_2 FILLER_21_2661 ();
 sg13g2_fill_1 FILLER_21_2663 ();
 sg13g2_fill_1 FILLER_21_2668 ();
 sg13g2_decap_8 FILLER_21_2673 ();
 sg13g2_fill_1 FILLER_21_2680 ();
 sg13g2_decap_8 FILLER_21_2706 ();
 sg13g2_decap_4 FILLER_21_2713 ();
 sg13g2_decap_4 FILLER_21_2744 ();
 sg13g2_fill_1 FILLER_21_2748 ();
 sg13g2_decap_8 FILLER_21_2761 ();
 sg13g2_fill_2 FILLER_21_2768 ();
 sg13g2_fill_2 FILLER_21_2805 ();
 sg13g2_fill_1 FILLER_21_2807 ();
 sg13g2_decap_8 FILLER_21_2822 ();
 sg13g2_fill_2 FILLER_21_2833 ();
 sg13g2_fill_1 FILLER_21_2835 ();
 sg13g2_fill_2 FILLER_21_2844 ();
 sg13g2_fill_1 FILLER_21_2846 ();
 sg13g2_fill_1 FILLER_21_2852 ();
 sg13g2_decap_8 FILLER_21_2857 ();
 sg13g2_decap_4 FILLER_21_2925 ();
 sg13g2_fill_2 FILLER_21_2939 ();
 sg13g2_fill_1 FILLER_21_2941 ();
 sg13g2_fill_2 FILLER_21_3004 ();
 sg13g2_fill_1 FILLER_21_3011 ();
 sg13g2_fill_2 FILLER_21_3021 ();
 sg13g2_decap_4 FILLER_21_3035 ();
 sg13g2_fill_1 FILLER_21_3049 ();
 sg13g2_decap_8 FILLER_21_3066 ();
 sg13g2_decap_8 FILLER_21_3073 ();
 sg13g2_fill_1 FILLER_21_3085 ();
 sg13g2_fill_2 FILLER_21_3090 ();
 sg13g2_fill_1 FILLER_21_3106 ();
 sg13g2_fill_1 FILLER_21_3114 ();
 sg13g2_decap_4 FILLER_21_3119 ();
 sg13g2_fill_1 FILLER_21_3123 ();
 sg13g2_decap_8 FILLER_21_3184 ();
 sg13g2_decap_4 FILLER_21_3191 ();
 sg13g2_fill_2 FILLER_21_3195 ();
 sg13g2_fill_2 FILLER_21_3202 ();
 sg13g2_fill_1 FILLER_21_3204 ();
 sg13g2_decap_8 FILLER_21_3209 ();
 sg13g2_fill_2 FILLER_21_3216 ();
 sg13g2_fill_1 FILLER_21_3218 ();
 sg13g2_fill_1 FILLER_21_3223 ();
 sg13g2_decap_8 FILLER_21_3259 ();
 sg13g2_fill_2 FILLER_21_3266 ();
 sg13g2_fill_1 FILLER_21_3276 ();
 sg13g2_decap_4 FILLER_21_3292 ();
 sg13g2_fill_1 FILLER_21_3296 ();
 sg13g2_fill_1 FILLER_21_3328 ();
 sg13g2_fill_2 FILLER_21_3360 ();
 sg13g2_fill_1 FILLER_21_3375 ();
 sg13g2_fill_1 FILLER_21_3380 ();
 sg13g2_decap_8 FILLER_21_3408 ();
 sg13g2_decap_8 FILLER_21_3415 ();
 sg13g2_fill_1 FILLER_21_3422 ();
 sg13g2_fill_2 FILLER_21_3433 ();
 sg13g2_fill_1 FILLER_21_3435 ();
 sg13g2_decap_4 FILLER_21_3441 ();
 sg13g2_fill_1 FILLER_21_3454 ();
 sg13g2_decap_8 FILLER_21_3489 ();
 sg13g2_decap_8 FILLER_21_3496 ();
 sg13g2_fill_2 FILLER_21_3529 ();
 sg13g2_decap_8 FILLER_21_3566 ();
 sg13g2_decap_8 FILLER_21_3573 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_4 FILLER_22_7 ();
 sg13g2_decap_4 FILLER_22_15 ();
 sg13g2_fill_2 FILLER_22_19 ();
 sg13g2_fill_2 FILLER_22_31 ();
 sg13g2_decap_4 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_93 ();
 sg13g2_decap_4 FILLER_22_100 ();
 sg13g2_fill_2 FILLER_22_108 ();
 sg13g2_fill_1 FILLER_22_123 ();
 sg13g2_fill_2 FILLER_22_132 ();
 sg13g2_fill_1 FILLER_22_155 ();
 sg13g2_fill_2 FILLER_22_205 ();
 sg13g2_decap_8 FILLER_22_233 ();
 sg13g2_fill_1 FILLER_22_240 ();
 sg13g2_decap_4 FILLER_22_255 ();
 sg13g2_fill_2 FILLER_22_259 ();
 sg13g2_fill_2 FILLER_22_274 ();
 sg13g2_fill_1 FILLER_22_276 ();
 sg13g2_fill_1 FILLER_22_313 ();
 sg13g2_fill_2 FILLER_22_318 ();
 sg13g2_fill_1 FILLER_22_320 ();
 sg13g2_fill_1 FILLER_22_342 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_decap_4 FILLER_22_406 ();
 sg13g2_decap_8 FILLER_22_445 ();
 sg13g2_fill_1 FILLER_22_452 ();
 sg13g2_decap_8 FILLER_22_462 ();
 sg13g2_decap_4 FILLER_22_469 ();
 sg13g2_fill_1 FILLER_22_473 ();
 sg13g2_fill_2 FILLER_22_509 ();
 sg13g2_fill_2 FILLER_22_516 ();
 sg13g2_fill_1 FILLER_22_518 ();
 sg13g2_decap_4 FILLER_22_580 ();
 sg13g2_fill_1 FILLER_22_584 ();
 sg13g2_fill_1 FILLER_22_698 ();
 sg13g2_decap_8 FILLER_22_750 ();
 sg13g2_decap_4 FILLER_22_757 ();
 sg13g2_fill_1 FILLER_22_761 ();
 sg13g2_fill_2 FILLER_22_777 ();
 sg13g2_fill_1 FILLER_22_779 ();
 sg13g2_decap_4 FILLER_22_806 ();
 sg13g2_decap_8 FILLER_22_831 ();
 sg13g2_fill_2 FILLER_22_838 ();
 sg13g2_fill_1 FILLER_22_840 ();
 sg13g2_fill_2 FILLER_22_867 ();
 sg13g2_decap_4 FILLER_22_905 ();
 sg13g2_fill_2 FILLER_22_909 ();
 sg13g2_fill_2 FILLER_22_955 ();
 sg13g2_fill_1 FILLER_22_957 ();
 sg13g2_decap_4 FILLER_22_976 ();
 sg13g2_fill_1 FILLER_22_980 ();
 sg13g2_fill_2 FILLER_22_1003 ();
 sg13g2_decap_8 FILLER_22_1056 ();
 sg13g2_decap_4 FILLER_22_1063 ();
 sg13g2_decap_4 FILLER_22_1080 ();
 sg13g2_fill_2 FILLER_22_1084 ();
 sg13g2_decap_8 FILLER_22_1119 ();
 sg13g2_fill_2 FILLER_22_1126 ();
 sg13g2_fill_1 FILLER_22_1128 ();
 sg13g2_fill_2 FILLER_22_1198 ();
 sg13g2_fill_2 FILLER_22_1217 ();
 sg13g2_fill_2 FILLER_22_1245 ();
 sg13g2_fill_1 FILLER_22_1247 ();
 sg13g2_fill_2 FILLER_22_1283 ();
 sg13g2_fill_1 FILLER_22_1285 ();
 sg13g2_fill_1 FILLER_22_1315 ();
 sg13g2_fill_1 FILLER_22_1334 ();
 sg13g2_fill_1 FILLER_22_1348 ();
 sg13g2_decap_4 FILLER_22_1373 ();
 sg13g2_fill_2 FILLER_22_1383 ();
 sg13g2_fill_1 FILLER_22_1385 ();
 sg13g2_decap_4 FILLER_22_1392 ();
 sg13g2_decap_4 FILLER_22_1401 ();
 sg13g2_fill_1 FILLER_22_1405 ();
 sg13g2_fill_1 FILLER_22_1432 ();
 sg13g2_fill_2 FILLER_22_1491 ();
 sg13g2_fill_1 FILLER_22_1493 ();
 sg13g2_fill_2 FILLER_22_1502 ();
 sg13g2_decap_8 FILLER_22_1526 ();
 sg13g2_decap_8 FILLER_22_1533 ();
 sg13g2_fill_2 FILLER_22_1597 ();
 sg13g2_fill_1 FILLER_22_1607 ();
 sg13g2_fill_2 FILLER_22_1643 ();
 sg13g2_fill_1 FILLER_22_1645 ();
 sg13g2_fill_2 FILLER_22_1659 ();
 sg13g2_fill_2 FILLER_22_1683 ();
 sg13g2_decap_8 FILLER_22_1698 ();
 sg13g2_decap_8 FILLER_22_1713 ();
 sg13g2_fill_1 FILLER_22_1733 ();
 sg13g2_fill_2 FILLER_22_1747 ();
 sg13g2_fill_2 FILLER_22_1775 ();
 sg13g2_fill_1 FILLER_22_1777 ();
 sg13g2_decap_4 FILLER_22_1786 ();
 sg13g2_decap_8 FILLER_22_1829 ();
 sg13g2_decap_8 FILLER_22_1836 ();
 sg13g2_fill_1 FILLER_22_1843 ();
 sg13g2_fill_1 FILLER_22_1862 ();
 sg13g2_decap_8 FILLER_22_1872 ();
 sg13g2_decap_8 FILLER_22_1879 ();
 sg13g2_fill_2 FILLER_22_1886 ();
 sg13g2_fill_1 FILLER_22_1888 ();
 sg13g2_decap_8 FILLER_22_1915 ();
 sg13g2_fill_1 FILLER_22_1922 ();
 sg13g2_decap_4 FILLER_22_1941 ();
 sg13g2_fill_1 FILLER_22_1966 ();
 sg13g2_fill_2 FILLER_22_1980 ();
 sg13g2_decap_8 FILLER_22_1986 ();
 sg13g2_decap_8 FILLER_22_1993 ();
 sg13g2_fill_2 FILLER_22_2000 ();
 sg13g2_decap_8 FILLER_22_2019 ();
 sg13g2_decap_8 FILLER_22_2026 ();
 sg13g2_decap_8 FILLER_22_2033 ();
 sg13g2_decap_8 FILLER_22_2040 ();
 sg13g2_decap_8 FILLER_22_2047 ();
 sg13g2_fill_2 FILLER_22_2054 ();
 sg13g2_fill_1 FILLER_22_2056 ();
 sg13g2_decap_4 FILLER_22_2073 ();
 sg13g2_fill_1 FILLER_22_2077 ();
 sg13g2_decap_4 FILLER_22_2089 ();
 sg13g2_fill_2 FILLER_22_2101 ();
 sg13g2_fill_1 FILLER_22_2103 ();
 sg13g2_fill_1 FILLER_22_2134 ();
 sg13g2_fill_2 FILLER_22_2204 ();
 sg13g2_decap_8 FILLER_22_2214 ();
 sg13g2_decap_8 FILLER_22_2221 ();
 sg13g2_fill_1 FILLER_22_2228 ();
 sg13g2_decap_8 FILLER_22_2239 ();
 sg13g2_decap_8 FILLER_22_2246 ();
 sg13g2_fill_2 FILLER_22_2253 ();
 sg13g2_fill_1 FILLER_22_2255 ();
 sg13g2_fill_1 FILLER_22_2265 ();
 sg13g2_decap_8 FILLER_22_2271 ();
 sg13g2_fill_2 FILLER_22_2278 ();
 sg13g2_fill_1 FILLER_22_2288 ();
 sg13g2_decap_8 FILLER_22_2320 ();
 sg13g2_decap_4 FILLER_22_2327 ();
 sg13g2_fill_1 FILLER_22_2331 ();
 sg13g2_decap_4 FILLER_22_2356 ();
 sg13g2_fill_2 FILLER_22_2360 ();
 sg13g2_decap_8 FILLER_22_2370 ();
 sg13g2_decap_4 FILLER_22_2377 ();
 sg13g2_fill_1 FILLER_22_2381 ();
 sg13g2_decap_8 FILLER_22_2395 ();
 sg13g2_fill_2 FILLER_22_2402 ();
 sg13g2_fill_1 FILLER_22_2404 ();
 sg13g2_fill_2 FILLER_22_2426 ();
 sg13g2_fill_1 FILLER_22_2434 ();
 sg13g2_decap_4 FILLER_22_2443 ();
 sg13g2_fill_2 FILLER_22_2452 ();
 sg13g2_fill_2 FILLER_22_2472 ();
 sg13g2_fill_1 FILLER_22_2474 ();
 sg13g2_decap_4 FILLER_22_2562 ();
 sg13g2_fill_1 FILLER_22_2566 ();
 sg13g2_decap_4 FILLER_22_2601 ();
 sg13g2_fill_2 FILLER_22_2605 ();
 sg13g2_decap_8 FILLER_22_2616 ();
 sg13g2_decap_8 FILLER_22_2623 ();
 sg13g2_fill_2 FILLER_22_2630 ();
 sg13g2_fill_1 FILLER_22_2649 ();
 sg13g2_fill_2 FILLER_22_2690 ();
 sg13g2_decap_8 FILLER_22_2756 ();
 sg13g2_decap_4 FILLER_22_2763 ();
 sg13g2_fill_2 FILLER_22_2802 ();
 sg13g2_fill_1 FILLER_22_2804 ();
 sg13g2_fill_2 FILLER_22_2844 ();
 sg13g2_fill_2 FILLER_22_2881 ();
 sg13g2_fill_1 FILLER_22_2883 ();
 sg13g2_fill_1 FILLER_22_2898 ();
 sg13g2_decap_4 FILLER_22_2920 ();
 sg13g2_fill_2 FILLER_22_2924 ();
 sg13g2_decap_4 FILLER_22_2942 ();
 sg13g2_fill_1 FILLER_22_2946 ();
 sg13g2_fill_2 FILLER_22_2955 ();
 sg13g2_fill_1 FILLER_22_2957 ();
 sg13g2_fill_2 FILLER_22_2971 ();
 sg13g2_fill_1 FILLER_22_2973 ();
 sg13g2_fill_2 FILLER_22_2979 ();
 sg13g2_decap_4 FILLER_22_3009 ();
 sg13g2_fill_2 FILLER_22_3048 ();
 sg13g2_decap_4 FILLER_22_3058 ();
 sg13g2_fill_1 FILLER_22_3062 ();
 sg13g2_decap_8 FILLER_22_3071 ();
 sg13g2_decap_8 FILLER_22_3112 ();
 sg13g2_decap_4 FILLER_22_3119 ();
 sg13g2_fill_1 FILLER_22_3123 ();
 sg13g2_decap_8 FILLER_22_3133 ();
 sg13g2_decap_8 FILLER_22_3140 ();
 sg13g2_fill_2 FILLER_22_3151 ();
 sg13g2_fill_1 FILLER_22_3153 ();
 sg13g2_fill_2 FILLER_22_3159 ();
 sg13g2_fill_2 FILLER_22_3166 ();
 sg13g2_fill_1 FILLER_22_3168 ();
 sg13g2_decap_8 FILLER_22_3173 ();
 sg13g2_decap_8 FILLER_22_3180 ();
 sg13g2_decap_8 FILLER_22_3187 ();
 sg13g2_fill_2 FILLER_22_3220 ();
 sg13g2_fill_2 FILLER_22_3246 ();
 sg13g2_fill_1 FILLER_22_3248 ();
 sg13g2_fill_2 FILLER_22_3280 ();
 sg13g2_fill_1 FILLER_22_3282 ();
 sg13g2_decap_8 FILLER_22_3287 ();
 sg13g2_decap_8 FILLER_22_3294 ();
 sg13g2_decap_8 FILLER_22_3301 ();
 sg13g2_decap_8 FILLER_22_3312 ();
 sg13g2_decap_8 FILLER_22_3319 ();
 sg13g2_decap_4 FILLER_22_3326 ();
 sg13g2_fill_2 FILLER_22_3357 ();
 sg13g2_fill_1 FILLER_22_3359 ();
 sg13g2_fill_2 FILLER_22_3365 ();
 sg13g2_decap_4 FILLER_22_3393 ();
 sg13g2_decap_4 FILLER_22_3414 ();
 sg13g2_fill_2 FILLER_22_3418 ();
 sg13g2_fill_2 FILLER_22_3425 ();
 sg13g2_fill_1 FILLER_22_3427 ();
 sg13g2_fill_2 FILLER_22_3439 ();
 sg13g2_fill_1 FILLER_22_3515 ();
 sg13g2_decap_4 FILLER_22_3525 ();
 sg13g2_fill_1 FILLER_22_3529 ();
 sg13g2_decap_4 FILLER_22_3534 ();
 sg13g2_fill_2 FILLER_22_3538 ();
 sg13g2_decap_4 FILLER_22_3545 ();
 sg13g2_decap_8 FILLER_22_3562 ();
 sg13g2_decap_8 FILLER_22_3569 ();
 sg13g2_decap_4 FILLER_22_3576 ();
 sg13g2_fill_2 FILLER_23_38 ();
 sg13g2_fill_1 FILLER_23_40 ();
 sg13g2_fill_2 FILLER_23_64 ();
 sg13g2_fill_1 FILLER_23_66 ();
 sg13g2_decap_8 FILLER_23_76 ();
 sg13g2_fill_1 FILLER_23_83 ();
 sg13g2_decap_8 FILLER_23_120 ();
 sg13g2_decap_8 FILLER_23_127 ();
 sg13g2_fill_2 FILLER_23_134 ();
 sg13g2_fill_1 FILLER_23_136 ();
 sg13g2_fill_2 FILLER_23_167 ();
 sg13g2_fill_1 FILLER_23_186 ();
 sg13g2_fill_2 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_208 ();
 sg13g2_fill_1 FILLER_23_215 ();
 sg13g2_decap_8 FILLER_23_229 ();
 sg13g2_decap_8 FILLER_23_236 ();
 sg13g2_decap_8 FILLER_23_247 ();
 sg13g2_fill_2 FILLER_23_254 ();
 sg13g2_fill_1 FILLER_23_286 ();
 sg13g2_fill_2 FILLER_23_323 ();
 sg13g2_decap_4 FILLER_23_366 ();
 sg13g2_decap_8 FILLER_23_401 ();
 sg13g2_decap_4 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_23_442 ();
 sg13g2_fill_2 FILLER_23_449 ();
 sg13g2_fill_1 FILLER_23_451 ();
 sg13g2_decap_8 FILLER_23_478 ();
 sg13g2_fill_2 FILLER_23_485 ();
 sg13g2_fill_2 FILLER_23_505 ();
 sg13g2_fill_1 FILLER_23_507 ();
 sg13g2_decap_4 FILLER_23_534 ();
 sg13g2_fill_1 FILLER_23_564 ();
 sg13g2_fill_1 FILLER_23_569 ();
 sg13g2_fill_1 FILLER_23_579 ();
 sg13g2_fill_2 FILLER_23_585 ();
 sg13g2_fill_1 FILLER_23_592 ();
 sg13g2_decap_8 FILLER_23_622 ();
 sg13g2_fill_1 FILLER_23_685 ();
 sg13g2_fill_2 FILLER_23_730 ();
 sg13g2_fill_1 FILLER_23_746 ();
 sg13g2_decap_4 FILLER_23_755 ();
 sg13g2_fill_1 FILLER_23_759 ();
 sg13g2_fill_2 FILLER_23_770 ();
 sg13g2_decap_4 FILLER_23_776 ();
 sg13g2_fill_1 FILLER_23_780 ();
 sg13g2_decap_8 FILLER_23_807 ();
 sg13g2_fill_2 FILLER_23_814 ();
 sg13g2_fill_1 FILLER_23_816 ();
 sg13g2_decap_8 FILLER_23_823 ();
 sg13g2_decap_4 FILLER_23_830 ();
 sg13g2_fill_2 FILLER_23_834 ();
 sg13g2_fill_2 FILLER_23_840 ();
 sg13g2_decap_4 FILLER_23_851 ();
 sg13g2_fill_2 FILLER_23_877 ();
 sg13g2_fill_1 FILLER_23_879 ();
 sg13g2_decap_8 FILLER_23_910 ();
 sg13g2_decap_4 FILLER_23_917 ();
 sg13g2_fill_1 FILLER_23_921 ();
 sg13g2_decap_8 FILLER_23_944 ();
 sg13g2_fill_2 FILLER_23_955 ();
 sg13g2_decap_4 FILLER_23_983 ();
 sg13g2_fill_2 FILLER_23_1013 ();
 sg13g2_decap_4 FILLER_23_1024 ();
 sg13g2_fill_1 FILLER_23_1033 ();
 sg13g2_fill_2 FILLER_23_1060 ();
 sg13g2_fill_1 FILLER_23_1062 ();
 sg13g2_decap_8 FILLER_23_1089 ();
 sg13g2_decap_4 FILLER_23_1096 ();
 sg13g2_decap_8 FILLER_23_1113 ();
 sg13g2_fill_1 FILLER_23_1146 ();
 sg13g2_fill_1 FILLER_23_1156 ();
 sg13g2_fill_2 FILLER_23_1192 ();
 sg13g2_fill_1 FILLER_23_1232 ();
 sg13g2_fill_2 FILLER_23_1289 ();
 sg13g2_fill_2 FILLER_23_1296 ();
 sg13g2_decap_4 FILLER_23_1358 ();
 sg13g2_fill_1 FILLER_23_1362 ();
 sg13g2_fill_1 FILLER_23_1375 ();
 sg13g2_decap_8 FILLER_23_1393 ();
 sg13g2_decap_8 FILLER_23_1400 ();
 sg13g2_fill_2 FILLER_23_1407 ();
 sg13g2_fill_2 FILLER_23_1414 ();
 sg13g2_fill_1 FILLER_23_1416 ();
 sg13g2_decap_4 FILLER_23_1421 ();
 sg13g2_fill_1 FILLER_23_1429 ();
 sg13g2_fill_2 FILLER_23_1435 ();
 sg13g2_fill_1 FILLER_23_1441 ();
 sg13g2_decap_8 FILLER_23_1484 ();
 sg13g2_decap_4 FILLER_23_1491 ();
 sg13g2_fill_1 FILLER_23_1495 ();
 sg13g2_decap_8 FILLER_23_1533 ();
 sg13g2_decap_4 FILLER_23_1540 ();
 sg13g2_decap_8 FILLER_23_1556 ();
 sg13g2_decap_8 FILLER_23_1563 ();
 sg13g2_fill_1 FILLER_23_1570 ();
 sg13g2_fill_1 FILLER_23_1589 ();
 sg13g2_decap_8 FILLER_23_1598 ();
 sg13g2_decap_8 FILLER_23_1605 ();
 sg13g2_decap_4 FILLER_23_1612 ();
 sg13g2_fill_2 FILLER_23_1616 ();
 sg13g2_decap_8 FILLER_23_1622 ();
 sg13g2_decap_8 FILLER_23_1629 ();
 sg13g2_decap_4 FILLER_23_1636 ();
 sg13g2_decap_8 FILLER_23_1648 ();
 sg13g2_fill_2 FILLER_23_1655 ();
 sg13g2_fill_2 FILLER_23_1661 ();
 sg13g2_fill_1 FILLER_23_1663 ();
 sg13g2_decap_8 FILLER_23_1694 ();
 sg13g2_fill_1 FILLER_23_1701 ();
 sg13g2_decap_4 FILLER_23_1706 ();
 sg13g2_fill_1 FILLER_23_1710 ();
 sg13g2_fill_2 FILLER_23_1744 ();
 sg13g2_decap_8 FILLER_23_1751 ();
 sg13g2_decap_8 FILLER_23_1766 ();
 sg13g2_fill_2 FILLER_23_1773 ();
 sg13g2_decap_8 FILLER_23_1801 ();
 sg13g2_decap_4 FILLER_23_1834 ();
 sg13g2_fill_2 FILLER_23_1838 ();
 sg13g2_decap_8 FILLER_23_1856 ();
 sg13g2_decap_8 FILLER_23_1889 ();
 sg13g2_decap_8 FILLER_23_1896 ();
 sg13g2_decap_4 FILLER_23_1903 ();
 sg13g2_decap_8 FILLER_23_1910 ();
 sg13g2_fill_1 FILLER_23_1917 ();
 sg13g2_decap_8 FILLER_23_1944 ();
 sg13g2_decap_8 FILLER_23_1951 ();
 sg13g2_decap_8 FILLER_23_1958 ();
 sg13g2_fill_2 FILLER_23_1965 ();
 sg13g2_fill_1 FILLER_23_1967 ();
 sg13g2_decap_4 FILLER_23_1981 ();
 sg13g2_fill_1 FILLER_23_1985 ();
 sg13g2_decap_8 FILLER_23_2041 ();
 sg13g2_decap_8 FILLER_23_2048 ();
 sg13g2_decap_8 FILLER_23_2055 ();
 sg13g2_decap_4 FILLER_23_2074 ();
 sg13g2_decap_8 FILLER_23_2086 ();
 sg13g2_fill_1 FILLER_23_2093 ();
 sg13g2_decap_8 FILLER_23_2129 ();
 sg13g2_decap_4 FILLER_23_2136 ();
 sg13g2_decap_4 FILLER_23_2153 ();
 sg13g2_fill_1 FILLER_23_2157 ();
 sg13g2_fill_2 FILLER_23_2162 ();
 sg13g2_fill_2 FILLER_23_2169 ();
 sg13g2_decap_8 FILLER_23_2179 ();
 sg13g2_decap_4 FILLER_23_2186 ();
 sg13g2_fill_2 FILLER_23_2198 ();
 sg13g2_decap_8 FILLER_23_2209 ();
 sg13g2_decap_8 FILLER_23_2216 ();
 sg13g2_fill_1 FILLER_23_2223 ();
 sg13g2_decap_4 FILLER_23_2232 ();
 sg13g2_fill_2 FILLER_23_2236 ();
 sg13g2_decap_4 FILLER_23_2255 ();
 sg13g2_fill_2 FILLER_23_2272 ();
 sg13g2_decap_4 FILLER_23_2283 ();
 sg13g2_fill_1 FILLER_23_2287 ();
 sg13g2_fill_2 FILLER_23_2293 ();
 sg13g2_decap_4 FILLER_23_2299 ();
 sg13g2_fill_2 FILLER_23_2303 ();
 sg13g2_decap_4 FILLER_23_2309 ();
 sg13g2_fill_1 FILLER_23_2313 ();
 sg13g2_decap_8 FILLER_23_2322 ();
 sg13g2_fill_2 FILLER_23_2329 ();
 sg13g2_fill_1 FILLER_23_2331 ();
 sg13g2_decap_8 FILLER_23_2336 ();
 sg13g2_decap_8 FILLER_23_2343 ();
 sg13g2_fill_1 FILLER_23_2350 ();
 sg13g2_decap_4 FILLER_23_2416 ();
 sg13g2_fill_1 FILLER_23_2420 ();
 sg13g2_decap_8 FILLER_23_2431 ();
 sg13g2_decap_8 FILLER_23_2438 ();
 sg13g2_fill_1 FILLER_23_2445 ();
 sg13g2_decap_8 FILLER_23_2465 ();
 sg13g2_fill_2 FILLER_23_2472 ();
 sg13g2_decap_8 FILLER_23_2500 ();
 sg13g2_fill_2 FILLER_23_2507 ();
 sg13g2_fill_1 FILLER_23_2509 ();
 sg13g2_decap_8 FILLER_23_2519 ();
 sg13g2_decap_4 FILLER_23_2526 ();
 sg13g2_fill_1 FILLER_23_2530 ();
 sg13g2_fill_1 FILLER_23_2545 ();
 sg13g2_decap_8 FILLER_23_2550 ();
 sg13g2_decap_8 FILLER_23_2557 ();
 sg13g2_fill_1 FILLER_23_2564 ();
 sg13g2_decap_8 FILLER_23_2570 ();
 sg13g2_fill_2 FILLER_23_2577 ();
 sg13g2_decap_4 FILLER_23_2582 ();
 sg13g2_fill_2 FILLER_23_2591 ();
 sg13g2_fill_1 FILLER_23_2634 ();
 sg13g2_decap_4 FILLER_23_2648 ();
 sg13g2_decap_4 FILLER_23_2656 ();
 sg13g2_fill_2 FILLER_23_2669 ();
 sg13g2_fill_1 FILLER_23_2671 ();
 sg13g2_decap_4 FILLER_23_2693 ();
 sg13g2_fill_2 FILLER_23_2697 ();
 sg13g2_decap_8 FILLER_23_2721 ();
 sg13g2_decap_4 FILLER_23_2728 ();
 sg13g2_fill_1 FILLER_23_2732 ();
 sg13g2_decap_8 FILLER_23_2745 ();
 sg13g2_fill_2 FILLER_23_2752 ();
 sg13g2_fill_1 FILLER_23_2754 ();
 sg13g2_decap_8 FILLER_23_2763 ();
 sg13g2_fill_2 FILLER_23_2770 ();
 sg13g2_fill_1 FILLER_23_2772 ();
 sg13g2_fill_2 FILLER_23_2778 ();
 sg13g2_fill_1 FILLER_23_2780 ();
 sg13g2_fill_1 FILLER_23_2816 ();
 sg13g2_fill_2 FILLER_23_2831 ();
 sg13g2_fill_2 FILLER_23_2850 ();
 sg13g2_fill_1 FILLER_23_2852 ();
 sg13g2_decap_8 FILLER_23_2869 ();
 sg13g2_fill_2 FILLER_23_2876 ();
 sg13g2_fill_1 FILLER_23_2878 ();
 sg13g2_decap_8 FILLER_23_2896 ();
 sg13g2_fill_1 FILLER_23_2903 ();
 sg13g2_fill_2 FILLER_23_2920 ();
 sg13g2_decap_8 FILLER_23_2940 ();
 sg13g2_fill_2 FILLER_23_2947 ();
 sg13g2_fill_1 FILLER_23_2949 ();
 sg13g2_decap_8 FILLER_23_3005 ();
 sg13g2_decap_8 FILLER_23_3012 ();
 sg13g2_decap_4 FILLER_23_3019 ();
 sg13g2_fill_2 FILLER_23_3023 ();
 sg13g2_fill_2 FILLER_23_3032 ();
 sg13g2_decap_8 FILLER_23_3038 ();
 sg13g2_fill_1 FILLER_23_3045 ();
 sg13g2_fill_2 FILLER_23_3063 ();
 sg13g2_decap_4 FILLER_23_3111 ();
 sg13g2_fill_1 FILLER_23_3115 ();
 sg13g2_fill_2 FILLER_23_3161 ();
 sg13g2_fill_1 FILLER_23_3199 ();
 sg13g2_decap_8 FILLER_23_3204 ();
 sg13g2_fill_2 FILLER_23_3263 ();
 sg13g2_fill_1 FILLER_23_3265 ();
 sg13g2_decap_4 FILLER_23_3292 ();
 sg13g2_fill_2 FILLER_23_3296 ();
 sg13g2_fill_1 FILLER_23_3324 ();
 sg13g2_decap_8 FILLER_23_3334 ();
 sg13g2_fill_2 FILLER_23_3341 ();
 sg13g2_fill_1 FILLER_23_3343 ();
 sg13g2_fill_2 FILLER_23_3375 ();
 sg13g2_decap_8 FILLER_23_3381 ();
 sg13g2_decap_4 FILLER_23_3388 ();
 sg13g2_fill_2 FILLER_23_3392 ();
 sg13g2_fill_2 FILLER_23_3434 ();
 sg13g2_fill_1 FILLER_23_3440 ();
 sg13g2_decap_4 FILLER_23_3450 ();
 sg13g2_fill_2 FILLER_23_3484 ();
 sg13g2_fill_1 FILLER_23_3486 ();
 sg13g2_decap_4 FILLER_23_3490 ();
 sg13g2_fill_2 FILLER_23_3494 ();
 sg13g2_fill_2 FILLER_23_3500 ();
 sg13g2_fill_2 FILLER_23_3516 ();
 sg13g2_fill_1 FILLER_23_3518 ();
 sg13g2_fill_2 FILLER_23_3545 ();
 sg13g2_decap_8 FILLER_23_3573 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_48 ();
 sg13g2_fill_1 FILLER_24_55 ();
 sg13g2_fill_2 FILLER_24_82 ();
 sg13g2_fill_1 FILLER_24_84 ();
 sg13g2_fill_1 FILLER_24_103 ();
 sg13g2_fill_2 FILLER_24_117 ();
 sg13g2_fill_2 FILLER_24_157 ();
 sg13g2_fill_2 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_fill_2 FILLER_24_291 ();
 sg13g2_fill_1 FILLER_24_306 ();
 sg13g2_decap_8 FILLER_24_324 ();
 sg13g2_fill_1 FILLER_24_331 ();
 sg13g2_fill_2 FILLER_24_359 ();
 sg13g2_fill_2 FILLER_24_380 ();
 sg13g2_fill_1 FILLER_24_382 ();
 sg13g2_decap_8 FILLER_24_409 ();
 sg13g2_decap_8 FILLER_24_416 ();
 sg13g2_decap_4 FILLER_24_423 ();
 sg13g2_fill_2 FILLER_24_440 ();
 sg13g2_fill_1 FILLER_24_442 ();
 sg13g2_decap_8 FILLER_24_469 ();
 sg13g2_fill_1 FILLER_24_502 ();
 sg13g2_decap_4 FILLER_24_512 ();
 sg13g2_fill_1 FILLER_24_528 ();
 sg13g2_fill_1 FILLER_24_538 ();
 sg13g2_fill_2 FILLER_24_548 ();
 sg13g2_fill_2 FILLER_24_559 ();
 sg13g2_fill_1 FILLER_24_561 ();
 sg13g2_fill_2 FILLER_24_574 ();
 sg13g2_fill_2 FILLER_24_606 ();
 sg13g2_fill_2 FILLER_24_616 ();
 sg13g2_fill_2 FILLER_24_623 ();
 sg13g2_fill_2 FILLER_24_651 ();
 sg13g2_decap_8 FILLER_24_696 ();
 sg13g2_fill_2 FILLER_24_703 ();
 sg13g2_fill_1 FILLER_24_709 ();
 sg13g2_fill_2 FILLER_24_776 ();
 sg13g2_fill_1 FILLER_24_778 ();
 sg13g2_fill_1 FILLER_24_783 ();
 sg13g2_decap_8 FILLER_24_797 ();
 sg13g2_decap_4 FILLER_24_804 ();
 sg13g2_fill_1 FILLER_24_808 ();
 sg13g2_decap_8 FILLER_24_817 ();
 sg13g2_fill_2 FILLER_24_824 ();
 sg13g2_fill_2 FILLER_24_861 ();
 sg13g2_fill_2 FILLER_24_889 ();
 sg13g2_fill_1 FILLER_24_891 ();
 sg13g2_fill_2 FILLER_24_918 ();
 sg13g2_decap_8 FILLER_24_961 ();
 sg13g2_decap_8 FILLER_24_972 ();
 sg13g2_decap_4 FILLER_24_979 ();
 sg13g2_fill_1 FILLER_24_983 ();
 sg13g2_fill_1 FILLER_24_1037 ();
 sg13g2_decap_4 FILLER_24_1090 ();
 sg13g2_fill_2 FILLER_24_1094 ();
 sg13g2_decap_8 FILLER_24_1122 ();
 sg13g2_fill_2 FILLER_24_1129 ();
 sg13g2_fill_2 FILLER_24_1135 ();
 sg13g2_decap_8 FILLER_24_1168 ();
 sg13g2_decap_4 FILLER_24_1175 ();
 sg13g2_fill_1 FILLER_24_1179 ();
 sg13g2_fill_2 FILLER_24_1211 ();
 sg13g2_fill_2 FILLER_24_1218 ();
 sg13g2_fill_1 FILLER_24_1269 ();
 sg13g2_fill_2 FILLER_24_1314 ();
 sg13g2_decap_8 FILLER_24_1342 ();
 sg13g2_decap_4 FILLER_24_1353 ();
 sg13g2_fill_1 FILLER_24_1357 ();
 sg13g2_fill_1 FILLER_24_1415 ();
 sg13g2_decap_8 FILLER_24_1426 ();
 sg13g2_fill_2 FILLER_24_1433 ();
 sg13g2_fill_2 FILLER_24_1446 ();
 sg13g2_fill_1 FILLER_24_1448 ();
 sg13g2_fill_2 FILLER_24_1457 ();
 sg13g2_fill_1 FILLER_24_1459 ();
 sg13g2_fill_2 FILLER_24_1464 ();
 sg13g2_fill_1 FILLER_24_1466 ();
 sg13g2_fill_2 FILLER_24_1472 ();
 sg13g2_fill_1 FILLER_24_1474 ();
 sg13g2_decap_4 FILLER_24_1480 ();
 sg13g2_decap_4 FILLER_24_1489 ();
 sg13g2_fill_1 FILLER_24_1493 ();
 sg13g2_decap_8 FILLER_24_1507 ();
 sg13g2_decap_4 FILLER_24_1514 ();
 sg13g2_fill_1 FILLER_24_1518 ();
 sg13g2_decap_4 FILLER_24_1536 ();
 sg13g2_fill_2 FILLER_24_1540 ();
 sg13g2_decap_8 FILLER_24_1608 ();
 sg13g2_fill_2 FILLER_24_1615 ();
 sg13g2_fill_1 FILLER_24_1617 ();
 sg13g2_fill_2 FILLER_24_1627 ();
 sg13g2_fill_1 FILLER_24_1629 ();
 sg13g2_decap_4 FILLER_24_1661 ();
 sg13g2_fill_1 FILLER_24_1665 ();
 sg13g2_fill_2 FILLER_24_1718 ();
 sg13g2_fill_1 FILLER_24_1729 ();
 sg13g2_decap_4 FILLER_24_1743 ();
 sg13g2_decap_8 FILLER_24_1773 ();
 sg13g2_decap_4 FILLER_24_1780 ();
 sg13g2_fill_2 FILLER_24_1784 ();
 sg13g2_fill_2 FILLER_24_1793 ();
 sg13g2_fill_2 FILLER_24_1803 ();
 sg13g2_fill_1 FILLER_24_1805 ();
 sg13g2_decap_4 FILLER_24_1815 ();
 sg13g2_fill_2 FILLER_24_1823 ();
 sg13g2_decap_8 FILLER_24_1828 ();
 sg13g2_fill_1 FILLER_24_1835 ();
 sg13g2_decap_8 FILLER_24_1840 ();
 sg13g2_decap_8 FILLER_24_1847 ();
 sg13g2_decap_4 FILLER_24_1854 ();
 sg13g2_decap_4 FILLER_24_1862 ();
 sg13g2_fill_1 FILLER_24_1866 ();
 sg13g2_fill_2 FILLER_24_1871 ();
 sg13g2_fill_1 FILLER_24_1873 ();
 sg13g2_fill_2 FILLER_24_1878 ();
 sg13g2_decap_4 FILLER_24_1903 ();
 sg13g2_decap_8 FILLER_24_1937 ();
 sg13g2_fill_2 FILLER_24_1970 ();
 sg13g2_decap_4 FILLER_24_1998 ();
 sg13g2_fill_2 FILLER_24_2010 ();
 sg13g2_fill_2 FILLER_24_2022 ();
 sg13g2_fill_1 FILLER_24_2024 ();
 sg13g2_fill_2 FILLER_24_2083 ();
 sg13g2_decap_8 FILLER_24_2089 ();
 sg13g2_decap_8 FILLER_24_2096 ();
 sg13g2_decap_4 FILLER_24_2103 ();
 sg13g2_fill_1 FILLER_24_2107 ();
 sg13g2_fill_1 FILLER_24_2113 ();
 sg13g2_fill_2 FILLER_24_2167 ();
 sg13g2_fill_1 FILLER_24_2204 ();
 sg13g2_fill_1 FILLER_24_2226 ();
 sg13g2_decap_4 FILLER_24_2236 ();
 sg13g2_decap_4 FILLER_24_2253 ();
 sg13g2_fill_2 FILLER_24_2283 ();
 sg13g2_fill_1 FILLER_24_2320 ();
 sg13g2_fill_2 FILLER_24_2369 ();
 sg13g2_decap_8 FILLER_24_2398 ();
 sg13g2_decap_8 FILLER_24_2405 ();
 sg13g2_fill_1 FILLER_24_2412 ();
 sg13g2_decap_4 FILLER_24_2432 ();
 sg13g2_fill_1 FILLER_24_2436 ();
 sg13g2_fill_2 FILLER_24_2457 ();
 sg13g2_decap_4 FILLER_24_2468 ();
 sg13g2_fill_1 FILLER_24_2472 ();
 sg13g2_decap_8 FILLER_24_2483 ();
 sg13g2_decap_8 FILLER_24_2490 ();
 sg13g2_decap_8 FILLER_24_2497 ();
 sg13g2_decap_4 FILLER_24_2504 ();
 sg13g2_fill_2 FILLER_24_2513 ();
 sg13g2_fill_1 FILLER_24_2515 ();
 sg13g2_fill_1 FILLER_24_2563 ();
 sg13g2_decap_8 FILLER_24_2582 ();
 sg13g2_decap_8 FILLER_24_2599 ();
 sg13g2_decap_4 FILLER_24_2631 ();
 sg13g2_fill_2 FILLER_24_2666 ();
 sg13g2_fill_1 FILLER_24_2668 ();
 sg13g2_fill_1 FILLER_24_2681 ();
 sg13g2_decap_8 FILLER_24_2688 ();
 sg13g2_decap_8 FILLER_24_2738 ();
 sg13g2_fill_2 FILLER_24_2771 ();
 sg13g2_fill_1 FILLER_24_2773 ();
 sg13g2_decap_8 FILLER_24_2790 ();
 sg13g2_decap_8 FILLER_24_2797 ();
 sg13g2_fill_1 FILLER_24_2811 ();
 sg13g2_decap_8 FILLER_24_2857 ();
 sg13g2_decap_8 FILLER_24_2864 ();
 sg13g2_decap_4 FILLER_24_2871 ();
 sg13g2_fill_2 FILLER_24_2875 ();
 sg13g2_fill_2 FILLER_24_2895 ();
 sg13g2_fill_1 FILLER_24_2897 ();
 sg13g2_decap_8 FILLER_24_2906 ();
 sg13g2_decap_4 FILLER_24_2913 ();
 sg13g2_fill_2 FILLER_24_2917 ();
 sg13g2_decap_4 FILLER_24_2935 ();
 sg13g2_fill_1 FILLER_24_2939 ();
 sg13g2_decap_4 FILLER_24_2954 ();
 sg13g2_fill_2 FILLER_24_2962 ();
 sg13g2_fill_1 FILLER_24_2964 ();
 sg13g2_decap_4 FILLER_24_3021 ();
 sg13g2_fill_1 FILLER_24_3025 ();
 sg13g2_fill_2 FILLER_24_3057 ();
 sg13g2_fill_1 FILLER_24_3059 ();
 sg13g2_decap_4 FILLER_24_3065 ();
 sg13g2_fill_1 FILLER_24_3069 ();
 sg13g2_fill_2 FILLER_24_3079 ();
 sg13g2_fill_2 FILLER_24_3095 ();
 sg13g2_decap_8 FILLER_24_3119 ();
 sg13g2_fill_2 FILLER_24_3130 ();
 sg13g2_decap_8 FILLER_24_3136 ();
 sg13g2_decap_8 FILLER_24_3143 ();
 sg13g2_decap_4 FILLER_24_3150 ();
 sg13g2_fill_2 FILLER_24_3154 ();
 sg13g2_fill_2 FILLER_24_3165 ();
 sg13g2_fill_1 FILLER_24_3167 ();
 sg13g2_fill_1 FILLER_24_3177 ();
 sg13g2_fill_2 FILLER_24_3204 ();
 sg13g2_fill_2 FILLER_24_3241 ();
 sg13g2_fill_1 FILLER_24_3243 ();
 sg13g2_fill_2 FILLER_24_3253 ();
 sg13g2_decap_8 FILLER_24_3263 ();
 sg13g2_decap_8 FILLER_24_3270 ();
 sg13g2_decap_8 FILLER_24_3280 ();
 sg13g2_fill_2 FILLER_24_3287 ();
 sg13g2_fill_2 FILLER_24_3307 ();
 sg13g2_fill_2 FILLER_24_3313 ();
 sg13g2_decap_4 FILLER_24_3351 ();
 sg13g2_fill_1 FILLER_24_3364 ();
 sg13g2_decap_8 FILLER_24_3374 ();
 sg13g2_decap_4 FILLER_24_3381 ();
 sg13g2_fill_1 FILLER_24_3385 ();
 sg13g2_fill_2 FILLER_24_3395 ();
 sg13g2_fill_2 FILLER_24_3415 ();
 sg13g2_fill_1 FILLER_24_3417 ();
 sg13g2_fill_2 FILLER_24_3423 ();
 sg13g2_fill_1 FILLER_24_3425 ();
 sg13g2_fill_2 FILLER_24_3444 ();
 sg13g2_fill_2 FILLER_24_3481 ();
 sg13g2_fill_1 FILLER_24_3483 ();
 sg13g2_fill_1 FILLER_24_3489 ();
 sg13g2_fill_2 FILLER_24_3498 ();
 sg13g2_decap_4 FILLER_24_3510 ();
 sg13g2_fill_2 FILLER_24_3528 ();
 sg13g2_fill_1 FILLER_24_3530 ();
 sg13g2_decap_4 FILLER_24_3536 ();
 sg13g2_fill_1 FILLER_24_3540 ();
 sg13g2_decap_4 FILLER_24_3545 ();
 sg13g2_fill_1 FILLER_24_3549 ();
 sg13g2_fill_2 FILLER_25_23 ();
 sg13g2_fill_1 FILLER_25_25 ();
 sg13g2_fill_2 FILLER_25_59 ();
 sg13g2_decap_8 FILLER_25_115 ();
 sg13g2_decap_8 FILLER_25_122 ();
 sg13g2_fill_1 FILLER_25_129 ();
 sg13g2_fill_1 FILLER_25_162 ();
 sg13g2_decap_4 FILLER_25_176 ();
 sg13g2_fill_1 FILLER_25_180 ();
 sg13g2_fill_2 FILLER_25_185 ();
 sg13g2_fill_1 FILLER_25_187 ();
 sg13g2_decap_4 FILLER_25_192 ();
 sg13g2_fill_1 FILLER_25_196 ();
 sg13g2_fill_2 FILLER_25_201 ();
 sg13g2_fill_1 FILLER_25_220 ();
 sg13g2_fill_2 FILLER_25_275 ();
 sg13g2_fill_1 FILLER_25_293 ();
 sg13g2_fill_2 FILLER_25_304 ();
 sg13g2_decap_4 FILLER_25_310 ();
 sg13g2_fill_1 FILLER_25_347 ();
 sg13g2_fill_2 FILLER_25_352 ();
 sg13g2_fill_1 FILLER_25_354 ();
 sg13g2_fill_2 FILLER_25_386 ();
 sg13g2_fill_1 FILLER_25_388 ();
 sg13g2_fill_1 FILLER_25_394 ();
 sg13g2_decap_4 FILLER_25_447 ();
 sg13g2_fill_2 FILLER_25_451 ();
 sg13g2_decap_8 FILLER_25_467 ();
 sg13g2_decap_8 FILLER_25_474 ();
 sg13g2_fill_2 FILLER_25_481 ();
 sg13g2_fill_1 FILLER_25_486 ();
 sg13g2_decap_8 FILLER_25_535 ();
 sg13g2_decap_8 FILLER_25_542 ();
 sg13g2_fill_2 FILLER_25_579 ();
 sg13g2_decap_8 FILLER_25_607 ();
 sg13g2_fill_2 FILLER_25_614 ();
 sg13g2_decap_8 FILLER_25_642 ();
 sg13g2_fill_1 FILLER_25_649 ();
 sg13g2_fill_1 FILLER_25_675 ();
 sg13g2_fill_2 FILLER_25_684 ();
 sg13g2_fill_1 FILLER_25_686 ();
 sg13g2_decap_4 FILLER_25_700 ();
 sg13g2_fill_2 FILLER_25_704 ();
 sg13g2_fill_2 FILLER_25_715 ();
 sg13g2_fill_2 FILLER_25_722 ();
 sg13g2_fill_1 FILLER_25_724 ();
 sg13g2_decap_8 FILLER_25_729 ();
 sg13g2_fill_2 FILLER_25_736 ();
 sg13g2_fill_1 FILLER_25_738 ();
 sg13g2_decap_4 FILLER_25_752 ();
 sg13g2_fill_1 FILLER_25_756 ();
 sg13g2_fill_2 FILLER_25_766 ();
 sg13g2_fill_2 FILLER_25_794 ();
 sg13g2_fill_1 FILLER_25_796 ();
 sg13g2_fill_2 FILLER_25_837 ();
 sg13g2_fill_1 FILLER_25_839 ();
 sg13g2_decap_8 FILLER_25_853 ();
 sg13g2_fill_1 FILLER_25_873 ();
 sg13g2_decap_8 FILLER_25_878 ();
 sg13g2_decap_4 FILLER_25_885 ();
 sg13g2_decap_8 FILLER_25_894 ();
 sg13g2_decap_8 FILLER_25_901 ();
 sg13g2_fill_1 FILLER_25_948 ();
 sg13g2_decap_8 FILLER_25_958 ();
 sg13g2_fill_1 FILLER_25_973 ();
 sg13g2_fill_1 FILLER_25_1000 ();
 sg13g2_fill_2 FILLER_25_1015 ();
 sg13g2_decap_4 FILLER_25_1110 ();
 sg13g2_fill_2 FILLER_25_1114 ();
 sg13g2_fill_2 FILLER_25_1142 ();
 sg13g2_fill_1 FILLER_25_1144 ();
 sg13g2_fill_2 FILLER_25_1163 ();
 sg13g2_decap_8 FILLER_25_1169 ();
 sg13g2_decap_8 FILLER_25_1176 ();
 sg13g2_decap_4 FILLER_25_1183 ();
 sg13g2_decap_8 FILLER_25_1195 ();
 sg13g2_fill_2 FILLER_25_1202 ();
 sg13g2_decap_8 FILLER_25_1207 ();
 sg13g2_fill_2 FILLER_25_1214 ();
 sg13g2_fill_1 FILLER_25_1249 ();
 sg13g2_fill_2 FILLER_25_1281 ();
 sg13g2_fill_1 FILLER_25_1283 ();
 sg13g2_decap_8 FILLER_25_1290 ();
 sg13g2_fill_2 FILLER_25_1310 ();
 sg13g2_decap_4 FILLER_25_1338 ();
 sg13g2_fill_1 FILLER_25_1342 ();
 sg13g2_fill_2 FILLER_25_1359 ();
 sg13g2_fill_1 FILLER_25_1361 ();
 sg13g2_decap_4 FILLER_25_1366 ();
 sg13g2_fill_2 FILLER_25_1370 ();
 sg13g2_decap_8 FILLER_25_1395 ();
 sg13g2_fill_2 FILLER_25_1402 ();
 sg13g2_fill_2 FILLER_25_1461 ();
 sg13g2_fill_1 FILLER_25_1463 ();
 sg13g2_fill_2 FILLER_25_1490 ();
 sg13g2_fill_2 FILLER_25_1544 ();
 sg13g2_fill_2 FILLER_25_1577 ();
 sg13g2_fill_2 FILLER_25_1605 ();
 sg13g2_decap_8 FILLER_25_1633 ();
 sg13g2_fill_2 FILLER_25_1644 ();
 sg13g2_fill_1 FILLER_25_1646 ();
 sg13g2_fill_1 FILLER_25_1661 ();
 sg13g2_decap_8 FILLER_25_1670 ();
 sg13g2_fill_2 FILLER_25_1677 ();
 sg13g2_decap_8 FILLER_25_1705 ();
 sg13g2_fill_2 FILLER_25_1712 ();
 sg13g2_decap_8 FILLER_25_1719 ();
 sg13g2_decap_8 FILLER_25_1726 ();
 sg13g2_decap_8 FILLER_25_1759 ();
 sg13g2_decap_4 FILLER_25_1766 ();
 sg13g2_decap_8 FILLER_25_1923 ();
 sg13g2_decap_8 FILLER_25_1930 ();
 sg13g2_decap_8 FILLER_25_1937 ();
 sg13g2_decap_8 FILLER_25_1944 ();
 sg13g2_fill_1 FILLER_25_1951 ();
 sg13g2_fill_1 FILLER_25_1961 ();
 sg13g2_fill_1 FILLER_25_1967 ();
 sg13g2_fill_1 FILLER_25_1996 ();
 sg13g2_decap_8 FILLER_25_2028 ();
 sg13g2_fill_1 FILLER_25_2035 ();
 sg13g2_decap_8 FILLER_25_2053 ();
 sg13g2_decap_4 FILLER_25_2060 ();
 sg13g2_fill_1 FILLER_25_2064 ();
 sg13g2_decap_4 FILLER_25_2069 ();
 sg13g2_fill_1 FILLER_25_2073 ();
 sg13g2_fill_2 FILLER_25_2100 ();
 sg13g2_fill_1 FILLER_25_2102 ();
 sg13g2_decap_8 FILLER_25_2129 ();
 sg13g2_decap_8 FILLER_25_2136 ();
 sg13g2_fill_1 FILLER_25_2147 ();
 sg13g2_decap_8 FILLER_25_2153 ();
 sg13g2_fill_2 FILLER_25_2165 ();
 sg13g2_fill_1 FILLER_25_2167 ();
 sg13g2_decap_8 FILLER_25_2172 ();
 sg13g2_fill_1 FILLER_25_2179 ();
 sg13g2_decap_8 FILLER_25_2184 ();
 sg13g2_fill_2 FILLER_25_2191 ();
 sg13g2_decap_8 FILLER_25_2217 ();
 sg13g2_decap_4 FILLER_25_2224 ();
 sg13g2_fill_1 FILLER_25_2228 ();
 sg13g2_decap_4 FILLER_25_2259 ();
 sg13g2_fill_2 FILLER_25_2272 ();
 sg13g2_fill_1 FILLER_25_2274 ();
 sg13g2_fill_1 FILLER_25_2279 ();
 sg13g2_decap_8 FILLER_25_2289 ();
 sg13g2_decap_8 FILLER_25_2300 ();
 sg13g2_fill_2 FILLER_25_2307 ();
 sg13g2_fill_1 FILLER_25_2309 ();
 sg13g2_fill_1 FILLER_25_2315 ();
 sg13g2_decap_8 FILLER_25_2329 ();
 sg13g2_decap_4 FILLER_25_2336 ();
 sg13g2_fill_1 FILLER_25_2340 ();
 sg13g2_fill_1 FILLER_25_2376 ();
 sg13g2_decap_4 FILLER_25_2391 ();
 sg13g2_fill_2 FILLER_25_2395 ();
 sg13g2_fill_2 FILLER_25_2405 ();
 sg13g2_fill_1 FILLER_25_2407 ();
 sg13g2_fill_2 FILLER_25_2432 ();
 sg13g2_fill_1 FILLER_25_2434 ();
 sg13g2_fill_1 FILLER_25_2442 ();
 sg13g2_fill_1 FILLER_25_2455 ();
 sg13g2_fill_2 FILLER_25_2466 ();
 sg13g2_decap_4 FILLER_25_2491 ();
 sg13g2_fill_2 FILLER_25_2495 ();
 sg13g2_fill_1 FILLER_25_2505 ();
 sg13g2_decap_4 FILLER_25_2566 ();
 sg13g2_fill_1 FILLER_25_2574 ();
 sg13g2_fill_1 FILLER_25_2610 ();
 sg13g2_fill_2 FILLER_25_2619 ();
 sg13g2_fill_1 FILLER_25_2629 ();
 sg13g2_decap_4 FILLER_25_2635 ();
 sg13g2_fill_2 FILLER_25_2639 ();
 sg13g2_fill_2 FILLER_25_2649 ();
 sg13g2_decap_8 FILLER_25_2655 ();
 sg13g2_decap_8 FILLER_25_2662 ();
 sg13g2_decap_4 FILLER_25_2669 ();
 sg13g2_fill_1 FILLER_25_2673 ();
 sg13g2_decap_8 FILLER_25_2692 ();
 sg13g2_decap_8 FILLER_25_2699 ();
 sg13g2_decap_4 FILLER_25_2710 ();
 sg13g2_fill_2 FILLER_25_2740 ();
 sg13g2_fill_1 FILLER_25_2742 ();
 sg13g2_fill_2 FILLER_25_2748 ();
 sg13g2_fill_1 FILLER_25_2750 ();
 sg13g2_decap_8 FILLER_25_2755 ();
 sg13g2_decap_8 FILLER_25_2762 ();
 sg13g2_fill_1 FILLER_25_2769 ();
 sg13g2_decap_8 FILLER_25_2775 ();
 sg13g2_fill_2 FILLER_25_2786 ();
 sg13g2_fill_2 FILLER_25_2796 ();
 sg13g2_fill_1 FILLER_25_2798 ();
 sg13g2_fill_1 FILLER_25_2826 ();
 sg13g2_decap_8 FILLER_25_2831 ();
 sg13g2_fill_2 FILLER_25_2838 ();
 sg13g2_fill_1 FILLER_25_2840 ();
 sg13g2_fill_1 FILLER_25_2886 ();
 sg13g2_fill_1 FILLER_25_2913 ();
 sg13g2_decap_8 FILLER_25_2922 ();
 sg13g2_fill_1 FILLER_25_2942 ();
 sg13g2_decap_4 FILLER_25_2956 ();
 sg13g2_fill_1 FILLER_25_2960 ();
 sg13g2_decap_8 FILLER_25_2966 ();
 sg13g2_decap_8 FILLER_25_2973 ();
 sg13g2_decap_4 FILLER_25_2980 ();
 sg13g2_fill_1 FILLER_25_2984 ();
 sg13g2_decap_8 FILLER_25_2993 ();
 sg13g2_fill_1 FILLER_25_3000 ();
 sg13g2_decap_4 FILLER_25_3055 ();
 sg13g2_fill_2 FILLER_25_3067 ();
 sg13g2_fill_1 FILLER_25_3069 ();
 sg13g2_fill_2 FILLER_25_3096 ();
 sg13g2_fill_2 FILLER_25_3145 ();
 sg13g2_fill_1 FILLER_25_3147 ();
 sg13g2_fill_1 FILLER_25_3161 ();
 sg13g2_decap_8 FILLER_25_3188 ();
 sg13g2_decap_4 FILLER_25_3208 ();
 sg13g2_fill_1 FILLER_25_3212 ();
 sg13g2_decap_8 FILLER_25_3232 ();
 sg13g2_decap_4 FILLER_25_3239 ();
 sg13g2_fill_2 FILLER_25_3243 ();
 sg13g2_decap_8 FILLER_25_3295 ();
 sg13g2_decap_8 FILLER_25_3302 ();
 sg13g2_decap_8 FILLER_25_3309 ();
 sg13g2_decap_4 FILLER_25_3320 ();
 sg13g2_fill_1 FILLER_25_3324 ();
 sg13g2_decap_4 FILLER_25_3340 ();
 sg13g2_fill_2 FILLER_25_3344 ();
 sg13g2_fill_1 FILLER_25_3366 ();
 sg13g2_fill_1 FILLER_25_3458 ();
 sg13g2_fill_2 FILLER_25_3464 ();
 sg13g2_fill_2 FILLER_25_3531 ();
 sg13g2_fill_1 FILLER_25_3533 ();
 sg13g2_fill_2 FILLER_25_3569 ();
 sg13g2_fill_1 FILLER_26_26 ();
 sg13g2_fill_2 FILLER_26_45 ();
 sg13g2_fill_2 FILLER_26_61 ();
 sg13g2_fill_2 FILLER_26_87 ();
 sg13g2_fill_1 FILLER_26_98 ();
 sg13g2_fill_2 FILLER_26_108 ();
 sg13g2_fill_1 FILLER_26_114 ();
 sg13g2_decap_8 FILLER_26_128 ();
 sg13g2_decap_8 FILLER_26_135 ();
 sg13g2_fill_1 FILLER_26_142 ();
 sg13g2_fill_2 FILLER_26_183 ();
 sg13g2_fill_1 FILLER_26_185 ();
 sg13g2_fill_2 FILLER_26_229 ();
 sg13g2_fill_1 FILLER_26_231 ();
 sg13g2_fill_2 FILLER_26_254 ();
 sg13g2_fill_1 FILLER_26_256 ();
 sg13g2_fill_2 FILLER_26_289 ();
 sg13g2_decap_4 FILLER_26_295 ();
 sg13g2_fill_1 FILLER_26_362 ();
 sg13g2_fill_1 FILLER_26_439 ();
 sg13g2_fill_1 FILLER_26_444 ();
 sg13g2_fill_2 FILLER_26_448 ();
 sg13g2_fill_1 FILLER_26_450 ();
 sg13g2_fill_2 FILLER_26_503 ();
 sg13g2_fill_1 FILLER_26_573 ();
 sg13g2_decap_8 FILLER_26_623 ();
 sg13g2_decap_8 FILLER_26_630 ();
 sg13g2_decap_8 FILLER_26_637 ();
 sg13g2_decap_8 FILLER_26_644 ();
 sg13g2_decap_8 FILLER_26_677 ();
 sg13g2_decap_4 FILLER_26_684 ();
 sg13g2_fill_1 FILLER_26_719 ();
 sg13g2_fill_2 FILLER_26_725 ();
 sg13g2_fill_1 FILLER_26_727 ();
 sg13g2_fill_2 FILLER_26_767 ();
 sg13g2_fill_1 FILLER_26_769 ();
 sg13g2_fill_2 FILLER_26_783 ();
 sg13g2_decap_8 FILLER_26_807 ();
 sg13g2_fill_2 FILLER_26_845 ();
 sg13g2_fill_2 FILLER_26_873 ();
 sg13g2_fill_1 FILLER_26_901 ();
 sg13g2_fill_2 FILLER_26_910 ();
 sg13g2_fill_1 FILLER_26_912 ();
 sg13g2_fill_2 FILLER_26_930 ();
 sg13g2_decap_4 FILLER_26_954 ();
 sg13g2_fill_2 FILLER_26_984 ();
 sg13g2_fill_2 FILLER_26_1032 ();
 sg13g2_decap_4 FILLER_26_1065 ();
 sg13g2_fill_2 FILLER_26_1069 ();
 sg13g2_fill_2 FILLER_26_1084 ();
 sg13g2_fill_1 FILLER_26_1086 ();
 sg13g2_fill_2 FILLER_26_1092 ();
 sg13g2_fill_1 FILLER_26_1094 ();
 sg13g2_fill_2 FILLER_26_1118 ();
 sg13g2_fill_1 FILLER_26_1120 ();
 sg13g2_decap_8 FILLER_26_1134 ();
 sg13g2_fill_2 FILLER_26_1141 ();
 sg13g2_fill_1 FILLER_26_1143 ();
 sg13g2_fill_2 FILLER_26_1174 ();
 sg13g2_fill_2 FILLER_26_1207 ();
 sg13g2_fill_2 FILLER_26_1235 ();
 sg13g2_fill_1 FILLER_26_1237 ();
 sg13g2_decap_4 FILLER_26_1243 ();
 sg13g2_fill_2 FILLER_26_1247 ();
 sg13g2_fill_2 FILLER_26_1280 ();
 sg13g2_fill_2 FILLER_26_1287 ();
 sg13g2_fill_1 FILLER_26_1289 ();
 sg13g2_fill_1 FILLER_26_1294 ();
 sg13g2_decap_4 FILLER_26_1304 ();
 sg13g2_fill_2 FILLER_26_1349 ();
 sg13g2_fill_1 FILLER_26_1351 ();
 sg13g2_decap_4 FILLER_26_1392 ();
 sg13g2_decap_8 FILLER_26_1401 ();
 sg13g2_fill_2 FILLER_26_1408 ();
 sg13g2_decap_4 FILLER_26_1415 ();
 sg13g2_fill_1 FILLER_26_1419 ();
 sg13g2_decap_8 FILLER_26_1429 ();
 sg13g2_decap_4 FILLER_26_1436 ();
 sg13g2_fill_1 FILLER_26_1458 ();
 sg13g2_decap_8 FILLER_26_1464 ();
 sg13g2_decap_4 FILLER_26_1471 ();
 sg13g2_fill_2 FILLER_26_1498 ();
 sg13g2_fill_2 FILLER_26_1525 ();
 sg13g2_fill_1 FILLER_26_1527 ();
 sg13g2_fill_1 FILLER_26_1536 ();
 sg13g2_fill_1 FILLER_26_1546 ();
 sg13g2_fill_2 FILLER_26_1551 ();
 sg13g2_fill_1 FILLER_26_1553 ();
 sg13g2_fill_2 FILLER_26_1570 ();
 sg13g2_fill_1 FILLER_26_1572 ();
 sg13g2_fill_2 FILLER_26_1592 ();
 sg13g2_fill_1 FILLER_26_1594 ();
 sg13g2_fill_1 FILLER_26_1612 ();
 sg13g2_fill_2 FILLER_26_1636 ();
 sg13g2_decap_4 FILLER_26_1676 ();
 sg13g2_fill_2 FILLER_26_1680 ();
 sg13g2_decap_8 FILLER_26_1685 ();
 sg13g2_decap_8 FILLER_26_1692 ();
 sg13g2_decap_4 FILLER_26_1699 ();
 sg13g2_fill_2 FILLER_26_1703 ();
 sg13g2_decap_8 FILLER_26_1731 ();
 sg13g2_decap_8 FILLER_26_1738 ();
 sg13g2_fill_2 FILLER_26_1745 ();
 sg13g2_decap_8 FILLER_26_1755 ();
 sg13g2_decap_4 FILLER_26_1762 ();
 sg13g2_fill_2 FILLER_26_1779 ();
 sg13g2_fill_1 FILLER_26_1781 ();
 sg13g2_decap_8 FILLER_26_1789 ();
 sg13g2_decap_8 FILLER_26_1799 ();
 sg13g2_decap_8 FILLER_26_1806 ();
 sg13g2_decap_8 FILLER_26_1821 ();
 sg13g2_decap_8 FILLER_26_1828 ();
 sg13g2_decap_8 FILLER_26_1835 ();
 sg13g2_decap_4 FILLER_26_1842 ();
 sg13g2_fill_2 FILLER_26_1846 ();
 sg13g2_fill_2 FILLER_26_1861 ();
 sg13g2_decap_8 FILLER_26_1866 ();
 sg13g2_fill_2 FILLER_26_1878 ();
 sg13g2_fill_2 FILLER_26_1913 ();
 sg13g2_fill_2 FILLER_26_1919 ();
 sg13g2_fill_1 FILLER_26_1921 ();
 sg13g2_fill_2 FILLER_26_1931 ();
 sg13g2_fill_1 FILLER_26_1969 ();
 sg13g2_decap_4 FILLER_26_1984 ();
 sg13g2_decap_8 FILLER_26_2050 ();
 sg13g2_decap_8 FILLER_26_2057 ();
 sg13g2_fill_1 FILLER_26_2064 ();
 sg13g2_decap_8 FILLER_26_2091 ();
 sg13g2_decap_4 FILLER_26_2098 ();
 sg13g2_decap_8 FILLER_26_2106 ();
 sg13g2_fill_1 FILLER_26_2113 ();
 sg13g2_fill_2 FILLER_26_2122 ();
 sg13g2_decap_4 FILLER_26_2145 ();
 sg13g2_decap_8 FILLER_26_2227 ();
 sg13g2_decap_4 FILLER_26_2234 ();
 sg13g2_fill_2 FILLER_26_2238 ();
 sg13g2_fill_2 FILLER_26_2262 ();
 sg13g2_fill_1 FILLER_26_2264 ();
 sg13g2_decap_8 FILLER_26_2291 ();
 sg13g2_fill_2 FILLER_26_2302 ();
 sg13g2_fill_2 FILLER_26_2339 ();
 sg13g2_fill_1 FILLER_26_2345 ();
 sg13g2_fill_2 FILLER_26_2350 ();
 sg13g2_fill_2 FILLER_26_2356 ();
 sg13g2_fill_1 FILLER_26_2358 ();
 sg13g2_fill_2 FILLER_26_2372 ();
 sg13g2_decap_4 FILLER_26_2395 ();
 sg13g2_fill_1 FILLER_26_2399 ();
 sg13g2_fill_1 FILLER_26_2405 ();
 sg13g2_decap_8 FILLER_26_2426 ();
 sg13g2_decap_4 FILLER_26_2433 ();
 sg13g2_fill_2 FILLER_26_2437 ();
 sg13g2_fill_2 FILLER_26_2443 ();
 sg13g2_fill_1 FILLER_26_2445 ();
 sg13g2_decap_4 FILLER_26_2474 ();
 sg13g2_decap_8 FILLER_26_2483 ();
 sg13g2_decap_8 FILLER_26_2490 ();
 sg13g2_fill_2 FILLER_26_2497 ();
 sg13g2_fill_1 FILLER_26_2499 ();
 sg13g2_fill_1 FILLER_26_2509 ();
 sg13g2_fill_1 FILLER_26_2528 ();
 sg13g2_decap_8 FILLER_26_2576 ();
 sg13g2_decap_8 FILLER_26_2583 ();
 sg13g2_decap_4 FILLER_26_2590 ();
 sg13g2_fill_1 FILLER_26_2594 ();
 sg13g2_decap_8 FILLER_26_2600 ();
 sg13g2_decap_4 FILLER_26_2607 ();
 sg13g2_fill_1 FILLER_26_2611 ();
 sg13g2_decap_4 FILLER_26_2622 ();
 sg13g2_fill_2 FILLER_26_2626 ();
 sg13g2_fill_1 FILLER_26_2644 ();
 sg13g2_decap_8 FILLER_26_2651 ();
 sg13g2_decap_8 FILLER_26_2658 ();
 sg13g2_decap_4 FILLER_26_2675 ();
 sg13g2_fill_2 FILLER_26_2679 ();
 sg13g2_decap_4 FILLER_26_2689 ();
 sg13g2_fill_2 FILLER_26_2693 ();
 sg13g2_fill_2 FILLER_26_2700 ();
 sg13g2_decap_8 FILLER_26_2710 ();
 sg13g2_fill_2 FILLER_26_2717 ();
 sg13g2_fill_1 FILLER_26_2719 ();
 sg13g2_fill_2 FILLER_26_2730 ();
 sg13g2_decap_8 FILLER_26_2763 ();
 sg13g2_decap_8 FILLER_26_2770 ();
 sg13g2_fill_2 FILLER_26_2791 ();
 sg13g2_fill_1 FILLER_26_2793 ();
 sg13g2_decap_4 FILLER_26_2800 ();
 sg13g2_fill_2 FILLER_26_2813 ();
 sg13g2_fill_1 FILLER_26_2815 ();
 sg13g2_fill_1 FILLER_26_2821 ();
 sg13g2_fill_1 FILLER_26_2827 ();
 sg13g2_decap_8 FILLER_26_2841 ();
 sg13g2_decap_4 FILLER_26_2848 ();
 sg13g2_decap_8 FILLER_26_2856 ();
 sg13g2_decap_8 FILLER_26_2863 ();
 sg13g2_fill_2 FILLER_26_2870 ();
 sg13g2_fill_1 FILLER_26_2877 ();
 sg13g2_fill_2 FILLER_26_2887 ();
 sg13g2_decap_8 FILLER_26_2920 ();
 sg13g2_decap_8 FILLER_26_2927 ();
 sg13g2_fill_1 FILLER_26_2934 ();
 sg13g2_decap_8 FILLER_26_2940 ();
 sg13g2_decap_8 FILLER_26_2947 ();
 sg13g2_fill_2 FILLER_26_2954 ();
 sg13g2_decap_8 FILLER_26_2964 ();
 sg13g2_fill_2 FILLER_26_2971 ();
 sg13g2_fill_1 FILLER_26_2973 ();
 sg13g2_decap_8 FILLER_26_3022 ();
 sg13g2_decap_8 FILLER_26_3065 ();
 sg13g2_decap_4 FILLER_26_3072 ();
 sg13g2_fill_2 FILLER_26_3076 ();
 sg13g2_fill_2 FILLER_26_3091 ();
 sg13g2_decap_8 FILLER_26_3134 ();
 sg13g2_decap_8 FILLER_26_3141 ();
 sg13g2_fill_1 FILLER_26_3148 ();
 sg13g2_decap_8 FILLER_26_3162 ();
 sg13g2_decap_4 FILLER_26_3169 ();
 sg13g2_fill_1 FILLER_26_3183 ();
 sg13g2_fill_2 FILLER_26_3194 ();
 sg13g2_fill_1 FILLER_26_3196 ();
 sg13g2_fill_1 FILLER_26_3210 ();
 sg13g2_decap_4 FILLER_26_3215 ();
 sg13g2_fill_2 FILLER_26_3219 ();
 sg13g2_fill_2 FILLER_26_3242 ();
 sg13g2_fill_2 FILLER_26_3253 ();
 sg13g2_fill_1 FILLER_26_3255 ();
 sg13g2_fill_1 FILLER_26_3260 ();
 sg13g2_decap_8 FILLER_26_3270 ();
 sg13g2_fill_2 FILLER_26_3277 ();
 sg13g2_fill_1 FILLER_26_3313 ();
 sg13g2_decap_8 FILLER_26_3348 ();
 sg13g2_decap_8 FILLER_26_3359 ();
 sg13g2_decap_4 FILLER_26_3366 ();
 sg13g2_decap_4 FILLER_26_3406 ();
 sg13g2_fill_2 FILLER_26_3410 ();
 sg13g2_fill_2 FILLER_26_3417 ();
 sg13g2_fill_1 FILLER_26_3419 ();
 sg13g2_fill_2 FILLER_26_3429 ();
 sg13g2_fill_1 FILLER_26_3431 ();
 sg13g2_fill_1 FILLER_26_3446 ();
 sg13g2_fill_2 FILLER_26_3473 ();
 sg13g2_fill_2 FILLER_26_3480 ();
 sg13g2_fill_1 FILLER_26_3482 ();
 sg13g2_fill_2 FILLER_26_3488 ();
 sg13g2_fill_1 FILLER_26_3490 ();
 sg13g2_fill_2 FILLER_26_3500 ();
 sg13g2_fill_1 FILLER_26_3502 ();
 sg13g2_fill_1 FILLER_26_3516 ();
 sg13g2_decap_4 FILLER_26_3526 ();
 sg13g2_fill_1 FILLER_26_3530 ();
 sg13g2_fill_1 FILLER_26_3544 ();
 sg13g2_decap_4 FILLER_26_3553 ();
 sg13g2_fill_1 FILLER_26_3557 ();
 sg13g2_decap_4 FILLER_26_3575 ();
 sg13g2_fill_1 FILLER_26_3579 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_fill_2 FILLER_27_14 ();
 sg13g2_fill_1 FILLER_27_16 ();
 sg13g2_fill_1 FILLER_27_41 ();
 sg13g2_fill_2 FILLER_27_53 ();
 sg13g2_fill_1 FILLER_27_90 ();
 sg13g2_fill_2 FILLER_27_139 ();
 sg13g2_decap_4 FILLER_27_145 ();
 sg13g2_decap_8 FILLER_27_179 ();
 sg13g2_decap_8 FILLER_27_186 ();
 sg13g2_fill_1 FILLER_27_193 ();
 sg13g2_decap_4 FILLER_27_198 ();
 sg13g2_fill_1 FILLER_27_202 ();
 sg13g2_fill_1 FILLER_27_221 ();
 sg13g2_decap_4 FILLER_27_227 ();
 sg13g2_fill_2 FILLER_27_231 ();
 sg13g2_fill_2 FILLER_27_243 ();
 sg13g2_fill_1 FILLER_27_259 ();
 sg13g2_decap_8 FILLER_27_336 ();
 sg13g2_fill_1 FILLER_27_343 ();
 sg13g2_fill_2 FILLER_27_347 ();
 sg13g2_decap_4 FILLER_27_358 ();
 sg13g2_fill_2 FILLER_27_362 ();
 sg13g2_fill_2 FILLER_27_390 ();
 sg13g2_fill_1 FILLER_27_424 ();
 sg13g2_fill_2 FILLER_27_482 ();
 sg13g2_fill_1 FILLER_27_493 ();
 sg13g2_decap_8 FILLER_27_546 ();
 sg13g2_decap_4 FILLER_27_553 ();
 sg13g2_fill_1 FILLER_27_561 ();
 sg13g2_decap_8 FILLER_27_599 ();
 sg13g2_fill_2 FILLER_27_606 ();
 sg13g2_decap_8 FILLER_27_612 ();
 sg13g2_fill_2 FILLER_27_619 ();
 sg13g2_decap_4 FILLER_27_625 ();
 sg13g2_fill_1 FILLER_27_629 ();
 sg13g2_fill_1 FILLER_27_668 ();
 sg13g2_decap_4 FILLER_27_699 ();
 sg13g2_fill_1 FILLER_27_703 ();
 sg13g2_decap_8 FILLER_27_708 ();
 sg13g2_fill_2 FILLER_27_715 ();
 sg13g2_fill_1 FILLER_27_717 ();
 sg13g2_decap_4 FILLER_27_757 ();
 sg13g2_fill_2 FILLER_27_761 ();
 sg13g2_fill_1 FILLER_27_828 ();
 sg13g2_decap_4 FILLER_27_842 ();
 sg13g2_decap_8 FILLER_27_863 ();
 sg13g2_fill_2 FILLER_27_870 ();
 sg13g2_fill_1 FILLER_27_872 ();
 sg13g2_decap_4 FILLER_27_879 ();
 sg13g2_fill_2 FILLER_27_883 ();
 sg13g2_fill_2 FILLER_27_889 ();
 sg13g2_fill_1 FILLER_27_891 ();
 sg13g2_fill_1 FILLER_27_896 ();
 sg13g2_decap_8 FILLER_27_906 ();
 sg13g2_fill_1 FILLER_27_913 ();
 sg13g2_decap_8 FILLER_27_918 ();
 sg13g2_fill_1 FILLER_27_925 ();
 sg13g2_fill_2 FILLER_27_972 ();
 sg13g2_fill_1 FILLER_27_974 ();
 sg13g2_fill_1 FILLER_27_988 ();
 sg13g2_fill_2 FILLER_27_997 ();
 sg13g2_fill_1 FILLER_27_999 ();
 sg13g2_fill_2 FILLER_27_1008 ();
 sg13g2_fill_1 FILLER_27_1010 ();
 sg13g2_fill_1 FILLER_27_1016 ();
 sg13g2_decap_4 FILLER_27_1021 ();
 sg13g2_fill_2 FILLER_27_1059 ();
 sg13g2_fill_1 FILLER_27_1070 ();
 sg13g2_fill_1 FILLER_27_1091 ();
 sg13g2_fill_1 FILLER_27_1097 ();
 sg13g2_fill_1 FILLER_27_1112 ();
 sg13g2_decap_4 FILLER_27_1144 ();
 sg13g2_fill_1 FILLER_27_1148 ();
 sg13g2_fill_1 FILLER_27_1178 ();
 sg13g2_fill_2 FILLER_27_1193 ();
 sg13g2_fill_2 FILLER_27_1215 ();
 sg13g2_fill_1 FILLER_27_1217 ();
 sg13g2_decap_8 FILLER_27_1243 ();
 sg13g2_fill_1 FILLER_27_1273 ();
 sg13g2_fill_2 FILLER_27_1305 ();
 sg13g2_fill_2 FILLER_27_1322 ();
 sg13g2_fill_1 FILLER_27_1324 ();
 sg13g2_fill_2 FILLER_27_1330 ();
 sg13g2_fill_1 FILLER_27_1332 ();
 sg13g2_fill_2 FILLER_27_1358 ();
 sg13g2_fill_1 FILLER_27_1360 ();
 sg13g2_decap_8 FILLER_27_1365 ();
 sg13g2_fill_2 FILLER_27_1372 ();
 sg13g2_fill_1 FILLER_27_1374 ();
 sg13g2_fill_2 FILLER_27_1379 ();
 sg13g2_fill_1 FILLER_27_1381 ();
 sg13g2_fill_2 FILLER_27_1396 ();
 sg13g2_fill_1 FILLER_27_1398 ();
 sg13g2_decap_4 FILLER_27_1411 ();
 sg13g2_fill_2 FILLER_27_1447 ();
 sg13g2_fill_1 FILLER_27_1449 ();
 sg13g2_decap_4 FILLER_27_1478 ();
 sg13g2_fill_1 FILLER_27_1496 ();
 sg13g2_decap_4 FILLER_27_1513 ();
 sg13g2_fill_1 FILLER_27_1517 ();
 sg13g2_fill_2 FILLER_27_1522 ();
 sg13g2_fill_2 FILLER_27_1542 ();
 sg13g2_fill_1 FILLER_27_1548 ();
 sg13g2_fill_2 FILLER_27_1573 ();
 sg13g2_fill_1 FILLER_27_1575 ();
 sg13g2_fill_2 FILLER_27_1613 ();
 sg13g2_fill_2 FILLER_27_1641 ();
 sg13g2_fill_2 FILLER_27_1671 ();
 sg13g2_decap_4 FILLER_27_1712 ();
 sg13g2_decap_8 FILLER_27_1720 ();
 sg13g2_fill_1 FILLER_27_1727 ();
 sg13g2_decap_4 FILLER_27_1732 ();
 sg13g2_decap_4 FILLER_27_1762 ();
 sg13g2_fill_2 FILLER_27_1766 ();
 sg13g2_decap_8 FILLER_27_1832 ();
 sg13g2_decap_4 FILLER_27_1905 ();
 sg13g2_fill_1 FILLER_27_1909 ();
 sg13g2_decap_8 FILLER_27_1920 ();
 sg13g2_decap_8 FILLER_27_1927 ();
 sg13g2_fill_2 FILLER_27_1942 ();
 sg13g2_fill_2 FILLER_27_1948 ();
 sg13g2_fill_2 FILLER_27_1959 ();
 sg13g2_fill_1 FILLER_27_1961 ();
 sg13g2_decap_8 FILLER_27_1973 ();
 sg13g2_decap_8 FILLER_27_1980 ();
 sg13g2_fill_2 FILLER_27_2010 ();
 sg13g2_fill_1 FILLER_27_2012 ();
 sg13g2_decap_8 FILLER_27_2040 ();
 sg13g2_fill_2 FILLER_27_2047 ();
 sg13g2_fill_1 FILLER_27_2049 ();
 sg13g2_fill_1 FILLER_27_2081 ();
 sg13g2_decap_8 FILLER_27_2117 ();
 sg13g2_decap_4 FILLER_27_2173 ();
 sg13g2_fill_1 FILLER_27_2177 ();
 sg13g2_fill_2 FILLER_27_2183 ();
 sg13g2_fill_1 FILLER_27_2204 ();
 sg13g2_decap_4 FILLER_27_2233 ();
 sg13g2_fill_1 FILLER_27_2237 ();
 sg13g2_decap_8 FILLER_27_2269 ();
 sg13g2_fill_1 FILLER_27_2276 ();
 sg13g2_fill_2 FILLER_27_2322 ();
 sg13g2_fill_1 FILLER_27_2324 ();
 sg13g2_fill_2 FILLER_27_2365 ();
 sg13g2_fill_1 FILLER_27_2367 ();
 sg13g2_decap_8 FILLER_27_2395 ();
 sg13g2_decap_4 FILLER_27_2402 ();
 sg13g2_fill_2 FILLER_27_2406 ();
 sg13g2_fill_1 FILLER_27_2429 ();
 sg13g2_fill_1 FILLER_27_2521 ();
 sg13g2_fill_2 FILLER_27_2565 ();
 sg13g2_fill_2 FILLER_27_2578 ();
 sg13g2_decap_4 FILLER_27_2593 ();
 sg13g2_fill_2 FILLER_27_2597 ();
 sg13g2_decap_8 FILLER_27_2621 ();
 sg13g2_fill_1 FILLER_27_2628 ();
 sg13g2_fill_2 FILLER_27_2634 ();
 sg13g2_fill_1 FILLER_27_2636 ();
 sg13g2_decap_4 FILLER_27_2645 ();
 sg13g2_fill_2 FILLER_27_2649 ();
 sg13g2_fill_1 FILLER_27_2672 ();
 sg13g2_decap_4 FILLER_27_2682 ();
 sg13g2_fill_1 FILLER_27_2686 ();
 sg13g2_fill_2 FILLER_27_2714 ();
 sg13g2_fill_1 FILLER_27_2716 ();
 sg13g2_fill_2 FILLER_27_2735 ();
 sg13g2_fill_1 FILLER_27_2737 ();
 sg13g2_fill_1 FILLER_27_2751 ();
 sg13g2_fill_1 FILLER_27_2788 ();
 sg13g2_fill_1 FILLER_27_2825 ();
 sg13g2_fill_1 FILLER_27_2852 ();
 sg13g2_fill_2 FILLER_27_2909 ();
 sg13g2_fill_1 FILLER_27_2911 ();
 sg13g2_fill_2 FILLER_27_2964 ();
 sg13g2_fill_1 FILLER_27_2966 ();
 sg13g2_decap_8 FILLER_27_2975 ();
 sg13g2_decap_4 FILLER_27_2982 ();
 sg13g2_decap_8 FILLER_27_2998 ();
 sg13g2_fill_1 FILLER_27_3005 ();
 sg13g2_fill_1 FILLER_27_3037 ();
 sg13g2_decap_4 FILLER_27_3057 ();
 sg13g2_fill_2 FILLER_27_3074 ();
 sg13g2_decap_8 FILLER_27_3144 ();
 sg13g2_fill_1 FILLER_27_3151 ();
 sg13g2_fill_1 FILLER_27_3191 ();
 sg13g2_fill_1 FILLER_27_3200 ();
 sg13g2_decap_8 FILLER_27_3227 ();
 sg13g2_decap_4 FILLER_27_3234 ();
 sg13g2_decap_8 FILLER_27_3269 ();
 sg13g2_fill_2 FILLER_27_3284 ();
 sg13g2_fill_1 FILLER_27_3286 ();
 sg13g2_fill_1 FILLER_27_3296 ();
 sg13g2_fill_2 FILLER_27_3301 ();
 sg13g2_fill_1 FILLER_27_3312 ();
 sg13g2_fill_1 FILLER_27_3327 ();
 sg13g2_fill_1 FILLER_27_3332 ();
 sg13g2_fill_2 FILLER_27_3337 ();
 sg13g2_fill_1 FILLER_27_3348 ();
 sg13g2_fill_1 FILLER_27_3384 ();
 sg13g2_fill_2 FILLER_27_3440 ();
 sg13g2_fill_2 FILLER_27_3455 ();
 sg13g2_decap_8 FILLER_27_3461 ();
 sg13g2_decap_4 FILLER_27_3468 ();
 sg13g2_fill_2 FILLER_27_3472 ();
 sg13g2_fill_2 FILLER_27_3489 ();
 sg13g2_fill_2 FILLER_27_3578 ();
 sg13g2_fill_2 FILLER_28_26 ();
 sg13g2_fill_1 FILLER_28_28 ();
 sg13g2_fill_1 FILLER_28_46 ();
 sg13g2_fill_1 FILLER_28_50 ();
 sg13g2_fill_2 FILLER_28_94 ();
 sg13g2_fill_1 FILLER_28_96 ();
 sg13g2_decap_4 FILLER_28_141 ();
 sg13g2_fill_2 FILLER_28_145 ();
 sg13g2_fill_2 FILLER_28_209 ();
 sg13g2_fill_1 FILLER_28_211 ();
 sg13g2_decap_4 FILLER_28_233 ();
 sg13g2_decap_8 FILLER_28_267 ();
 sg13g2_fill_1 FILLER_28_274 ();
 sg13g2_fill_1 FILLER_28_285 ();
 sg13g2_decap_4 FILLER_28_364 ();
 sg13g2_fill_1 FILLER_28_387 ();
 sg13g2_fill_2 FILLER_28_402 ();
 sg13g2_fill_2 FILLER_28_414 ();
 sg13g2_fill_1 FILLER_28_434 ();
 sg13g2_fill_2 FILLER_28_440 ();
 sg13g2_fill_1 FILLER_28_442 ();
 sg13g2_fill_1 FILLER_28_465 ();
 sg13g2_fill_1 FILLER_28_502 ();
 sg13g2_fill_1 FILLER_28_509 ();
 sg13g2_fill_1 FILLER_28_521 ();
 sg13g2_fill_2 FILLER_28_526 ();
 sg13g2_fill_1 FILLER_28_538 ();
 sg13g2_fill_2 FILLER_28_562 ();
 sg13g2_fill_1 FILLER_28_564 ();
 sg13g2_fill_2 FILLER_28_569 ();
 sg13g2_fill_1 FILLER_28_583 ();
 sg13g2_fill_2 FILLER_28_636 ();
 sg13g2_fill_1 FILLER_28_648 ();
 sg13g2_decap_8 FILLER_28_666 ();
 sg13g2_decap_8 FILLER_28_673 ();
 sg13g2_fill_2 FILLER_28_693 ();
 sg13g2_fill_1 FILLER_28_695 ();
 sg13g2_decap_4 FILLER_28_701 ();
 sg13g2_fill_1 FILLER_28_705 ();
 sg13g2_decap_4 FILLER_28_710 ();
 sg13g2_decap_4 FILLER_28_752 ();
 sg13g2_fill_1 FILLER_28_756 ();
 sg13g2_decap_8 FILLER_28_783 ();
 sg13g2_decap_8 FILLER_28_790 ();
 sg13g2_fill_2 FILLER_28_797 ();
 sg13g2_fill_1 FILLER_28_799 ();
 sg13g2_decap_8 FILLER_28_804 ();
 sg13g2_decap_4 FILLER_28_811 ();
 sg13g2_fill_2 FILLER_28_815 ();
 sg13g2_decap_4 FILLER_28_821 ();
 sg13g2_decap_8 FILLER_28_860 ();
 sg13g2_decap_4 FILLER_28_867 ();
 sg13g2_fill_2 FILLER_28_871 ();
 sg13g2_fill_1 FILLER_28_977 ();
 sg13g2_fill_2 FILLER_28_1004 ();
 sg13g2_fill_1 FILLER_28_1006 ();
 sg13g2_fill_2 FILLER_28_1033 ();
 sg13g2_fill_2 FILLER_28_1054 ();
 sg13g2_fill_2 FILLER_28_1070 ();
 sg13g2_fill_1 FILLER_28_1072 ();
 sg13g2_decap_4 FILLER_28_1079 ();
 sg13g2_fill_1 FILLER_28_1083 ();
 sg13g2_fill_1 FILLER_28_1088 ();
 sg13g2_fill_1 FILLER_28_1094 ();
 sg13g2_decap_8 FILLER_28_1099 ();
 sg13g2_fill_2 FILLER_28_1106 ();
 sg13g2_fill_1 FILLER_28_1114 ();
 sg13g2_fill_1 FILLER_28_1130 ();
 sg13g2_decap_8 FILLER_28_1144 ();
 sg13g2_fill_1 FILLER_28_1151 ();
 sg13g2_fill_2 FILLER_28_1158 ();
 sg13g2_fill_1 FILLER_28_1160 ();
 sg13g2_fill_2 FILLER_28_1175 ();
 sg13g2_fill_1 FILLER_28_1177 ();
 sg13g2_fill_1 FILLER_28_1183 ();
 sg13g2_decap_8 FILLER_28_1211 ();
 sg13g2_decap_4 FILLER_28_1279 ();
 sg13g2_fill_1 FILLER_28_1283 ();
 sg13g2_fill_1 FILLER_28_1310 ();
 sg13g2_decap_4 FILLER_28_1328 ();
 sg13g2_fill_1 FILLER_28_1394 ();
 sg13g2_decap_4 FILLER_28_1407 ();
 sg13g2_decap_8 FILLER_28_1423 ();
 sg13g2_decap_8 FILLER_28_1430 ();
 sg13g2_decap_8 FILLER_28_1453 ();
 sg13g2_fill_1 FILLER_28_1460 ();
 sg13g2_fill_2 FILLER_28_1496 ();
 sg13g2_fill_1 FILLER_28_1559 ();
 sg13g2_fill_2 FILLER_28_1568 ();
 sg13g2_fill_1 FILLER_28_1570 ();
 sg13g2_fill_2 FILLER_28_1640 ();
 sg13g2_fill_2 FILLER_28_1713 ();
 sg13g2_fill_1 FILLER_28_1715 ();
 sg13g2_decap_8 FILLER_28_1772 ();
 sg13g2_decap_4 FILLER_28_1779 ();
 sg13g2_fill_1 FILLER_28_1783 ();
 sg13g2_decap_4 FILLER_28_1789 ();
 sg13g2_decap_8 FILLER_28_1819 ();
 sg13g2_decap_8 FILLER_28_1861 ();
 sg13g2_decap_8 FILLER_28_1868 ();
 sg13g2_decap_8 FILLER_28_1879 ();
 sg13g2_decap_8 FILLER_28_1893 ();
 sg13g2_decap_4 FILLER_28_1900 ();
 sg13g2_fill_2 FILLER_28_1904 ();
 sg13g2_fill_2 FILLER_28_1929 ();
 sg13g2_fill_1 FILLER_28_1931 ();
 sg13g2_decap_4 FILLER_28_1943 ();
 sg13g2_fill_1 FILLER_28_1947 ();
 sg13g2_fill_1 FILLER_28_1951 ();
 sg13g2_decap_4 FILLER_28_1974 ();
 sg13g2_decap_4 FILLER_28_1982 ();
 sg13g2_fill_1 FILLER_28_1986 ();
 sg13g2_decap_4 FILLER_28_2006 ();
 sg13g2_fill_1 FILLER_28_2010 ();
 sg13g2_fill_2 FILLER_28_2051 ();
 sg13g2_fill_2 FILLER_28_2058 ();
 sg13g2_decap_8 FILLER_28_2091 ();
 sg13g2_fill_1 FILLER_28_2098 ();
 sg13g2_decap_8 FILLER_28_2103 ();
 sg13g2_decap_4 FILLER_28_2110 ();
 sg13g2_decap_8 FILLER_28_2144 ();
 sg13g2_fill_1 FILLER_28_2215 ();
 sg13g2_fill_2 FILLER_28_2264 ();
 sg13g2_fill_1 FILLER_28_2266 ();
 sg13g2_fill_1 FILLER_28_2285 ();
 sg13g2_fill_1 FILLER_28_2303 ();
 sg13g2_fill_2 FILLER_28_2334 ();
 sg13g2_fill_1 FILLER_28_2336 ();
 sg13g2_fill_1 FILLER_28_2372 ();
 sg13g2_decap_8 FILLER_28_2394 ();
 sg13g2_fill_2 FILLER_28_2401 ();
 sg13g2_fill_2 FILLER_28_2412 ();
 sg13g2_fill_2 FILLER_28_2418 ();
 sg13g2_fill_2 FILLER_28_2429 ();
 sg13g2_fill_1 FILLER_28_2431 ();
 sg13g2_decap_4 FILLER_28_2437 ();
 sg13g2_fill_2 FILLER_28_2449 ();
 sg13g2_fill_1 FILLER_28_2460 ();
 sg13g2_fill_2 FILLER_28_2474 ();
 sg13g2_fill_1 FILLER_28_2476 ();
 sg13g2_fill_2 FILLER_28_2495 ();
 sg13g2_fill_2 FILLER_28_2596 ();
 sg13g2_fill_1 FILLER_28_2598 ();
 sg13g2_fill_1 FILLER_28_2625 ();
 sg13g2_fill_2 FILLER_28_2652 ();
 sg13g2_decap_8 FILLER_28_2680 ();
 sg13g2_decap_8 FILLER_28_2687 ();
 sg13g2_fill_2 FILLER_28_2694 ();
 sg13g2_fill_1 FILLER_28_2696 ();
 sg13g2_decap_4 FILLER_28_2702 ();
 sg13g2_fill_2 FILLER_28_2711 ();
 sg13g2_fill_1 FILLER_28_2713 ();
 sg13g2_decap_8 FILLER_28_2718 ();
 sg13g2_decap_8 FILLER_28_2725 ();
 sg13g2_fill_1 FILLER_28_2732 ();
 sg13g2_fill_2 FILLER_28_2759 ();
 sg13g2_fill_1 FILLER_28_2761 ();
 sg13g2_fill_2 FILLER_28_2772 ();
 sg13g2_fill_1 FILLER_28_2774 ();
 sg13g2_decap_8 FILLER_28_2779 ();
 sg13g2_decap_8 FILLER_28_2786 ();
 sg13g2_decap_8 FILLER_28_2793 ();
 sg13g2_fill_2 FILLER_28_2800 ();
 sg13g2_decap_8 FILLER_28_2837 ();
 sg13g2_decap_8 FILLER_28_2844 ();
 sg13g2_decap_8 FILLER_28_2851 ();
 sg13g2_fill_2 FILLER_28_2858 ();
 sg13g2_fill_1 FILLER_28_2936 ();
 sg13g2_decap_4 FILLER_28_2977 ();
 sg13g2_fill_1 FILLER_28_2981 ();
 sg13g2_fill_1 FILLER_28_2987 ();
 sg13g2_fill_2 FILLER_28_2996 ();
 sg13g2_fill_2 FILLER_28_3012 ();
 sg13g2_fill_2 FILLER_28_3040 ();
 sg13g2_decap_8 FILLER_28_3055 ();
 sg13g2_decap_4 FILLER_28_3062 ();
 sg13g2_fill_1 FILLER_28_3066 ();
 sg13g2_decap_8 FILLER_28_3075 ();
 sg13g2_decap_4 FILLER_28_3082 ();
 sg13g2_fill_1 FILLER_28_3086 ();
 sg13g2_decap_8 FILLER_28_3091 ();
 sg13g2_decap_8 FILLER_28_3098 ();
 sg13g2_decap_8 FILLER_28_3105 ();
 sg13g2_fill_2 FILLER_28_3116 ();
 sg13g2_decap_8 FILLER_28_3127 ();
 sg13g2_fill_2 FILLER_28_3134 ();
 sg13g2_fill_2 FILLER_28_3165 ();
 sg13g2_decap_8 FILLER_28_3175 ();
 sg13g2_decap_8 FILLER_28_3182 ();
 sg13g2_decap_4 FILLER_28_3209 ();
 sg13g2_fill_1 FILLER_28_3213 ();
 sg13g2_fill_1 FILLER_28_3219 ();
 sg13g2_decap_8 FILLER_28_3228 ();
 sg13g2_decap_4 FILLER_28_3235 ();
 sg13g2_fill_2 FILLER_28_3251 ();
 sg13g2_fill_2 FILLER_28_3267 ();
 sg13g2_decap_8 FILLER_28_3281 ();
 sg13g2_fill_1 FILLER_28_3288 ();
 sg13g2_decap_4 FILLER_28_3339 ();
 sg13g2_fill_1 FILLER_28_3343 ();
 sg13g2_fill_2 FILLER_28_3353 ();
 sg13g2_fill_1 FILLER_28_3355 ();
 sg13g2_decap_8 FILLER_28_3369 ();
 sg13g2_decap_8 FILLER_28_3376 ();
 sg13g2_decap_8 FILLER_28_3383 ();
 sg13g2_decap_4 FILLER_28_3390 ();
 sg13g2_fill_2 FILLER_28_3394 ();
 sg13g2_decap_8 FILLER_28_3400 ();
 sg13g2_decap_8 FILLER_28_3407 ();
 sg13g2_fill_2 FILLER_28_3414 ();
 sg13g2_fill_1 FILLER_28_3435 ();
 sg13g2_fill_2 FILLER_28_3467 ();
 sg13g2_fill_1 FILLER_28_3480 ();
 sg13g2_decap_8 FILLER_28_3502 ();
 sg13g2_decap_8 FILLER_28_3509 ();
 sg13g2_fill_1 FILLER_28_3520 ();
 sg13g2_decap_8 FILLER_28_3538 ();
 sg13g2_decap_8 FILLER_28_3545 ();
 sg13g2_decap_8 FILLER_28_3552 ();
 sg13g2_fill_2 FILLER_28_3559 ();
 sg13g2_fill_1 FILLER_28_3561 ();
 sg13g2_decap_8 FILLER_28_3566 ();
 sg13g2_decap_8 FILLER_28_3573 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_4 FILLER_29_7 ();
 sg13g2_decap_4 FILLER_29_15 ();
 sg13g2_fill_2 FILLER_29_66 ();
 sg13g2_fill_1 FILLER_29_68 ();
 sg13g2_fill_1 FILLER_29_138 ();
 sg13g2_decap_4 FILLER_29_156 ();
 sg13g2_decap_8 FILLER_29_182 ();
 sg13g2_fill_1 FILLER_29_189 ();
 sg13g2_fill_1 FILLER_29_212 ();
 sg13g2_fill_1 FILLER_29_231 ();
 sg13g2_fill_2 FILLER_29_245 ();
 sg13g2_fill_1 FILLER_29_247 ();
 sg13g2_decap_4 FILLER_29_293 ();
 sg13g2_decap_8 FILLER_29_301 ();
 sg13g2_fill_2 FILLER_29_331 ();
 sg13g2_fill_2 FILLER_29_368 ();
 sg13g2_fill_2 FILLER_29_382 ();
 sg13g2_fill_1 FILLER_29_424 ();
 sg13g2_fill_2 FILLER_29_433 ();
 sg13g2_fill_2 FILLER_29_484 ();
 sg13g2_fill_1 FILLER_29_486 ();
 sg13g2_fill_2 FILLER_29_491 ();
 sg13g2_fill_1 FILLER_29_493 ();
 sg13g2_fill_2 FILLER_29_548 ();
 sg13g2_fill_1 FILLER_29_573 ();
 sg13g2_fill_2 FILLER_29_586 ();
 sg13g2_fill_1 FILLER_29_588 ();
 sg13g2_fill_1 FILLER_29_614 ();
 sg13g2_fill_1 FILLER_29_721 ();
 sg13g2_decap_8 FILLER_29_762 ();
 sg13g2_decap_4 FILLER_29_769 ();
 sg13g2_fill_2 FILLER_29_773 ();
 sg13g2_decap_4 FILLER_29_801 ();
 sg13g2_fill_1 FILLER_29_805 ();
 sg13g2_decap_4 FILLER_29_892 ();
 sg13g2_fill_2 FILLER_29_922 ();
 sg13g2_fill_1 FILLER_29_924 ();
 sg13g2_fill_2 FILLER_29_934 ();
 sg13g2_fill_1 FILLER_29_936 ();
 sg13g2_fill_2 FILLER_29_948 ();
 sg13g2_fill_2 FILLER_29_959 ();
 sg13g2_fill_1 FILLER_29_988 ();
 sg13g2_fill_1 FILLER_29_1003 ();
 sg13g2_decap_4 FILLER_29_1009 ();
 sg13g2_fill_1 FILLER_29_1017 ();
 sg13g2_fill_1 FILLER_29_1022 ();
 sg13g2_fill_1 FILLER_29_1037 ();
 sg13g2_fill_2 FILLER_29_1048 ();
 sg13g2_fill_1 FILLER_29_1050 ();
 sg13g2_fill_1 FILLER_29_1058 ();
 sg13g2_decap_8 FILLER_29_1064 ();
 sg13g2_fill_2 FILLER_29_1071 ();
 sg13g2_decap_8 FILLER_29_1077 ();
 sg13g2_decap_8 FILLER_29_1115 ();
 sg13g2_decap_8 FILLER_29_1122 ();
 sg13g2_fill_2 FILLER_29_1159 ();
 sg13g2_fill_1 FILLER_29_1161 ();
 sg13g2_decap_4 FILLER_29_1211 ();
 sg13g2_fill_1 FILLER_29_1215 ();
 sg13g2_fill_2 FILLER_29_1230 ();
 sg13g2_fill_1 FILLER_29_1232 ();
 sg13g2_fill_2 FILLER_29_1248 ();
 sg13g2_decap_4 FILLER_29_1284 ();
 sg13g2_fill_2 FILLER_29_1293 ();
 sg13g2_decap_8 FILLER_29_1299 ();
 sg13g2_fill_2 FILLER_29_1306 ();
 sg13g2_fill_1 FILLER_29_1320 ();
 sg13g2_decap_4 FILLER_29_1324 ();
 sg13g2_decap_4 FILLER_29_1333 ();
 sg13g2_fill_2 FILLER_29_1337 ();
 sg13g2_decap_8 FILLER_29_1369 ();
 sg13g2_fill_2 FILLER_29_1376 ();
 sg13g2_fill_1 FILLER_29_1378 ();
 sg13g2_fill_1 FILLER_29_1383 ();
 sg13g2_decap_8 FILLER_29_1389 ();
 sg13g2_decap_4 FILLER_29_1396 ();
 sg13g2_fill_2 FILLER_29_1400 ();
 sg13g2_decap_8 FILLER_29_1412 ();
 sg13g2_fill_2 FILLER_29_1419 ();
 sg13g2_decap_4 FILLER_29_1438 ();
 sg13g2_fill_1 FILLER_29_1442 ();
 sg13g2_fill_2 FILLER_29_1448 ();
 sg13g2_fill_1 FILLER_29_1467 ();
 sg13g2_fill_1 FILLER_29_1486 ();
 sg13g2_decap_4 FILLER_29_1492 ();
 sg13g2_fill_1 FILLER_29_1496 ();
 sg13g2_decap_8 FILLER_29_1516 ();
 sg13g2_decap_8 FILLER_29_1523 ();
 sg13g2_decap_4 FILLER_29_1530 ();
 sg13g2_decap_8 FILLER_29_1542 ();
 sg13g2_fill_2 FILLER_29_1566 ();
 sg13g2_fill_2 FILLER_29_1580 ();
 sg13g2_fill_1 FILLER_29_1626 ();
 sg13g2_fill_2 FILLER_29_1639 ();
 sg13g2_fill_1 FILLER_29_1690 ();
 sg13g2_decap_8 FILLER_29_1726 ();
 sg13g2_decap_8 FILLER_29_1733 ();
 sg13g2_decap_8 FILLER_29_1740 ();
 sg13g2_decap_4 FILLER_29_1747 ();
 sg13g2_fill_2 FILLER_29_1751 ();
 sg13g2_decap_8 FILLER_29_1795 ();
 sg13g2_fill_2 FILLER_29_1802 ();
 sg13g2_decap_4 FILLER_29_1808 ();
 sg13g2_decap_4 FILLER_29_1817 ();
 sg13g2_fill_1 FILLER_29_1821 ();
 sg13g2_decap_8 FILLER_29_1859 ();
 sg13g2_fill_1 FILLER_29_1866 ();
 sg13g2_decap_8 FILLER_29_1871 ();
 sg13g2_decap_4 FILLER_29_1878 ();
 sg13g2_decap_8 FILLER_29_1905 ();
 sg13g2_decap_4 FILLER_29_1912 ();
 sg13g2_fill_2 FILLER_29_1916 ();
 sg13g2_decap_8 FILLER_29_1923 ();
 sg13g2_decap_8 FILLER_29_1930 ();
 sg13g2_fill_1 FILLER_29_1947 ();
 sg13g2_fill_1 FILLER_29_1982 ();
 sg13g2_decap_8 FILLER_29_1988 ();
 sg13g2_fill_1 FILLER_29_2000 ();
 sg13g2_decap_8 FILLER_29_2009 ();
 sg13g2_decap_4 FILLER_29_2016 ();
 sg13g2_fill_2 FILLER_29_2030 ();
 sg13g2_fill_1 FILLER_29_2032 ();
 sg13g2_fill_2 FILLER_29_2042 ();
 sg13g2_fill_1 FILLER_29_2044 ();
 sg13g2_fill_1 FILLER_29_2073 ();
 sg13g2_decap_4 FILLER_29_2084 ();
 sg13g2_decap_8 FILLER_29_2114 ();
 sg13g2_fill_2 FILLER_29_2121 ();
 sg13g2_fill_1 FILLER_29_2123 ();
 sg13g2_decap_8 FILLER_29_2128 ();
 sg13g2_decap_8 FILLER_29_2135 ();
 sg13g2_fill_2 FILLER_29_2142 ();
 sg13g2_fill_1 FILLER_29_2144 ();
 sg13g2_fill_2 FILLER_29_2150 ();
 sg13g2_fill_1 FILLER_29_2152 ();
 sg13g2_decap_8 FILLER_29_2157 ();
 sg13g2_decap_4 FILLER_29_2164 ();
 sg13g2_fill_2 FILLER_29_2168 ();
 sg13g2_decap_8 FILLER_29_2174 ();
 sg13g2_decap_8 FILLER_29_2181 ();
 sg13g2_decap_8 FILLER_29_2188 ();
 sg13g2_decap_4 FILLER_29_2195 ();
 sg13g2_decap_8 FILLER_29_2220 ();
 sg13g2_decap_8 FILLER_29_2231 ();
 sg13g2_fill_1 FILLER_29_2317 ();
 sg13g2_fill_2 FILLER_29_2322 ();
 sg13g2_fill_1 FILLER_29_2324 ();
 sg13g2_fill_2 FILLER_29_2348 ();
 sg13g2_fill_1 FILLER_29_2364 ();
 sg13g2_decap_8 FILLER_29_2388 ();
 sg13g2_decap_8 FILLER_29_2395 ();
 sg13g2_fill_2 FILLER_29_2402 ();
 sg13g2_fill_1 FILLER_29_2487 ();
 sg13g2_fill_2 FILLER_29_2524 ();
 sg13g2_fill_2 FILLER_29_2530 ();
 sg13g2_fill_1 FILLER_29_2607 ();
 sg13g2_decap_4 FILLER_29_2613 ();
 sg13g2_fill_1 FILLER_29_2617 ();
 sg13g2_fill_2 FILLER_29_2631 ();
 sg13g2_fill_1 FILLER_29_2633 ();
 sg13g2_decap_4 FILLER_29_2643 ();
 sg13g2_fill_2 FILLER_29_2674 ();
 sg13g2_fill_1 FILLER_29_2698 ();
 sg13g2_fill_1 FILLER_29_2743 ();
 sg13g2_fill_2 FILLER_29_2748 ();
 sg13g2_fill_1 FILLER_29_2763 ();
 sg13g2_fill_1 FILLER_29_2790 ();
 sg13g2_fill_1 FILLER_29_2825 ();
 sg13g2_decap_8 FILLER_29_2860 ();
 sg13g2_fill_1 FILLER_29_2867 ();
 sg13g2_fill_1 FILLER_29_2873 ();
 sg13g2_fill_1 FILLER_29_2878 ();
 sg13g2_decap_8 FILLER_29_2897 ();
 sg13g2_fill_2 FILLER_29_2904 ();
 sg13g2_decap_8 FILLER_29_2926 ();
 sg13g2_fill_2 FILLER_29_2933 ();
 sg13g2_fill_1 FILLER_29_3004 ();
 sg13g2_fill_2 FILLER_29_3035 ();
 sg13g2_fill_1 FILLER_29_3037 ();
 sg13g2_fill_1 FILLER_29_3070 ();
 sg13g2_decap_4 FILLER_29_3097 ();
 sg13g2_fill_1 FILLER_29_3101 ();
 sg13g2_fill_2 FILLER_29_3107 ();
 sg13g2_fill_2 FILLER_29_3117 ();
 sg13g2_fill_2 FILLER_29_3133 ();
 sg13g2_decap_8 FILLER_29_3143 ();
 sg13g2_fill_2 FILLER_29_3150 ();
 sg13g2_fill_1 FILLER_29_3152 ();
 sg13g2_decap_8 FILLER_29_3158 ();
 sg13g2_decap_4 FILLER_29_3165 ();
 sg13g2_fill_1 FILLER_29_3169 ();
 sg13g2_decap_8 FILLER_29_3178 ();
 sg13g2_decap_4 FILLER_29_3185 ();
 sg13g2_fill_2 FILLER_29_3189 ();
 sg13g2_decap_8 FILLER_29_3196 ();
 sg13g2_fill_1 FILLER_29_3203 ();
 sg13g2_fill_1 FILLER_29_3246 ();
 sg13g2_decap_8 FILLER_29_3272 ();
 sg13g2_decap_8 FILLER_29_3279 ();
 sg13g2_fill_1 FILLER_29_3290 ();
 sg13g2_decap_4 FILLER_29_3319 ();
 sg13g2_fill_2 FILLER_29_3323 ();
 sg13g2_fill_2 FILLER_29_3337 ();
 sg13g2_fill_1 FILLER_29_3339 ();
 sg13g2_fill_1 FILLER_29_3376 ();
 sg13g2_fill_2 FILLER_29_3385 ();
 sg13g2_fill_1 FILLER_29_3387 ();
 sg13g2_decap_4 FILLER_29_3410 ();
 sg13g2_fill_2 FILLER_29_3414 ();
 sg13g2_decap_4 FILLER_29_3420 ();
 sg13g2_fill_2 FILLER_29_3424 ();
 sg13g2_decap_8 FILLER_29_3434 ();
 sg13g2_decap_8 FILLER_29_3441 ();
 sg13g2_decap_4 FILLER_29_3448 ();
 sg13g2_decap_8 FILLER_29_3461 ();
 sg13g2_decap_8 FILLER_29_3468 ();
 sg13g2_fill_1 FILLER_29_3475 ();
 sg13g2_fill_2 FILLER_29_3481 ();
 sg13g2_fill_1 FILLER_29_3483 ();
 sg13g2_fill_2 FILLER_29_3490 ();
 sg13g2_fill_2 FILLER_29_3500 ();
 sg13g2_fill_2 FILLER_29_3520 ();
 sg13g2_fill_2 FILLER_29_3527 ();
 sg13g2_fill_1 FILLER_29_3529 ();
 sg13g2_decap_4 FILLER_29_3539 ();
 sg13g2_fill_1 FILLER_29_3543 ();
 sg13g2_fill_1 FILLER_29_3579 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_7 ();
 sg13g2_fill_2 FILLER_30_27 ();
 sg13g2_decap_8 FILLER_30_58 ();
 sg13g2_fill_2 FILLER_30_65 ();
 sg13g2_fill_1 FILLER_30_67 ();
 sg13g2_fill_2 FILLER_30_82 ();
 sg13g2_fill_2 FILLER_30_110 ();
 sg13g2_decap_4 FILLER_30_122 ();
 sg13g2_fill_1 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_163 ();
 sg13g2_fill_2 FILLER_30_170 ();
 sg13g2_fill_2 FILLER_30_193 ();
 sg13g2_fill_2 FILLER_30_247 ();
 sg13g2_fill_1 FILLER_30_249 ();
 sg13g2_fill_2 FILLER_30_254 ();
 sg13g2_fill_1 FILLER_30_256 ();
 sg13g2_fill_2 FILLER_30_261 ();
 sg13g2_fill_1 FILLER_30_263 ();
 sg13g2_decap_8 FILLER_30_289 ();
 sg13g2_fill_1 FILLER_30_296 ();
 sg13g2_fill_2 FILLER_30_330 ();
 sg13g2_decap_8 FILLER_30_336 ();
 sg13g2_fill_2 FILLER_30_343 ();
 sg13g2_fill_1 FILLER_30_345 ();
 sg13g2_decap_4 FILLER_30_350 ();
 sg13g2_fill_2 FILLER_30_365 ();
 sg13g2_decap_8 FILLER_30_395 ();
 sg13g2_decap_8 FILLER_30_402 ();
 sg13g2_fill_2 FILLER_30_450 ();
 sg13g2_fill_1 FILLER_30_452 ();
 sg13g2_fill_1 FILLER_30_458 ();
 sg13g2_fill_2 FILLER_30_467 ();
 sg13g2_fill_2 FILLER_30_474 ();
 sg13g2_fill_1 FILLER_30_476 ();
 sg13g2_decap_8 FILLER_30_481 ();
 sg13g2_decap_8 FILLER_30_488 ();
 sg13g2_decap_4 FILLER_30_495 ();
 sg13g2_fill_2 FILLER_30_499 ();
 sg13g2_fill_2 FILLER_30_527 ();
 sg13g2_decap_4 FILLER_30_538 ();
 sg13g2_fill_1 FILLER_30_542 ();
 sg13g2_decap_8 FILLER_30_554 ();
 sg13g2_decap_4 FILLER_30_561 ();
 sg13g2_fill_1 FILLER_30_565 ();
 sg13g2_decap_8 FILLER_30_571 ();
 sg13g2_decap_4 FILLER_30_578 ();
 sg13g2_fill_1 FILLER_30_582 ();
 sg13g2_fill_2 FILLER_30_599 ();
 sg13g2_fill_1 FILLER_30_601 ();
 sg13g2_fill_2 FILLER_30_641 ();
 sg13g2_decap_8 FILLER_30_661 ();
 sg13g2_decap_8 FILLER_30_668 ();
 sg13g2_decap_4 FILLER_30_675 ();
 sg13g2_fill_2 FILLER_30_736 ();
 sg13g2_fill_2 FILLER_30_765 ();
 sg13g2_fill_1 FILLER_30_771 ();
 sg13g2_fill_1 FILLER_30_784 ();
 sg13g2_fill_2 FILLER_30_798 ();
 sg13g2_fill_1 FILLER_30_800 ();
 sg13g2_fill_1 FILLER_30_823 ();
 sg13g2_fill_1 FILLER_30_837 ();
 sg13g2_fill_2 FILLER_30_856 ();
 sg13g2_fill_2 FILLER_30_871 ();
 sg13g2_decap_8 FILLER_30_877 ();
 sg13g2_decap_8 FILLER_30_884 ();
 sg13g2_decap_8 FILLER_30_891 ();
 sg13g2_decap_4 FILLER_30_898 ();
 sg13g2_decap_8 FILLER_30_923 ();
 sg13g2_fill_2 FILLER_30_939 ();
 sg13g2_fill_2 FILLER_30_947 ();
 sg13g2_fill_1 FILLER_30_949 ();
 sg13g2_fill_1 FILLER_30_958 ();
 sg13g2_fill_2 FILLER_30_968 ();
 sg13g2_fill_1 FILLER_30_982 ();
 sg13g2_fill_2 FILLER_30_1038 ();
 sg13g2_decap_4 FILLER_30_1049 ();
 sg13g2_fill_1 FILLER_30_1053 ();
 sg13g2_decap_4 FILLER_30_1088 ();
 sg13g2_decap_8 FILLER_30_1125 ();
 sg13g2_fill_1 FILLER_30_1142 ();
 sg13g2_decap_8 FILLER_30_1172 ();
 sg13g2_decap_4 FILLER_30_1189 ();
 sg13g2_fill_2 FILLER_30_1193 ();
 sg13g2_fill_2 FILLER_30_1230 ();
 sg13g2_fill_2 FILLER_30_1248 ();
 sg13g2_decap_8 FILLER_30_1288 ();
 sg13g2_decap_8 FILLER_30_1295 ();
 sg13g2_decap_8 FILLER_30_1302 ();
 sg13g2_fill_2 FILLER_30_1309 ();
 sg13g2_fill_1 FILLER_30_1311 ();
 sg13g2_fill_2 FILLER_30_1316 ();
 sg13g2_decap_8 FILLER_30_1342 ();
 sg13g2_decap_8 FILLER_30_1353 ();
 sg13g2_decap_8 FILLER_30_1360 ();
 sg13g2_decap_4 FILLER_30_1367 ();
 sg13g2_decap_4 FILLER_30_1390 ();
 sg13g2_fill_2 FILLER_30_1394 ();
 sg13g2_fill_2 FILLER_30_1404 ();
 sg13g2_decap_4 FILLER_30_1416 ();
 sg13g2_fill_1 FILLER_30_1420 ();
 sg13g2_fill_2 FILLER_30_1429 ();
 sg13g2_fill_1 FILLER_30_1431 ();
 sg13g2_fill_1 FILLER_30_1469 ();
 sg13g2_decap_4 FILLER_30_1514 ();
 sg13g2_fill_2 FILLER_30_1548 ();
 sg13g2_fill_1 FILLER_30_1550 ();
 sg13g2_decap_4 FILLER_30_1556 ();
 sg13g2_fill_1 FILLER_30_1560 ();
 sg13g2_decap_4 FILLER_30_1571 ();
 sg13g2_fill_2 FILLER_30_1575 ();
 sg13g2_fill_2 FILLER_30_1602 ();
 sg13g2_fill_1 FILLER_30_1604 ();
 sg13g2_fill_1 FILLER_30_1623 ();
 sg13g2_fill_1 FILLER_30_1631 ();
 sg13g2_fill_2 FILLER_30_1669 ();
 sg13g2_decap_8 FILLER_30_1706 ();
 sg13g2_decap_8 FILLER_30_1713 ();
 sg13g2_fill_1 FILLER_30_1720 ();
 sg13g2_decap_4 FILLER_30_1731 ();
 sg13g2_fill_1 FILLER_30_1748 ();
 sg13g2_decap_8 FILLER_30_1753 ();
 sg13g2_decap_8 FILLER_30_1760 ();
 sg13g2_decap_4 FILLER_30_1767 ();
 sg13g2_decap_8 FILLER_30_1775 ();
 sg13g2_decap_4 FILLER_30_1796 ();
 sg13g2_fill_1 FILLER_30_1800 ();
 sg13g2_decap_4 FILLER_30_1841 ();
 sg13g2_fill_1 FILLER_30_1845 ();
 sg13g2_fill_2 FILLER_30_1854 ();
 sg13g2_fill_2 FILLER_30_1882 ();
 sg13g2_fill_1 FILLER_30_1887 ();
 sg13g2_fill_1 FILLER_30_1934 ();
 sg13g2_decap_8 FILLER_30_1940 ();
 sg13g2_decap_4 FILLER_30_1947 ();
 sg13g2_fill_2 FILLER_30_1951 ();
 sg13g2_decap_4 FILLER_30_1961 ();
 sg13g2_fill_2 FILLER_30_1979 ();
 sg13g2_decap_8 FILLER_30_2016 ();
 sg13g2_fill_2 FILLER_30_2023 ();
 sg13g2_fill_2 FILLER_30_2051 ();
 sg13g2_decap_4 FILLER_30_2105 ();
 sg13g2_decap_4 FILLER_30_2113 ();
 sg13g2_fill_1 FILLER_30_2117 ();
 sg13g2_decap_8 FILLER_30_2222 ();
 sg13g2_decap_8 FILLER_30_2229 ();
 sg13g2_decap_8 FILLER_30_2236 ();
 sg13g2_decap_8 FILLER_30_2243 ();
 sg13g2_decap_4 FILLER_30_2250 ();
 sg13g2_decap_8 FILLER_30_2267 ();
 sg13g2_decap_8 FILLER_30_2274 ();
 sg13g2_decap_8 FILLER_30_2281 ();
 sg13g2_decap_8 FILLER_30_2292 ();
 sg13g2_decap_4 FILLER_30_2299 ();
 sg13g2_fill_1 FILLER_30_2303 ();
 sg13g2_fill_1 FILLER_30_2330 ();
 sg13g2_decap_4 FILLER_30_2436 ();
 sg13g2_fill_2 FILLER_30_2440 ();
 sg13g2_decap_8 FILLER_30_2450 ();
 sg13g2_decap_8 FILLER_30_2457 ();
 sg13g2_fill_1 FILLER_30_2464 ();
 sg13g2_fill_1 FILLER_30_2470 ();
 sg13g2_decap_4 FILLER_30_2475 ();
 sg13g2_fill_1 FILLER_30_2479 ();
 sg13g2_decap_8 FILLER_30_2484 ();
 sg13g2_fill_1 FILLER_30_2503 ();
 sg13g2_fill_1 FILLER_30_2508 ();
 sg13g2_fill_2 FILLER_30_2518 ();
 sg13g2_fill_1 FILLER_30_2520 ();
 sg13g2_decap_8 FILLER_30_2547 ();
 sg13g2_decap_8 FILLER_30_2567 ();
 sg13g2_decap_8 FILLER_30_2574 ();
 sg13g2_fill_1 FILLER_30_2581 ();
 sg13g2_fill_1 FILLER_30_2603 ();
 sg13g2_decap_4 FILLER_30_2609 ();
 sg13g2_decap_4 FILLER_30_2673 ();
 sg13g2_fill_2 FILLER_30_2712 ();
 sg13g2_decap_8 FILLER_30_2803 ();
 sg13g2_decap_8 FILLER_30_2814 ();
 sg13g2_fill_2 FILLER_30_2821 ();
 sg13g2_decap_4 FILLER_30_2853 ();
 sg13g2_decap_8 FILLER_30_2902 ();
 sg13g2_decap_4 FILLER_30_2909 ();
 sg13g2_fill_1 FILLER_30_2920 ();
 sg13g2_decap_8 FILLER_30_2940 ();
 sg13g2_decap_8 FILLER_30_2947 ();
 sg13g2_decap_8 FILLER_30_2954 ();
 sg13g2_decap_4 FILLER_30_2961 ();
 sg13g2_fill_1 FILLER_30_2965 ();
 sg13g2_decap_8 FILLER_30_2970 ();
 sg13g2_fill_2 FILLER_30_2977 ();
 sg13g2_fill_1 FILLER_30_2979 ();
 sg13g2_decap_4 FILLER_30_2994 ();
 sg13g2_decap_8 FILLER_30_3003 ();
 sg13g2_decap_4 FILLER_30_3010 ();
 sg13g2_fill_2 FILLER_30_3014 ();
 sg13g2_decap_8 FILLER_30_3020 ();
 sg13g2_fill_2 FILLER_30_3027 ();
 sg13g2_fill_1 FILLER_30_3034 ();
 sg13g2_decap_8 FILLER_30_3058 ();
 sg13g2_decap_4 FILLER_30_3065 ();
 sg13g2_fill_1 FILLER_30_3069 ();
 sg13g2_fill_2 FILLER_30_3079 ();
 sg13g2_fill_1 FILLER_30_3081 ();
 sg13g2_fill_2 FILLER_30_3095 ();
 sg13g2_fill_1 FILLER_30_3097 ();
 sg13g2_decap_4 FILLER_30_3164 ();
 sg13g2_fill_2 FILLER_30_3199 ();
 sg13g2_decap_4 FILLER_30_3210 ();
 sg13g2_decap_4 FILLER_30_3219 ();
 sg13g2_decap_4 FILLER_30_3231 ();
 sg13g2_fill_1 FILLER_30_3235 ();
 sg13g2_fill_2 FILLER_30_3245 ();
 sg13g2_fill_1 FILLER_30_3247 ();
 sg13g2_decap_8 FILLER_30_3262 ();
 sg13g2_fill_2 FILLER_30_3269 ();
 sg13g2_fill_2 FILLER_30_3276 ();
 sg13g2_fill_1 FILLER_30_3278 ();
 sg13g2_fill_2 FILLER_30_3287 ();
 sg13g2_fill_1 FILLER_30_3289 ();
 sg13g2_fill_1 FILLER_30_3304 ();
 sg13g2_fill_2 FILLER_30_3314 ();
 sg13g2_fill_2 FILLER_30_3320 ();
 sg13g2_decap_8 FILLER_30_3330 ();
 sg13g2_decap_8 FILLER_30_3337 ();
 sg13g2_fill_2 FILLER_30_3344 ();
 sg13g2_fill_2 FILLER_30_3364 ();
 sg13g2_fill_1 FILLER_30_3366 ();
 sg13g2_fill_1 FILLER_30_3428 ();
 sg13g2_decap_4 FILLER_30_3455 ();
 sg13g2_fill_1 FILLER_30_3473 ();
 sg13g2_fill_1 FILLER_30_3479 ();
 sg13g2_decap_4 FILLER_30_3501 ();
 sg13g2_fill_2 FILLER_30_3531 ();
 sg13g2_fill_2 FILLER_30_3559 ();
 sg13g2_decap_4 FILLER_30_3574 ();
 sg13g2_fill_2 FILLER_30_3578 ();
 sg13g2_decap_4 FILLER_31_34 ();
 sg13g2_fill_1 FILLER_31_38 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_fill_2 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_83 ();
 sg13g2_fill_2 FILLER_31_90 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_fill_1 FILLER_31_147 ();
 sg13g2_fill_1 FILLER_31_152 ();
 sg13g2_fill_1 FILLER_31_163 ();
 sg13g2_fill_2 FILLER_31_194 ();
 sg13g2_fill_1 FILLER_31_196 ();
 sg13g2_fill_2 FILLER_31_205 ();
 sg13g2_fill_2 FILLER_31_211 ();
 sg13g2_fill_1 FILLER_31_218 ();
 sg13g2_decap_8 FILLER_31_223 ();
 sg13g2_decap_8 FILLER_31_264 ();
 sg13g2_decap_8 FILLER_31_271 ();
 sg13g2_decap_4 FILLER_31_278 ();
 sg13g2_fill_2 FILLER_31_282 ();
 sg13g2_fill_2 FILLER_31_309 ();
 sg13g2_decap_8 FILLER_31_315 ();
 sg13g2_fill_2 FILLER_31_322 ();
 sg13g2_fill_1 FILLER_31_324 ();
 sg13g2_fill_2 FILLER_31_368 ();
 sg13g2_fill_1 FILLER_31_396 ();
 sg13g2_fill_1 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_433 ();
 sg13g2_fill_1 FILLER_31_443 ();
 sg13g2_fill_2 FILLER_31_458 ();
 sg13g2_fill_1 FILLER_31_460 ();
 sg13g2_decap_8 FILLER_31_492 ();
 sg13g2_decap_4 FILLER_31_499 ();
 sg13g2_fill_2 FILLER_31_503 ();
 sg13g2_fill_2 FILLER_31_514 ();
 sg13g2_fill_1 FILLER_31_516 ();
 sg13g2_decap_4 FILLER_31_522 ();
 sg13g2_fill_1 FILLER_31_526 ();
 sg13g2_decap_4 FILLER_31_532 ();
 sg13g2_fill_1 FILLER_31_536 ();
 sg13g2_fill_2 FILLER_31_543 ();
 sg13g2_fill_1 FILLER_31_545 ();
 sg13g2_decap_4 FILLER_31_556 ();
 sg13g2_fill_1 FILLER_31_560 ();
 sg13g2_decap_8 FILLER_31_612 ();
 sg13g2_decap_8 FILLER_31_619 ();
 sg13g2_decap_4 FILLER_31_626 ();
 sg13g2_fill_2 FILLER_31_630 ();
 sg13g2_fill_2 FILLER_31_711 ();
 sg13g2_fill_1 FILLER_31_738 ();
 sg13g2_decap_4 FILLER_31_789 ();
 sg13g2_fill_1 FILLER_31_793 ();
 sg13g2_fill_2 FILLER_31_851 ();
 sg13g2_decap_4 FILLER_31_884 ();
 sg13g2_decap_8 FILLER_31_892 ();
 sg13g2_decap_8 FILLER_31_899 ();
 sg13g2_fill_2 FILLER_31_906 ();
 sg13g2_fill_1 FILLER_31_934 ();
 sg13g2_fill_2 FILLER_31_956 ();
 sg13g2_fill_1 FILLER_31_987 ();
 sg13g2_fill_2 FILLER_31_1018 ();
 sg13g2_fill_1 FILLER_31_1020 ();
 sg13g2_decap_4 FILLER_31_1035 ();
 sg13g2_fill_1 FILLER_31_1039 ();
 sg13g2_fill_2 FILLER_31_1160 ();
 sg13g2_decap_4 FILLER_31_1204 ();
 sg13g2_fill_2 FILLER_31_1208 ();
 sg13g2_decap_4 FILLER_31_1233 ();
 sg13g2_fill_2 FILLER_31_1250 ();
 sg13g2_fill_1 FILLER_31_1256 ();
 sg13g2_fill_1 FILLER_31_1270 ();
 sg13g2_fill_2 FILLER_31_1275 ();
 sg13g2_fill_1 FILLER_31_1277 ();
 sg13g2_decap_8 FILLER_31_1359 ();
 sg13g2_decap_8 FILLER_31_1366 ();
 sg13g2_fill_2 FILLER_31_1373 ();
 sg13g2_fill_1 FILLER_31_1382 ();
 sg13g2_decap_8 FILLER_31_1390 ();
 sg13g2_fill_1 FILLER_31_1397 ();
 sg13g2_decap_4 FILLER_31_1403 ();
 sg13g2_fill_2 FILLER_31_1407 ();
 sg13g2_fill_2 FILLER_31_1427 ();
 sg13g2_decap_8 FILLER_31_1455 ();
 sg13g2_fill_2 FILLER_31_1462 ();
 sg13g2_fill_1 FILLER_31_1472 ();
 sg13g2_fill_2 FILLER_31_1494 ();
 sg13g2_fill_1 FILLER_31_1496 ();
 sg13g2_decap_4 FILLER_31_1552 ();
 sg13g2_fill_1 FILLER_31_1582 ();
 sg13g2_fill_2 FILLER_31_1601 ();
 sg13g2_fill_2 FILLER_31_1629 ();
 sg13g2_fill_1 FILLER_31_1669 ();
 sg13g2_decap_8 FILLER_31_1696 ();
 sg13g2_decap_4 FILLER_31_1729 ();
 sg13g2_fill_2 FILLER_31_1733 ();
 sg13g2_fill_2 FILLER_31_1765 ();
 sg13g2_fill_1 FILLER_31_1767 ();
 sg13g2_fill_2 FILLER_31_1811 ();
 sg13g2_fill_1 FILLER_31_1813 ();
 sg13g2_fill_2 FILLER_31_1834 ();
 sg13g2_decap_8 FILLER_31_1862 ();
 sg13g2_decap_8 FILLER_31_1869 ();
 sg13g2_fill_2 FILLER_31_1876 ();
 sg13g2_fill_1 FILLER_31_1878 ();
 sg13g2_fill_1 FILLER_31_1897 ();
 sg13g2_fill_2 FILLER_31_1911 ();
 sg13g2_decap_8 FILLER_31_1918 ();
 sg13g2_fill_1 FILLER_31_1925 ();
 sg13g2_fill_2 FILLER_31_1959 ();
 sg13g2_fill_1 FILLER_31_1961 ();
 sg13g2_fill_2 FILLER_31_1977 ();
 sg13g2_decap_8 FILLER_31_1983 ();
 sg13g2_decap_8 FILLER_31_1990 ();
 sg13g2_fill_1 FILLER_31_1997 ();
 sg13g2_decap_4 FILLER_31_2017 ();
 sg13g2_decap_4 FILLER_31_2026 ();
 sg13g2_decap_8 FILLER_31_2058 ();
 sg13g2_fill_2 FILLER_31_2065 ();
 sg13g2_fill_2 FILLER_31_2127 ();
 sg13g2_fill_1 FILLER_31_2133 ();
 sg13g2_decap_8 FILLER_31_2138 ();
 sg13g2_decap_8 FILLER_31_2145 ();
 sg13g2_decap_8 FILLER_31_2152 ();
 sg13g2_decap_8 FILLER_31_2159 ();
 sg13g2_decap_4 FILLER_31_2166 ();
 sg13g2_fill_2 FILLER_31_2170 ();
 sg13g2_decap_8 FILLER_31_2176 ();
 sg13g2_fill_2 FILLER_31_2183 ();
 sg13g2_fill_1 FILLER_31_2185 ();
 sg13g2_decap_8 FILLER_31_2194 ();
 sg13g2_fill_2 FILLER_31_2201 ();
 sg13g2_fill_1 FILLER_31_2203 ();
 sg13g2_decap_4 FILLER_31_2256 ();
 sg13g2_fill_2 FILLER_31_2260 ();
 sg13g2_decap_8 FILLER_31_2294 ();
 sg13g2_decap_8 FILLER_31_2301 ();
 sg13g2_decap_4 FILLER_31_2330 ();
 sg13g2_fill_2 FILLER_31_2334 ();
 sg13g2_decap_8 FILLER_31_2357 ();
 sg13g2_decap_8 FILLER_31_2364 ();
 sg13g2_decap_4 FILLER_31_2375 ();
 sg13g2_fill_2 FILLER_31_2379 ();
 sg13g2_fill_2 FILLER_31_2399 ();
 sg13g2_fill_2 FILLER_31_2410 ();
 sg13g2_fill_1 FILLER_31_2554 ();
 sg13g2_fill_2 FILLER_31_2564 ();
 sg13g2_fill_1 FILLER_31_2566 ();
 sg13g2_fill_2 FILLER_31_2585 ();
 sg13g2_decap_8 FILLER_31_2626 ();
 sg13g2_decap_8 FILLER_31_2633 ();
 sg13g2_decap_8 FILLER_31_2640 ();
 sg13g2_fill_2 FILLER_31_2647 ();
 sg13g2_decap_4 FILLER_31_2653 ();
 sg13g2_fill_2 FILLER_31_2657 ();
 sg13g2_fill_1 FILLER_31_2672 ();
 sg13g2_fill_2 FILLER_31_2677 ();
 sg13g2_fill_1 FILLER_31_2683 ();
 sg13g2_decap_8 FILLER_31_2701 ();
 sg13g2_fill_2 FILLER_31_2708 ();
 sg13g2_decap_8 FILLER_31_2714 ();
 sg13g2_fill_2 FILLER_31_2721 ();
 sg13g2_fill_1 FILLER_31_2723 ();
 sg13g2_decap_8 FILLER_31_2736 ();
 sg13g2_fill_2 FILLER_31_2743 ();
 sg13g2_fill_1 FILLER_31_2785 ();
 sg13g2_decap_4 FILLER_31_2804 ();
 sg13g2_fill_2 FILLER_31_2808 ();
 sg13g2_fill_2 FILLER_31_2841 ();
 sg13g2_fill_1 FILLER_31_2843 ();
 sg13g2_decap_4 FILLER_31_2859 ();
 sg13g2_fill_1 FILLER_31_2863 ();
 sg13g2_decap_8 FILLER_31_2872 ();
 sg13g2_decap_8 FILLER_31_2879 ();
 sg13g2_decap_8 FILLER_31_2886 ();
 sg13g2_fill_2 FILLER_31_2893 ();
 sg13g2_fill_1 FILLER_31_2895 ();
 sg13g2_fill_2 FILLER_31_2901 ();
 sg13g2_fill_2 FILLER_31_2916 ();
 sg13g2_fill_1 FILLER_31_2918 ();
 sg13g2_fill_2 FILLER_31_2934 ();
 sg13g2_decap_4 FILLER_31_3019 ();
 sg13g2_fill_2 FILLER_31_3023 ();
 sg13g2_fill_2 FILLER_31_3051 ();
 sg13g2_fill_1 FILLER_31_3053 ();
 sg13g2_decap_4 FILLER_31_3085 ();
 sg13g2_fill_2 FILLER_31_3115 ();
 sg13g2_decap_4 FILLER_31_3121 ();
 sg13g2_fill_2 FILLER_31_3139 ();
 sg13g2_fill_1 FILLER_31_3141 ();
 sg13g2_decap_8 FILLER_31_3163 ();
 sg13g2_fill_1 FILLER_31_3179 ();
 sg13g2_fill_1 FILLER_31_3222 ();
 sg13g2_decap_4 FILLER_31_3232 ();
 sg13g2_fill_1 FILLER_31_3236 ();
 sg13g2_decap_4 FILLER_31_3263 ();
 sg13g2_fill_1 FILLER_31_3267 ();
 sg13g2_fill_2 FILLER_31_3303 ();
 sg13g2_decap_8 FILLER_31_3331 ();
 sg13g2_decap_4 FILLER_31_3368 ();
 sg13g2_fill_1 FILLER_31_3372 ();
 sg13g2_decap_4 FILLER_31_3386 ();
 sg13g2_fill_2 FILLER_31_3390 ();
 sg13g2_decap_8 FILLER_31_3410 ();
 sg13g2_decap_8 FILLER_31_3417 ();
 sg13g2_fill_2 FILLER_31_3424 ();
 sg13g2_fill_1 FILLER_31_3439 ();
 sg13g2_decap_8 FILLER_31_3444 ();
 sg13g2_decap_8 FILLER_31_3451 ();
 sg13g2_fill_2 FILLER_31_3473 ();
 sg13g2_fill_1 FILLER_31_3475 ();
 sg13g2_decap_8 FILLER_31_3489 ();
 sg13g2_fill_2 FILLER_31_3496 ();
 sg13g2_fill_1 FILLER_31_3498 ();
 sg13g2_decap_8 FILLER_31_3504 ();
 sg13g2_decap_8 FILLER_31_3511 ();
 sg13g2_decap_8 FILLER_31_3518 ();
 sg13g2_fill_2 FILLER_31_3525 ();
 sg13g2_fill_2 FILLER_31_3531 ();
 sg13g2_decap_8 FILLER_31_3559 ();
 sg13g2_decap_8 FILLER_31_3566 ();
 sg13g2_decap_8 FILLER_31_3573 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_7 ();
 sg13g2_fill_1 FILLER_32_9 ();
 sg13g2_fill_2 FILLER_32_55 ();
 sg13g2_fill_1 FILLER_32_57 ();
 sg13g2_fill_1 FILLER_32_67 ();
 sg13g2_fill_2 FILLER_32_80 ();
 sg13g2_fill_1 FILLER_32_82 ();
 sg13g2_fill_1 FILLER_32_115 ();
 sg13g2_fill_1 FILLER_32_129 ();
 sg13g2_fill_1 FILLER_32_139 ();
 sg13g2_fill_1 FILLER_32_150 ();
 sg13g2_fill_1 FILLER_32_200 ();
 sg13g2_fill_2 FILLER_32_206 ();
 sg13g2_fill_2 FILLER_32_234 ();
 sg13g2_decap_4 FILLER_32_293 ();
 sg13g2_decap_8 FILLER_32_302 ();
 sg13g2_fill_1 FILLER_32_340 ();
 sg13g2_fill_1 FILLER_32_346 ();
 sg13g2_decap_4 FILLER_32_356 ();
 sg13g2_fill_1 FILLER_32_360 ();
 sg13g2_fill_2 FILLER_32_368 ();
 sg13g2_fill_2 FILLER_32_403 ();
 sg13g2_fill_2 FILLER_32_460 ();
 sg13g2_fill_2 FILLER_32_475 ();
 sg13g2_decap_4 FILLER_32_513 ();
 sg13g2_fill_2 FILLER_32_517 ();
 sg13g2_decap_4 FILLER_32_530 ();
 sg13g2_fill_1 FILLER_32_534 ();
 sg13g2_decap_8 FILLER_32_539 ();
 sg13g2_fill_2 FILLER_32_546 ();
 sg13g2_fill_1 FILLER_32_548 ();
 sg13g2_fill_2 FILLER_32_559 ();
 sg13g2_fill_1 FILLER_32_561 ();
 sg13g2_fill_2 FILLER_32_571 ();
 sg13g2_fill_1 FILLER_32_573 ();
 sg13g2_decap_4 FILLER_32_587 ();
 sg13g2_fill_2 FILLER_32_596 ();
 sg13g2_fill_1 FILLER_32_598 ();
 sg13g2_decap_4 FILLER_32_603 ();
 sg13g2_fill_1 FILLER_32_607 ();
 sg13g2_fill_1 FILLER_32_648 ();
 sg13g2_decap_8 FILLER_32_654 ();
 sg13g2_decap_8 FILLER_32_661 ();
 sg13g2_decap_4 FILLER_32_668 ();
 sg13g2_fill_1 FILLER_32_721 ();
 sg13g2_fill_1 FILLER_32_735 ();
 sg13g2_fill_2 FILLER_32_745 ();
 sg13g2_fill_1 FILLER_32_747 ();
 sg13g2_decap_8 FILLER_32_798 ();
 sg13g2_fill_2 FILLER_32_805 ();
 sg13g2_fill_1 FILLER_32_807 ();
 sg13g2_fill_1 FILLER_32_812 ();
 sg13g2_fill_2 FILLER_32_847 ();
 sg13g2_fill_1 FILLER_32_849 ();
 sg13g2_fill_2 FILLER_32_855 ();
 sg13g2_fill_2 FILLER_32_865 ();
 sg13g2_fill_2 FILLER_32_876 ();
 sg13g2_decap_8 FILLER_32_904 ();
 sg13g2_decap_8 FILLER_32_911 ();
 sg13g2_fill_1 FILLER_32_918 ();
 sg13g2_fill_2 FILLER_32_951 ();
 sg13g2_fill_2 FILLER_32_1008 ();
 sg13g2_fill_2 FILLER_32_1019 ();
 sg13g2_decap_4 FILLER_32_1042 ();
 sg13g2_fill_2 FILLER_32_1046 ();
 sg13g2_fill_2 FILLER_32_1052 ();
 sg13g2_decap_4 FILLER_32_1058 ();
 sg13g2_fill_2 FILLER_32_1071 ();
 sg13g2_fill_1 FILLER_32_1073 ();
 sg13g2_decap_8 FILLER_32_1146 ();
 sg13g2_decap_4 FILLER_32_1153 ();
 sg13g2_decap_8 FILLER_32_1183 ();
 sg13g2_decap_8 FILLER_32_1190 ();
 sg13g2_fill_2 FILLER_32_1197 ();
 sg13g2_decap_4 FILLER_32_1225 ();
 sg13g2_fill_1 FILLER_32_1237 ();
 sg13g2_fill_2 FILLER_32_1253 ();
 sg13g2_fill_1 FILLER_32_1255 ();
 sg13g2_decap_8 FILLER_32_1287 ();
 sg13g2_fill_2 FILLER_32_1294 ();
 sg13g2_decap_4 FILLER_32_1306 ();
 sg13g2_fill_2 FILLER_32_1315 ();
 sg13g2_fill_1 FILLER_32_1325 ();
 sg13g2_decap_8 FILLER_32_1357 ();
 sg13g2_fill_2 FILLER_32_1398 ();
 sg13g2_decap_8 FILLER_32_1408 ();
 sg13g2_fill_2 FILLER_32_1415 ();
 sg13g2_fill_1 FILLER_32_1417 ();
 sg13g2_fill_2 FILLER_32_1428 ();
 sg13g2_fill_1 FILLER_32_1430 ();
 sg13g2_decap_8 FILLER_32_1461 ();
 sg13g2_fill_2 FILLER_32_1468 ();
 sg13g2_fill_1 FILLER_32_1510 ();
 sg13g2_fill_1 FILLER_32_1520 ();
 sg13g2_fill_1 FILLER_32_1534 ();
 sg13g2_fill_1 FILLER_32_1543 ();
 sg13g2_decap_4 FILLER_32_1549 ();
 sg13g2_fill_2 FILLER_32_1553 ();
 sg13g2_fill_1 FILLER_32_1560 ();
 sg13g2_fill_2 FILLER_32_1614 ();
 sg13g2_fill_1 FILLER_32_1642 ();
 sg13g2_fill_2 FILLER_32_1678 ();
 sg13g2_decap_8 FILLER_32_1706 ();
 sg13g2_fill_1 FILLER_32_1713 ();
 sg13g2_decap_8 FILLER_32_1722 ();
 sg13g2_decap_4 FILLER_32_1729 ();
 sg13g2_fill_2 FILLER_32_1741 ();
 sg13g2_decap_8 FILLER_32_1748 ();
 sg13g2_decap_8 FILLER_32_1755 ();
 sg13g2_fill_2 FILLER_32_1762 ();
 sg13g2_fill_1 FILLER_32_1764 ();
 sg13g2_fill_2 FILLER_32_1782 ();
 sg13g2_decap_8 FILLER_32_1789 ();
 sg13g2_decap_8 FILLER_32_1796 ();
 sg13g2_decap_8 FILLER_32_1803 ();
 sg13g2_fill_2 FILLER_32_1810 ();
 sg13g2_fill_1 FILLER_32_1812 ();
 sg13g2_decap_4 FILLER_32_1817 ();
 sg13g2_fill_1 FILLER_32_1821 ();
 sg13g2_fill_1 FILLER_32_1830 ();
 sg13g2_decap_4 FILLER_32_1836 ();
 sg13g2_fill_2 FILLER_32_1840 ();
 sg13g2_fill_2 FILLER_32_1851 ();
 sg13g2_fill_1 FILLER_32_1853 ();
 sg13g2_fill_2 FILLER_32_1892 ();
 sg13g2_decap_4 FILLER_32_1913 ();
 sg13g2_fill_1 FILLER_32_1917 ();
 sg13g2_decap_8 FILLER_32_1922 ();
 sg13g2_decap_8 FILLER_32_1929 ();
 sg13g2_fill_2 FILLER_32_1940 ();
 sg13g2_fill_2 FILLER_32_1946 ();
 sg13g2_decap_4 FILLER_32_1953 ();
 sg13g2_fill_2 FILLER_32_1957 ();
 sg13g2_decap_4 FILLER_32_2013 ();
 sg13g2_fill_1 FILLER_32_2017 ();
 sg13g2_decap_4 FILLER_32_2028 ();
 sg13g2_fill_1 FILLER_32_2041 ();
 sg13g2_decap_4 FILLER_32_2106 ();
 sg13g2_fill_2 FILLER_32_2110 ();
 sg13g2_fill_2 FILLER_32_2121 ();
 sg13g2_fill_2 FILLER_32_2127 ();
 sg13g2_decap_8 FILLER_32_2134 ();
 sg13g2_fill_1 FILLER_32_2141 ();
 sg13g2_decap_4 FILLER_32_2172 ();
 sg13g2_fill_1 FILLER_32_2176 ();
 sg13g2_decap_8 FILLER_32_2201 ();
 sg13g2_decap_4 FILLER_32_2208 ();
 sg13g2_fill_1 FILLER_32_2224 ();
 sg13g2_decap_4 FILLER_32_2230 ();
 sg13g2_fill_2 FILLER_32_2234 ();
 sg13g2_decap_4 FILLER_32_2240 ();
 sg13g2_fill_2 FILLER_32_2244 ();
 sg13g2_decap_8 FILLER_32_2258 ();
 sg13g2_decap_8 FILLER_32_2265 ();
 sg13g2_decap_8 FILLER_32_2272 ();
 sg13g2_decap_4 FILLER_32_2283 ();
 sg13g2_fill_1 FILLER_32_2287 ();
 sg13g2_decap_4 FILLER_32_2320 ();
 sg13g2_fill_1 FILLER_32_2324 ();
 sg13g2_decap_8 FILLER_32_2355 ();
 sg13g2_decap_8 FILLER_32_2362 ();
 sg13g2_fill_2 FILLER_32_2369 ();
 sg13g2_fill_2 FILLER_32_2398 ();
 sg13g2_fill_1 FILLER_32_2400 ();
 sg13g2_fill_2 FILLER_32_2414 ();
 sg13g2_fill_1 FILLER_32_2416 ();
 sg13g2_decap_8 FILLER_32_2422 ();
 sg13g2_decap_4 FILLER_32_2429 ();
 sg13g2_fill_1 FILLER_32_2433 ();
 sg13g2_decap_4 FILLER_32_2438 ();
 sg13g2_fill_2 FILLER_32_2447 ();
 sg13g2_fill_1 FILLER_32_2449 ();
 sg13g2_decap_4 FILLER_32_2463 ();
 sg13g2_fill_2 FILLER_32_2467 ();
 sg13g2_fill_1 FILLER_32_2516 ();
 sg13g2_decap_8 FILLER_32_2531 ();
 sg13g2_fill_2 FILLER_32_2564 ();
 sg13g2_fill_1 FILLER_32_2566 ();
 sg13g2_fill_2 FILLER_32_2602 ();
 sg13g2_decap_8 FILLER_32_2636 ();
 sg13g2_fill_2 FILLER_32_2643 ();
 sg13g2_decap_4 FILLER_32_2658 ();
 sg13g2_fill_1 FILLER_32_2662 ();
 sg13g2_fill_2 FILLER_32_2694 ();
 sg13g2_decap_4 FILLER_32_2774 ();
 sg13g2_fill_2 FILLER_32_2778 ();
 sg13g2_decap_4 FILLER_32_2804 ();
 sg13g2_fill_1 FILLER_32_2808 ();
 sg13g2_decap_4 FILLER_32_2819 ();
 sg13g2_decap_8 FILLER_32_2831 ();
 sg13g2_decap_8 FILLER_32_2838 ();
 sg13g2_fill_2 FILLER_32_2845 ();
 sg13g2_fill_2 FILLER_32_2856 ();
 sg13g2_fill_1 FILLER_32_2858 ();
 sg13g2_fill_2 FILLER_32_2864 ();
 sg13g2_fill_2 FILLER_32_2870 ();
 sg13g2_fill_1 FILLER_32_2890 ();
 sg13g2_fill_2 FILLER_32_2896 ();
 sg13g2_decap_8 FILLER_32_2916 ();
 sg13g2_fill_1 FILLER_32_2923 ();
 sg13g2_decap_4 FILLER_32_2933 ();
 sg13g2_fill_2 FILLER_32_2950 ();
 sg13g2_fill_1 FILLER_32_2952 ();
 sg13g2_fill_1 FILLER_32_2962 ();
 sg13g2_decap_8 FILLER_32_2968 ();
 sg13g2_decap_8 FILLER_32_2979 ();
 sg13g2_decap_8 FILLER_32_2986 ();
 sg13g2_decap_4 FILLER_32_2993 ();
 sg13g2_fill_1 FILLER_32_2997 ();
 sg13g2_decap_4 FILLER_32_3022 ();
 sg13g2_fill_2 FILLER_32_3026 ();
 sg13g2_decap_8 FILLER_32_3041 ();
 sg13g2_decap_4 FILLER_32_3048 ();
 sg13g2_fill_1 FILLER_32_3069 ();
 sg13g2_fill_1 FILLER_32_3074 ();
 sg13g2_fill_2 FILLER_32_3084 ();
 sg13g2_fill_1 FILLER_32_3086 ();
 sg13g2_fill_2 FILLER_32_3096 ();
 sg13g2_decap_4 FILLER_32_3142 ();
 sg13g2_decap_8 FILLER_32_3157 ();
 sg13g2_decap_8 FILLER_32_3164 ();
 sg13g2_fill_2 FILLER_32_3171 ();
 sg13g2_fill_1 FILLER_32_3183 ();
 sg13g2_decap_4 FILLER_32_3244 ();
 sg13g2_decap_8 FILLER_32_3252 ();
 sg13g2_decap_4 FILLER_32_3259 ();
 sg13g2_decap_4 FILLER_32_3276 ();
 sg13g2_fill_1 FILLER_32_3280 ();
 sg13g2_decap_4 FILLER_32_3286 ();
 sg13g2_fill_1 FILLER_32_3290 ();
 sg13g2_decap_8 FILLER_32_3317 ();
 sg13g2_decap_8 FILLER_32_3332 ();
 sg13g2_decap_8 FILLER_32_3339 ();
 sg13g2_fill_1 FILLER_32_3346 ();
 sg13g2_fill_1 FILLER_32_3355 ();
 sg13g2_decap_8 FILLER_32_3374 ();
 sg13g2_decap_8 FILLER_32_3381 ();
 sg13g2_fill_2 FILLER_32_3388 ();
 sg13g2_fill_1 FILLER_32_3390 ();
 sg13g2_fill_1 FILLER_32_3399 ();
 sg13g2_decap_8 FILLER_32_3404 ();
 sg13g2_decap_8 FILLER_32_3424 ();
 sg13g2_decap_4 FILLER_32_3431 ();
 sg13g2_fill_1 FILLER_32_3435 ();
 sg13g2_decap_8 FILLER_32_3449 ();
 sg13g2_decap_8 FILLER_32_3456 ();
 sg13g2_fill_2 FILLER_32_3463 ();
 sg13g2_fill_1 FILLER_32_3465 ();
 sg13g2_decap_4 FILLER_32_3492 ();
 sg13g2_fill_1 FILLER_32_3522 ();
 sg13g2_decap_8 FILLER_32_3554 ();
 sg13g2_decap_8 FILLER_32_3561 ();
 sg13g2_decap_8 FILLER_32_3568 ();
 sg13g2_decap_4 FILLER_32_3575 ();
 sg13g2_fill_1 FILLER_32_3579 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_4 FILLER_33_7 ();
 sg13g2_fill_1 FILLER_33_15 ();
 sg13g2_decap_4 FILLER_33_38 ();
 sg13g2_fill_2 FILLER_33_42 ();
 sg13g2_fill_2 FILLER_33_48 ();
 sg13g2_fill_1 FILLER_33_50 ();
 sg13g2_fill_2 FILLER_33_60 ();
 sg13g2_fill_2 FILLER_33_70 ();
 sg13g2_fill_1 FILLER_33_72 ();
 sg13g2_fill_1 FILLER_33_90 ();
 sg13g2_fill_1 FILLER_33_113 ();
 sg13g2_fill_2 FILLER_33_183 ();
 sg13g2_fill_1 FILLER_33_185 ();
 sg13g2_fill_1 FILLER_33_195 ();
 sg13g2_fill_2 FILLER_33_259 ();
 sg13g2_fill_1 FILLER_33_310 ();
 sg13g2_fill_1 FILLER_33_348 ();
 sg13g2_fill_2 FILLER_33_366 ();
 sg13g2_decap_4 FILLER_33_386 ();
 sg13g2_fill_2 FILLER_33_390 ();
 sg13g2_fill_1 FILLER_33_424 ();
 sg13g2_fill_1 FILLER_33_469 ();
 sg13g2_decap_8 FILLER_33_507 ();
 sg13g2_fill_1 FILLER_33_514 ();
 sg13g2_decap_8 FILLER_33_541 ();
 sg13g2_fill_2 FILLER_33_548 ();
 sg13g2_decap_8 FILLER_33_558 ();
 sg13g2_fill_1 FILLER_33_663 ();
 sg13g2_fill_1 FILLER_33_699 ();
 sg13g2_fill_2 FILLER_33_714 ();
 sg13g2_fill_2 FILLER_33_729 ();
 sg13g2_fill_2 FILLER_33_746 ();
 sg13g2_fill_2 FILLER_33_765 ();
 sg13g2_decap_4 FILLER_33_772 ();
 sg13g2_fill_2 FILLER_33_795 ();
 sg13g2_fill_2 FILLER_33_812 ();
 sg13g2_decap_8 FILLER_33_819 ();
 sg13g2_decap_4 FILLER_33_826 ();
 sg13g2_decap_4 FILLER_33_845 ();
 sg13g2_fill_2 FILLER_33_849 ();
 sg13g2_decap_8 FILLER_33_892 ();
 sg13g2_decap_4 FILLER_33_899 ();
 sg13g2_fill_1 FILLER_33_903 ();
 sg13g2_fill_1 FILLER_33_939 ();
 sg13g2_decap_4 FILLER_33_973 ();
 sg13g2_fill_1 FILLER_33_977 ();
 sg13g2_decap_8 FILLER_33_1008 ();
 sg13g2_fill_1 FILLER_33_1015 ();
 sg13g2_fill_2 FILLER_33_1094 ();
 sg13g2_fill_1 FILLER_33_1096 ();
 sg13g2_fill_2 FILLER_33_1125 ();
 sg13g2_fill_2 FILLER_33_1162 ();
 sg13g2_fill_1 FILLER_33_1164 ();
 sg13g2_decap_4 FILLER_33_1200 ();
 sg13g2_fill_2 FILLER_33_1217 ();
 sg13g2_fill_1 FILLER_33_1219 ();
 sg13g2_decap_4 FILLER_33_1233 ();
 sg13g2_decap_4 FILLER_33_1242 ();
 sg13g2_fill_1 FILLER_33_1246 ();
 sg13g2_fill_1 FILLER_33_1251 ();
 sg13g2_decap_8 FILLER_33_1260 ();
 sg13g2_decap_8 FILLER_33_1267 ();
 sg13g2_decap_4 FILLER_33_1274 ();
 sg13g2_fill_1 FILLER_33_1323 ();
 sg13g2_fill_1 FILLER_33_1350 ();
 sg13g2_fill_1 FILLER_33_1408 ();
 sg13g2_decap_8 FILLER_33_1435 ();
 sg13g2_fill_2 FILLER_33_1442 ();
 sg13g2_fill_2 FILLER_33_1449 ();
 sg13g2_fill_1 FILLER_33_1451 ();
 sg13g2_fill_1 FILLER_33_1456 ();
 sg13g2_fill_2 FILLER_33_1483 ();
 sg13g2_fill_2 FILLER_33_1520 ();
 sg13g2_fill_2 FILLER_33_1548 ();
 sg13g2_fill_2 FILLER_33_1558 ();
 sg13g2_fill_1 FILLER_33_1583 ();
 sg13g2_fill_1 FILLER_33_1595 ();
 sg13g2_fill_2 FILLER_33_1605 ();
 sg13g2_fill_2 FILLER_33_1626 ();
 sg13g2_fill_1 FILLER_33_1642 ();
 sg13g2_fill_2 FILLER_33_1688 ();
 sg13g2_fill_1 FILLER_33_1690 ();
 sg13g2_decap_8 FILLER_33_1695 ();
 sg13g2_fill_1 FILLER_33_1702 ();
 sg13g2_decap_4 FILLER_33_1729 ();
 sg13g2_fill_1 FILLER_33_1733 ();
 sg13g2_decap_8 FILLER_33_1760 ();
 sg13g2_fill_1 FILLER_33_1767 ();
 sg13g2_fill_1 FILLER_33_1787 ();
 sg13g2_decap_8 FILLER_33_1796 ();
 sg13g2_fill_2 FILLER_33_1803 ();
 sg13g2_fill_2 FILLER_33_1813 ();
 sg13g2_decap_4 FILLER_33_1820 ();
 sg13g2_fill_1 FILLER_33_1824 ();
 sg13g2_fill_2 FILLER_33_1830 ();
 sg13g2_fill_1 FILLER_33_1832 ();
 sg13g2_fill_1 FILLER_33_1837 ();
 sg13g2_fill_2 FILLER_33_1853 ();
 sg13g2_fill_1 FILLER_33_1855 ();
 sg13g2_fill_2 FILLER_33_1862 ();
 sg13g2_fill_1 FILLER_33_1890 ();
 sg13g2_decap_8 FILLER_33_1896 ();
 sg13g2_fill_1 FILLER_33_1903 ();
 sg13g2_decap_4 FILLER_33_1921 ();
 sg13g2_fill_2 FILLER_33_1925 ();
 sg13g2_decap_8 FILLER_33_1931 ();
 sg13g2_decap_4 FILLER_33_1938 ();
 sg13g2_fill_1 FILLER_33_1942 ();
 sg13g2_decap_8 FILLER_33_1951 ();
 sg13g2_decap_4 FILLER_33_1958 ();
 sg13g2_fill_1 FILLER_33_1962 ();
 sg13g2_fill_1 FILLER_33_1993 ();
 sg13g2_decap_8 FILLER_33_2009 ();
 sg13g2_fill_1 FILLER_33_2016 ();
 sg13g2_fill_1 FILLER_33_2052 ();
 sg13g2_decap_4 FILLER_33_2057 ();
 sg13g2_decap_8 FILLER_33_2067 ();
 sg13g2_fill_2 FILLER_33_2074 ();
 sg13g2_fill_1 FILLER_33_2076 ();
 sg13g2_decap_8 FILLER_33_2081 ();
 sg13g2_decap_4 FILLER_33_2088 ();
 sg13g2_fill_2 FILLER_33_2114 ();
 sg13g2_fill_1 FILLER_33_2116 ();
 sg13g2_fill_1 FILLER_33_2125 ();
 sg13g2_decap_8 FILLER_33_2139 ();
 sg13g2_decap_4 FILLER_33_2146 ();
 sg13g2_fill_2 FILLER_33_2168 ();
 sg13g2_fill_1 FILLER_33_2170 ();
 sg13g2_decap_8 FILLER_33_2200 ();
 sg13g2_decap_8 FILLER_33_2207 ();
 sg13g2_fill_2 FILLER_33_2214 ();
 sg13g2_fill_1 FILLER_33_2216 ();
 sg13g2_fill_1 FILLER_33_2242 ();
 sg13g2_fill_1 FILLER_33_2269 ();
 sg13g2_decap_4 FILLER_33_2301 ();
 sg13g2_decap_8 FILLER_33_2309 ();
 sg13g2_decap_8 FILLER_33_2316 ();
 sg13g2_decap_8 FILLER_33_2323 ();
 sg13g2_decap_8 FILLER_33_2330 ();
 sg13g2_fill_1 FILLER_33_2363 ();
 sg13g2_fill_1 FILLER_33_2421 ();
 sg13g2_fill_2 FILLER_33_2448 ();
 sg13g2_fill_1 FILLER_33_2450 ();
 sg13g2_decap_4 FILLER_33_2460 ();
 sg13g2_fill_2 FILLER_33_2464 ();
 sg13g2_decap_8 FILLER_33_2492 ();
 sg13g2_fill_1 FILLER_33_2499 ();
 sg13g2_fill_1 FILLER_33_2504 ();
 sg13g2_decap_8 FILLER_33_2508 ();
 sg13g2_fill_1 FILLER_33_2515 ();
 sg13g2_fill_1 FILLER_33_2523 ();
 sg13g2_decap_8 FILLER_33_2528 ();
 sg13g2_decap_8 FILLER_33_2535 ();
 sg13g2_decap_8 FILLER_33_2542 ();
 sg13g2_fill_1 FILLER_33_2549 ();
 sg13g2_decap_8 FILLER_33_2554 ();
 sg13g2_decap_8 FILLER_33_2561 ();
 sg13g2_fill_1 FILLER_33_2568 ();
 sg13g2_decap_4 FILLER_33_2604 ();
 sg13g2_fill_1 FILLER_33_2608 ();
 sg13g2_fill_2 FILLER_33_2618 ();
 sg13g2_fill_1 FILLER_33_2620 ();
 sg13g2_decap_8 FILLER_33_2625 ();
 sg13g2_fill_2 FILLER_33_2632 ();
 sg13g2_decap_8 FILLER_33_2691 ();
 sg13g2_decap_8 FILLER_33_2698 ();
 sg13g2_fill_2 FILLER_33_2705 ();
 sg13g2_decap_4 FILLER_33_2711 ();
 sg13g2_fill_1 FILLER_33_2715 ();
 sg13g2_decap_8 FILLER_33_2720 ();
 sg13g2_decap_4 FILLER_33_2727 ();
 sg13g2_fill_1 FILLER_33_2731 ();
 sg13g2_fill_1 FILLER_33_2741 ();
 sg13g2_fill_2 FILLER_33_2759 ();
 sg13g2_fill_2 FILLER_33_2770 ();
 sg13g2_fill_1 FILLER_33_2772 ();
 sg13g2_fill_2 FILLER_33_2813 ();
 sg13g2_fill_1 FILLER_33_2823 ();
 sg13g2_decap_8 FILLER_33_2841 ();
 sg13g2_fill_2 FILLER_33_2848 ();
 sg13g2_fill_2 FILLER_33_2868 ();
 sg13g2_fill_2 FILLER_33_2875 ();
 sg13g2_decap_8 FILLER_33_2889 ();
 sg13g2_fill_1 FILLER_33_2900 ();
 sg13g2_fill_2 FILLER_33_2920 ();
 sg13g2_fill_1 FILLER_33_2922 ();
 sg13g2_fill_2 FILLER_33_2940 ();
 sg13g2_fill_2 FILLER_33_2968 ();
 sg13g2_fill_1 FILLER_33_2970 ();
 sg13g2_decap_8 FILLER_33_2975 ();
 sg13g2_decap_8 FILLER_33_2995 ();
 sg13g2_fill_2 FILLER_33_3037 ();
 sg13g2_fill_1 FILLER_33_3039 ();
 sg13g2_decap_8 FILLER_33_3046 ();
 sg13g2_decap_8 FILLER_33_3053 ();
 sg13g2_fill_1 FILLER_33_3060 ();
 sg13g2_decap_4 FILLER_33_3069 ();
 sg13g2_fill_1 FILLER_33_3073 ();
 sg13g2_decap_4 FILLER_33_3121 ();
 sg13g2_fill_2 FILLER_33_3125 ();
 sg13g2_decap_8 FILLER_33_3131 ();
 sg13g2_fill_1 FILLER_33_3138 ();
 sg13g2_decap_8 FILLER_33_3157 ();
 sg13g2_fill_1 FILLER_33_3174 ();
 sg13g2_decap_4 FILLER_33_3190 ();
 sg13g2_fill_2 FILLER_33_3194 ();
 sg13g2_decap_8 FILLER_33_3201 ();
 sg13g2_fill_2 FILLER_33_3208 ();
 sg13g2_fill_1 FILLER_33_3210 ();
 sg13g2_fill_1 FILLER_33_3224 ();
 sg13g2_decap_8 FILLER_33_3233 ();
 sg13g2_decap_4 FILLER_33_3240 ();
 sg13g2_fill_2 FILLER_33_3244 ();
 sg13g2_decap_4 FILLER_33_3293 ();
 sg13g2_fill_1 FILLER_33_3297 ();
 sg13g2_fill_2 FILLER_33_3313 ();
 sg13g2_fill_1 FILLER_33_3366 ();
 sg13g2_fill_2 FILLER_33_3376 ();
 sg13g2_fill_1 FILLER_33_3378 ();
 sg13g2_fill_2 FILLER_33_3400 ();
 sg13g2_fill_1 FILLER_33_3402 ();
 sg13g2_fill_2 FILLER_33_3429 ();
 sg13g2_fill_1 FILLER_33_3431 ();
 sg13g2_fill_2 FILLER_33_3462 ();
 sg13g2_fill_2 FILLER_33_3490 ();
 sg13g2_fill_1 FILLER_33_3531 ();
 sg13g2_decap_8 FILLER_33_3545 ();
 sg13g2_decap_8 FILLER_33_3552 ();
 sg13g2_decap_8 FILLER_33_3559 ();
 sg13g2_decap_8 FILLER_33_3566 ();
 sg13g2_decap_8 FILLER_33_3573 ();
 sg13g2_decap_8 FILLER_34_26 ();
 sg13g2_decap_8 FILLER_34_33 ();
 sg13g2_fill_2 FILLER_34_40 ();
 sg13g2_fill_1 FILLER_34_52 ();
 sg13g2_fill_2 FILLER_34_84 ();
 sg13g2_fill_2 FILLER_34_97 ();
 sg13g2_decap_8 FILLER_34_138 ();
 sg13g2_decap_4 FILLER_34_145 ();
 sg13g2_fill_1 FILLER_34_158 ();
 sg13g2_fill_2 FILLER_34_187 ();
 sg13g2_fill_2 FILLER_34_215 ();
 sg13g2_fill_1 FILLER_34_217 ();
 sg13g2_fill_2 FILLER_34_232 ();
 sg13g2_fill_1 FILLER_34_234 ();
 sg13g2_fill_1 FILLER_34_247 ();
 sg13g2_decap_8 FILLER_34_256 ();
 sg13g2_fill_2 FILLER_34_263 ();
 sg13g2_fill_2 FILLER_34_283 ();
 sg13g2_fill_1 FILLER_34_285 ();
 sg13g2_fill_1 FILLER_34_300 ();
 sg13g2_decap_4 FILLER_34_355 ();
 sg13g2_fill_1 FILLER_34_359 ();
 sg13g2_fill_2 FILLER_34_413 ();
 sg13g2_fill_1 FILLER_34_415 ();
 sg13g2_decap_4 FILLER_34_424 ();
 sg13g2_fill_2 FILLER_34_457 ();
 sg13g2_decap_8 FILLER_34_518 ();
 sg13g2_fill_1 FILLER_34_525 ();
 sg13g2_decap_8 FILLER_34_530 ();
 sg13g2_fill_2 FILLER_34_565 ();
 sg13g2_fill_2 FILLER_34_600 ();
 sg13g2_fill_1 FILLER_34_602 ();
 sg13g2_fill_1 FILLER_34_608 ();
 sg13g2_decap_8 FILLER_34_649 ();
 sg13g2_decap_4 FILLER_34_656 ();
 sg13g2_fill_1 FILLER_34_686 ();
 sg13g2_fill_1 FILLER_34_705 ();
 sg13g2_fill_1 FILLER_34_741 ();
 sg13g2_fill_1 FILLER_34_751 ();
 sg13g2_fill_1 FILLER_34_757 ();
 sg13g2_fill_2 FILLER_34_824 ();
 sg13g2_fill_1 FILLER_34_826 ();
 sg13g2_fill_1 FILLER_34_837 ();
 sg13g2_decap_8 FILLER_34_908 ();
 sg13g2_decap_4 FILLER_34_919 ();
 sg13g2_fill_1 FILLER_34_923 ();
 sg13g2_decap_8 FILLER_34_973 ();
 sg13g2_decap_4 FILLER_34_980 ();
 sg13g2_fill_2 FILLER_34_984 ();
 sg13g2_fill_2 FILLER_34_995 ();
 sg13g2_fill_1 FILLER_34_997 ();
 sg13g2_decap_4 FILLER_34_1003 ();
 sg13g2_fill_2 FILLER_34_1007 ();
 sg13g2_fill_2 FILLER_34_1044 ();
 sg13g2_fill_2 FILLER_34_1074 ();
 sg13g2_fill_1 FILLER_34_1076 ();
 sg13g2_fill_2 FILLER_34_1105 ();
 sg13g2_fill_1 FILLER_34_1138 ();
 sg13g2_decap_4 FILLER_34_1166 ();
 sg13g2_decap_4 FILLER_34_1192 ();
 sg13g2_fill_2 FILLER_34_1196 ();
 sg13g2_fill_1 FILLER_34_1235 ();
 sg13g2_fill_1 FILLER_34_1242 ();
 sg13g2_decap_4 FILLER_34_1248 ();
 sg13g2_fill_2 FILLER_34_1257 ();
 sg13g2_fill_1 FILLER_34_1259 ();
 sg13g2_fill_1 FILLER_34_1265 ();
 sg13g2_decap_4 FILLER_34_1292 ();
 sg13g2_fill_1 FILLER_34_1301 ();
 sg13g2_decap_8 FILLER_34_1306 ();
 sg13g2_decap_4 FILLER_34_1313 ();
 sg13g2_fill_1 FILLER_34_1317 ();
 sg13g2_decap_8 FILLER_34_1343 ();
 sg13g2_decap_8 FILLER_34_1350 ();
 sg13g2_fill_1 FILLER_34_1357 ();
 sg13g2_decap_8 FILLER_34_1402 ();
 sg13g2_decap_8 FILLER_34_1414 ();
 sg13g2_fill_1 FILLER_34_1421 ();
 sg13g2_fill_2 FILLER_34_1432 ();
 sg13g2_fill_2 FILLER_34_1439 ();
 sg13g2_fill_1 FILLER_34_1474 ();
 sg13g2_fill_2 FILLER_34_1498 ();
 sg13g2_fill_1 FILLER_34_1500 ();
 sg13g2_fill_2 FILLER_34_1508 ();
 sg13g2_fill_1 FILLER_34_1510 ();
 sg13g2_fill_2 FILLER_34_1521 ();
 sg13g2_fill_2 FILLER_34_1532 ();
 sg13g2_fill_1 FILLER_34_1534 ();
 sg13g2_fill_1 FILLER_34_1544 ();
 sg13g2_fill_2 FILLER_34_1555 ();
 sg13g2_fill_1 FILLER_34_1656 ();
 sg13g2_fill_2 FILLER_34_1667 ();
 sg13g2_fill_2 FILLER_34_1673 ();
 sg13g2_fill_1 FILLER_34_1684 ();
 sg13g2_decap_8 FILLER_34_1694 ();
 sg13g2_decap_4 FILLER_34_1714 ();
 sg13g2_decap_4 FILLER_34_1726 ();
 sg13g2_fill_2 FILLER_34_1730 ();
 sg13g2_fill_2 FILLER_34_1736 ();
 sg13g2_fill_1 FILLER_34_1738 ();
 sg13g2_fill_1 FILLER_34_1744 ();
 sg13g2_fill_2 FILLER_34_1749 ();
 sg13g2_fill_1 FILLER_34_1751 ();
 sg13g2_decap_8 FILLER_34_1767 ();
 sg13g2_fill_2 FILLER_34_1774 ();
 sg13g2_fill_2 FILLER_34_1781 ();
 sg13g2_fill_2 FILLER_34_1807 ();
 sg13g2_fill_1 FILLER_34_1835 ();
 sg13g2_decap_8 FILLER_34_1851 ();
 sg13g2_fill_2 FILLER_34_1858 ();
 sg13g2_decap_8 FILLER_34_1865 ();
 sg13g2_fill_2 FILLER_34_1872 ();
 sg13g2_fill_1 FILLER_34_1902 ();
 sg13g2_fill_2 FILLER_34_1914 ();
 sg13g2_fill_1 FILLER_34_1916 ();
 sg13g2_fill_1 FILLER_34_1943 ();
 sg13g2_decap_4 FILLER_34_1948 ();
 sg13g2_fill_2 FILLER_34_1952 ();
 sg13g2_decap_8 FILLER_34_1964 ();
 sg13g2_decap_4 FILLER_34_1971 ();
 sg13g2_fill_2 FILLER_34_1975 ();
 sg13g2_decap_4 FILLER_34_2001 ();
 sg13g2_fill_2 FILLER_34_2005 ();
 sg13g2_decap_8 FILLER_34_2011 ();
 sg13g2_decap_8 FILLER_34_2018 ();
 sg13g2_fill_2 FILLER_34_2025 ();
 sg13g2_fill_1 FILLER_34_2027 ();
 sg13g2_decap_8 FILLER_34_2032 ();
 sg13g2_fill_2 FILLER_34_2047 ();
 sg13g2_fill_1 FILLER_34_2049 ();
 sg13g2_decap_8 FILLER_34_2070 ();
 sg13g2_decap_8 FILLER_34_2077 ();
 sg13g2_fill_2 FILLER_34_2084 ();
 sg13g2_fill_1 FILLER_34_2086 ();
 sg13g2_decap_4 FILLER_34_2120 ();
 sg13g2_fill_1 FILLER_34_2124 ();
 sg13g2_fill_2 FILLER_34_2137 ();
 sg13g2_fill_1 FILLER_34_2139 ();
 sg13g2_fill_2 FILLER_34_2154 ();
 sg13g2_fill_1 FILLER_34_2156 ();
 sg13g2_decap_8 FILLER_34_2165 ();
 sg13g2_decap_8 FILLER_34_2172 ();
 sg13g2_fill_2 FILLER_34_2179 ();
 sg13g2_fill_1 FILLER_34_2181 ();
 sg13g2_decap_8 FILLER_34_2195 ();
 sg13g2_decap_8 FILLER_34_2202 ();
 sg13g2_decap_8 FILLER_34_2209 ();
 sg13g2_fill_1 FILLER_34_2216 ();
 sg13g2_decap_8 FILLER_34_2225 ();
 sg13g2_decap_8 FILLER_34_2232 ();
 sg13g2_decap_8 FILLER_34_2239 ();
 sg13g2_decap_4 FILLER_34_2246 ();
 sg13g2_decap_8 FILLER_34_2255 ();
 sg13g2_decap_8 FILLER_34_2262 ();
 sg13g2_decap_8 FILLER_34_2269 ();
 sg13g2_decap_4 FILLER_34_2276 ();
 sg13g2_fill_1 FILLER_34_2280 ();
 sg13g2_decap_4 FILLER_34_2285 ();
 sg13g2_fill_1 FILLER_34_2289 ();
 sg13g2_fill_1 FILLER_34_2312 ();
 sg13g2_decap_8 FILLER_34_2333 ();
 sg13g2_decap_4 FILLER_34_2340 ();
 sg13g2_fill_1 FILLER_34_2344 ();
 sg13g2_fill_1 FILLER_34_2358 ();
 sg13g2_fill_2 FILLER_34_2368 ();
 sg13g2_fill_1 FILLER_34_2370 ();
 sg13g2_decap_4 FILLER_34_2376 ();
 sg13g2_fill_1 FILLER_34_2380 ();
 sg13g2_fill_2 FILLER_34_2404 ();
 sg13g2_fill_2 FILLER_34_2419 ();
 sg13g2_fill_1 FILLER_34_2444 ();
 sg13g2_decap_8 FILLER_34_2475 ();
 sg13g2_decap_8 FILLER_34_2482 ();
 sg13g2_decap_4 FILLER_34_2489 ();
 sg13g2_fill_1 FILLER_34_2493 ();
 sg13g2_decap_8 FILLER_34_2498 ();
 sg13g2_decap_8 FILLER_34_2505 ();
 sg13g2_fill_2 FILLER_34_2512 ();
 sg13g2_decap_8 FILLER_34_2570 ();
 sg13g2_decap_4 FILLER_34_2577 ();
 sg13g2_fill_2 FILLER_34_2581 ();
 sg13g2_fill_2 FILLER_34_2612 ();
 sg13g2_decap_8 FILLER_34_2640 ();
 sg13g2_decap_4 FILLER_34_2647 ();
 sg13g2_fill_2 FILLER_34_2651 ();
 sg13g2_fill_1 FILLER_34_2692 ();
 sg13g2_decap_4 FILLER_34_2701 ();
 sg13g2_fill_1 FILLER_34_2705 ();
 sg13g2_fill_1 FILLER_34_2732 ();
 sg13g2_fill_1 FILLER_34_2747 ();
 sg13g2_fill_1 FILLER_34_2779 ();
 sg13g2_fill_1 FILLER_34_2800 ();
 sg13g2_decap_4 FILLER_34_2809 ();
 sg13g2_decap_4 FILLER_34_2865 ();
 sg13g2_decap_8 FILLER_34_2882 ();
 sg13g2_fill_1 FILLER_34_2889 ();
 sg13g2_decap_8 FILLER_34_2895 ();
 sg13g2_fill_1 FILLER_34_2902 ();
 sg13g2_fill_1 FILLER_34_2938 ();
 sg13g2_fill_1 FILLER_34_2952 ();
 sg13g2_fill_2 FILLER_34_2957 ();
 sg13g2_fill_1 FILLER_34_2959 ();
 sg13g2_decap_8 FILLER_34_2986 ();
 sg13g2_decap_8 FILLER_34_2993 ();
 sg13g2_fill_2 FILLER_34_3000 ();
 sg13g2_fill_1 FILLER_34_3002 ();
 sg13g2_fill_1 FILLER_34_3021 ();
 sg13g2_fill_2 FILLER_34_3027 ();
 sg13g2_fill_1 FILLER_34_3039 ();
 sg13g2_fill_2 FILLER_34_3054 ();
 sg13g2_fill_2 FILLER_34_3117 ();
 sg13g2_fill_1 FILLER_34_3119 ();
 sg13g2_fill_2 FILLER_34_3174 ();
 sg13g2_fill_1 FILLER_34_3176 ();
 sg13g2_fill_2 FILLER_34_3192 ();
 sg13g2_fill_1 FILLER_34_3194 ();
 sg13g2_fill_1 FILLER_34_3208 ();
 sg13g2_fill_2 FILLER_34_3240 ();
 sg13g2_decap_8 FILLER_34_3268 ();
 sg13g2_fill_2 FILLER_34_3275 ();
 sg13g2_fill_1 FILLER_34_3313 ();
 sg13g2_decap_8 FILLER_34_3334 ();
 sg13g2_fill_2 FILLER_34_3341 ();
 sg13g2_fill_2 FILLER_34_3348 ();
 sg13g2_fill_1 FILLER_34_3350 ();
 sg13g2_fill_2 FILLER_34_3365 ();
 sg13g2_fill_1 FILLER_34_3367 ();
 sg13g2_fill_1 FILLER_34_3394 ();
 sg13g2_decap_8 FILLER_34_3426 ();
 sg13g2_fill_2 FILLER_34_3433 ();
 sg13g2_fill_1 FILLER_34_3439 ();
 sg13g2_decap_8 FILLER_34_3455 ();
 sg13g2_fill_2 FILLER_34_3462 ();
 sg13g2_fill_2 FILLER_34_3473 ();
 sg13g2_fill_1 FILLER_34_3479 ();
 sg13g2_fill_1 FILLER_34_3489 ();
 sg13g2_decap_8 FILLER_34_3547 ();
 sg13g2_decap_8 FILLER_34_3554 ();
 sg13g2_decap_8 FILLER_34_3561 ();
 sg13g2_decap_8 FILLER_34_3568 ();
 sg13g2_decap_4 FILLER_34_3575 ();
 sg13g2_fill_1 FILLER_34_3579 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_fill_2 FILLER_35_14 ();
 sg13g2_fill_1 FILLER_35_16 ();
 sg13g2_fill_2 FILLER_35_43 ();
 sg13g2_fill_2 FILLER_35_50 ();
 sg13g2_fill_1 FILLER_35_69 ();
 sg13g2_fill_2 FILLER_35_96 ();
 sg13g2_fill_2 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_118 ();
 sg13g2_fill_2 FILLER_35_125 ();
 sg13g2_decap_8 FILLER_35_135 ();
 sg13g2_fill_2 FILLER_35_142 ();
 sg13g2_fill_1 FILLER_35_144 ();
 sg13g2_fill_1 FILLER_35_171 ();
 sg13g2_decap_8 FILLER_35_263 ();
 sg13g2_fill_2 FILLER_35_308 ();
 sg13g2_fill_1 FILLER_35_326 ();
 sg13g2_fill_1 FILLER_35_332 ();
 sg13g2_decap_8 FILLER_35_351 ();
 sg13g2_fill_1 FILLER_35_358 ();
 sg13g2_decap_4 FILLER_35_363 ();
 sg13g2_fill_1 FILLER_35_367 ();
 sg13g2_fill_2 FILLER_35_373 ();
 sg13g2_fill_2 FILLER_35_388 ();
 sg13g2_fill_1 FILLER_35_390 ();
 sg13g2_decap_4 FILLER_35_425 ();
 sg13g2_fill_2 FILLER_35_429 ();
 sg13g2_fill_2 FILLER_35_436 ();
 sg13g2_fill_1 FILLER_35_438 ();
 sg13g2_decap_4 FILLER_35_444 ();
 sg13g2_fill_1 FILLER_35_448 ();
 sg13g2_fill_2 FILLER_35_488 ();
 sg13g2_fill_2 FILLER_35_499 ();
 sg13g2_fill_2 FILLER_35_514 ();
 sg13g2_fill_1 FILLER_35_558 ();
 sg13g2_fill_2 FILLER_35_562 ();
 sg13g2_fill_2 FILLER_35_586 ();
 sg13g2_fill_1 FILLER_35_588 ();
 sg13g2_fill_2 FILLER_35_602 ();
 sg13g2_fill_1 FILLER_35_604 ();
 sg13g2_decap_8 FILLER_35_610 ();
 sg13g2_fill_1 FILLER_35_617 ();
 sg13g2_decap_4 FILLER_35_635 ();
 sg13g2_fill_2 FILLER_35_643 ();
 sg13g2_fill_2 FILLER_35_669 ();
 sg13g2_fill_1 FILLER_35_689 ();
 sg13g2_fill_1 FILLER_35_704 ();
 sg13g2_fill_1 FILLER_35_717 ();
 sg13g2_fill_1 FILLER_35_735 ();
 sg13g2_decap_4 FILLER_35_754 ();
 sg13g2_decap_8 FILLER_35_784 ();
 sg13g2_decap_4 FILLER_35_791 ();
 sg13g2_fill_1 FILLER_35_795 ();
 sg13g2_decap_8 FILLER_35_801 ();
 sg13g2_decap_8 FILLER_35_808 ();
 sg13g2_decap_8 FILLER_35_820 ();
 sg13g2_fill_2 FILLER_35_827 ();
 sg13g2_fill_1 FILLER_35_829 ();
 sg13g2_fill_2 FILLER_35_840 ();
 sg13g2_decap_8 FILLER_35_847 ();
 sg13g2_fill_2 FILLER_35_854 ();
 sg13g2_fill_1 FILLER_35_856 ();
 sg13g2_fill_2 FILLER_35_862 ();
 sg13g2_fill_1 FILLER_35_876 ();
 sg13g2_decap_8 FILLER_35_883 ();
 sg13g2_decap_8 FILLER_35_890 ();
 sg13g2_fill_2 FILLER_35_897 ();
 sg13g2_fill_1 FILLER_35_899 ();
 sg13g2_fill_2 FILLER_35_908 ();
 sg13g2_decap_4 FILLER_35_915 ();
 sg13g2_fill_2 FILLER_35_919 ();
 sg13g2_fill_1 FILLER_35_933 ();
 sg13g2_fill_1 FILLER_35_946 ();
 sg13g2_fill_1 FILLER_35_956 ();
 sg13g2_decap_8 FILLER_35_974 ();
 sg13g2_decap_4 FILLER_35_1015 ();
 sg13g2_fill_1 FILLER_35_1019 ();
 sg13g2_decap_8 FILLER_35_1024 ();
 sg13g2_decap_4 FILLER_35_1031 ();
 sg13g2_fill_1 FILLER_35_1035 ();
 sg13g2_decap_4 FILLER_35_1053 ();
 sg13g2_fill_1 FILLER_35_1057 ();
 sg13g2_fill_1 FILLER_35_1088 ();
 sg13g2_decap_4 FILLER_35_1117 ();
 sg13g2_fill_1 FILLER_35_1121 ();
 sg13g2_decap_8 FILLER_35_1126 ();
 sg13g2_decap_8 FILLER_35_1133 ();
 sg13g2_decap_4 FILLER_35_1140 ();
 sg13g2_fill_1 FILLER_35_1144 ();
 sg13g2_decap_4 FILLER_35_1153 ();
 sg13g2_fill_1 FILLER_35_1157 ();
 sg13g2_fill_1 FILLER_35_1163 ();
 sg13g2_fill_1 FILLER_35_1208 ();
 sg13g2_decap_4 FILLER_35_1254 ();
 sg13g2_fill_2 FILLER_35_1275 ();
 sg13g2_decap_8 FILLER_35_1281 ();
 sg13g2_decap_4 FILLER_35_1288 ();
 sg13g2_fill_1 FILLER_35_1292 ();
 sg13g2_decap_4 FILLER_35_1301 ();
 sg13g2_fill_1 FILLER_35_1305 ();
 sg13g2_decap_8 FILLER_35_1311 ();
 sg13g2_decap_8 FILLER_35_1318 ();
 sg13g2_decap_4 FILLER_35_1325 ();
 sg13g2_fill_2 FILLER_35_1329 ();
 sg13g2_decap_4 FILLER_35_1345 ();
 sg13g2_decap_8 FILLER_35_1379 ();
 sg13g2_decap_4 FILLER_35_1386 ();
 sg13g2_fill_1 FILLER_35_1445 ();
 sg13g2_decap_4 FILLER_35_1454 ();
 sg13g2_fill_2 FILLER_35_1468 ();
 sg13g2_fill_1 FILLER_35_1470 ();
 sg13g2_fill_2 FILLER_35_1518 ();
 sg13g2_fill_1 FILLER_35_1520 ();
 sg13g2_decap_4 FILLER_35_1531 ();
 sg13g2_fill_2 FILLER_35_1573 ();
 sg13g2_fill_1 FILLER_35_1575 ();
 sg13g2_fill_2 FILLER_35_1580 ();
 sg13g2_fill_2 FILLER_35_1608 ();
 sg13g2_fill_2 FILLER_35_1641 ();
 sg13g2_fill_1 FILLER_35_1652 ();
 sg13g2_decap_8 FILLER_35_1656 ();
 sg13g2_decap_8 FILLER_35_1663 ();
 sg13g2_decap_4 FILLER_35_1670 ();
 sg13g2_fill_1 FILLER_35_1674 ();
 sg13g2_decap_4 FILLER_35_1701 ();
 sg13g2_fill_1 FILLER_35_1705 ();
 sg13g2_fill_2 FILLER_35_1714 ();
 sg13g2_fill_1 FILLER_35_1716 ();
 sg13g2_fill_1 FILLER_35_1748 ();
 sg13g2_fill_2 FILLER_35_1774 ();
 sg13g2_fill_2 FILLER_35_1781 ();
 sg13g2_fill_1 FILLER_35_1783 ();
 sg13g2_decap_8 FILLER_35_1788 ();
 sg13g2_fill_2 FILLER_35_1795 ();
 sg13g2_fill_1 FILLER_35_1797 ();
 sg13g2_decap_8 FILLER_35_1806 ();
 sg13g2_fill_1 FILLER_35_1813 ();
 sg13g2_decap_8 FILLER_35_1818 ();
 sg13g2_decap_4 FILLER_35_1825 ();
 sg13g2_fill_2 FILLER_35_1851 ();
 sg13g2_decap_8 FILLER_35_1857 ();
 sg13g2_decap_8 FILLER_35_1877 ();
 sg13g2_fill_1 FILLER_35_1884 ();
 sg13g2_fill_1 FILLER_35_1913 ();
 sg13g2_fill_2 FILLER_35_1959 ();
 sg13g2_decap_8 FILLER_35_2038 ();
 sg13g2_decap_8 FILLER_35_2045 ();
 sg13g2_decap_4 FILLER_35_2076 ();
 sg13g2_decap_8 FILLER_35_2108 ();
 sg13g2_decap_8 FILLER_35_2115 ();
 sg13g2_fill_2 FILLER_35_2122 ();
 sg13g2_decap_4 FILLER_35_2139 ();
 sg13g2_decap_8 FILLER_35_2156 ();
 sg13g2_decap_8 FILLER_35_2168 ();
 sg13g2_fill_2 FILLER_35_2175 ();
 sg13g2_fill_2 FILLER_35_2210 ();
 sg13g2_fill_2 FILLER_35_2231 ();
 sg13g2_fill_1 FILLER_35_2233 ();
 sg13g2_decap_4 FILLER_35_2243 ();
 sg13g2_fill_2 FILLER_35_2247 ();
 sg13g2_decap_4 FILLER_35_2257 ();
 sg13g2_decap_4 FILLER_35_2264 ();
 sg13g2_decap_4 FILLER_35_2291 ();
 sg13g2_fill_2 FILLER_35_2295 ();
 sg13g2_decap_4 FILLER_35_2302 ();
 sg13g2_decap_4 FILLER_35_2315 ();
 sg13g2_fill_1 FILLER_35_2319 ();
 sg13g2_decap_4 FILLER_35_2349 ();
 sg13g2_fill_1 FILLER_35_2353 ();
 sg13g2_fill_2 FILLER_35_2364 ();
 sg13g2_fill_2 FILLER_35_2381 ();
 sg13g2_fill_1 FILLER_35_2383 ();
 sg13g2_fill_2 FILLER_35_2402 ();
 sg13g2_fill_1 FILLER_35_2404 ();
 sg13g2_decap_8 FILLER_35_2538 ();
 sg13g2_decap_4 FILLER_35_2545 ();
 sg13g2_fill_1 FILLER_35_2549 ();
 sg13g2_fill_1 FILLER_35_2554 ();
 sg13g2_fill_1 FILLER_35_2581 ();
 sg13g2_fill_2 FILLER_35_2587 ();
 sg13g2_fill_2 FILLER_35_2602 ();
 sg13g2_fill_1 FILLER_35_2624 ();
 sg13g2_fill_1 FILLER_35_2629 ();
 sg13g2_decap_4 FILLER_35_2640 ();
 sg13g2_fill_1 FILLER_35_2644 ();
 sg13g2_decap_8 FILLER_35_2650 ();
 sg13g2_decap_8 FILLER_35_2661 ();
 sg13g2_decap_8 FILLER_35_2668 ();
 sg13g2_fill_1 FILLER_35_2675 ();
 sg13g2_decap_4 FILLER_35_2684 ();
 sg13g2_fill_1 FILLER_35_2688 ();
 sg13g2_fill_2 FILLER_35_2720 ();
 sg13g2_fill_1 FILLER_35_2727 ();
 sg13g2_fill_1 FILLER_35_2732 ();
 sg13g2_decap_4 FILLER_35_2819 ();
 sg13g2_fill_1 FILLER_35_2823 ();
 sg13g2_decap_4 FILLER_35_2828 ();
 sg13g2_fill_1 FILLER_35_2832 ();
 sg13g2_fill_2 FILLER_35_2838 ();
 sg13g2_fill_1 FILLER_35_2840 ();
 sg13g2_decap_4 FILLER_35_2846 ();
 sg13g2_decap_4 FILLER_35_2858 ();
 sg13g2_fill_1 FILLER_35_2862 ();
 sg13g2_decap_8 FILLER_35_2895 ();
 sg13g2_decap_4 FILLER_35_2902 ();
 sg13g2_fill_1 FILLER_35_2915 ();
 sg13g2_decap_8 FILLER_35_2920 ();
 sg13g2_fill_2 FILLER_35_2953 ();
 sg13g2_fill_2 FILLER_35_2964 ();
 sg13g2_fill_1 FILLER_35_2966 ();
 sg13g2_fill_2 FILLER_35_2984 ();
 sg13g2_decap_4 FILLER_35_3056 ();
 sg13g2_fill_2 FILLER_35_3073 ();
 sg13g2_fill_1 FILLER_35_3075 ();
 sg13g2_decap_8 FILLER_35_3080 ();
 sg13g2_decap_8 FILLER_35_3087 ();
 sg13g2_decap_8 FILLER_35_3094 ();
 sg13g2_fill_2 FILLER_35_3101 ();
 sg13g2_fill_2 FILLER_35_3112 ();
 sg13g2_fill_1 FILLER_35_3118 ();
 sg13g2_fill_2 FILLER_35_3128 ();
 sg13g2_fill_1 FILLER_35_3130 ();
 sg13g2_fill_2 FILLER_35_3135 ();
 sg13g2_decap_4 FILLER_35_3168 ();
 sg13g2_fill_1 FILLER_35_3172 ();
 sg13g2_fill_2 FILLER_35_3182 ();
 sg13g2_fill_2 FILLER_35_3190 ();
 sg13g2_fill_2 FILLER_35_3197 ();
 sg13g2_decap_8 FILLER_35_3216 ();
 sg13g2_fill_1 FILLER_35_3232 ();
 sg13g2_decap_8 FILLER_35_3237 ();
 sg13g2_decap_4 FILLER_35_3244 ();
 sg13g2_fill_1 FILLER_35_3248 ();
 sg13g2_decap_8 FILLER_35_3263 ();
 sg13g2_decap_4 FILLER_35_3301 ();
 sg13g2_fill_2 FILLER_35_3305 ();
 sg13g2_decap_4 FILLER_35_3316 ();
 sg13g2_fill_1 FILLER_35_3320 ();
 sg13g2_decap_8 FILLER_35_3334 ();
 sg13g2_fill_2 FILLER_35_3341 ();
 sg13g2_fill_1 FILLER_35_3351 ();
 sg13g2_fill_2 FILLER_35_3387 ();
 sg13g2_fill_1 FILLER_35_3389 ();
 sg13g2_decap_4 FILLER_35_3421 ();
 sg13g2_decap_8 FILLER_35_3491 ();
 sg13g2_fill_2 FILLER_35_3498 ();
 sg13g2_fill_1 FILLER_35_3500 ();
 sg13g2_decap_8 FILLER_35_3505 ();
 sg13g2_decap_8 FILLER_35_3512 ();
 sg13g2_decap_8 FILLER_35_3519 ();
 sg13g2_decap_8 FILLER_35_3526 ();
 sg13g2_decap_8 FILLER_35_3533 ();
 sg13g2_decap_8 FILLER_35_3540 ();
 sg13g2_decap_8 FILLER_35_3547 ();
 sg13g2_decap_8 FILLER_35_3554 ();
 sg13g2_decap_8 FILLER_35_3561 ();
 sg13g2_decap_8 FILLER_35_3568 ();
 sg13g2_decap_4 FILLER_35_3575 ();
 sg13g2_fill_1 FILLER_35_3579 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_fill_1 FILLER_36_21 ();
 sg13g2_fill_2 FILLER_36_70 ();
 sg13g2_fill_2 FILLER_36_82 ();
 sg13g2_fill_2 FILLER_36_88 ();
 sg13g2_fill_2 FILLER_36_107 ();
 sg13g2_fill_2 FILLER_36_114 ();
 sg13g2_fill_1 FILLER_36_116 ();
 sg13g2_decap_8 FILLER_36_130 ();
 sg13g2_fill_1 FILLER_36_137 ();
 sg13g2_fill_2 FILLER_36_142 ();
 sg13g2_fill_1 FILLER_36_144 ();
 sg13g2_fill_1 FILLER_36_150 ();
 sg13g2_decap_8 FILLER_36_176 ();
 sg13g2_decap_4 FILLER_36_183 ();
 sg13g2_fill_1 FILLER_36_218 ();
 sg13g2_fill_2 FILLER_36_246 ();
 sg13g2_fill_2 FILLER_36_252 ();
 sg13g2_fill_1 FILLER_36_258 ();
 sg13g2_decap_8 FILLER_36_264 ();
 sg13g2_decap_8 FILLER_36_271 ();
 sg13g2_decap_4 FILLER_36_278 ();
 sg13g2_fill_2 FILLER_36_287 ();
 sg13g2_fill_1 FILLER_36_289 ();
 sg13g2_decap_8 FILLER_36_300 ();
 sg13g2_fill_2 FILLER_36_307 ();
 sg13g2_fill_1 FILLER_36_319 ();
 sg13g2_decap_4 FILLER_36_343 ();
 sg13g2_fill_2 FILLER_36_347 ();
 sg13g2_fill_2 FILLER_36_375 ();
 sg13g2_fill_1 FILLER_36_386 ();
 sg13g2_decap_8 FILLER_36_413 ();
 sg13g2_fill_1 FILLER_36_420 ();
 sg13g2_fill_1 FILLER_36_441 ();
 sg13g2_decap_8 FILLER_36_452 ();
 sg13g2_decap_4 FILLER_36_459 ();
 sg13g2_fill_2 FILLER_36_463 ();
 sg13g2_fill_2 FILLER_36_481 ();
 sg13g2_fill_1 FILLER_36_483 ();
 sg13g2_fill_2 FILLER_36_493 ();
 sg13g2_fill_1 FILLER_36_495 ();
 sg13g2_fill_1 FILLER_36_563 ();
 sg13g2_fill_2 FILLER_36_625 ();
 sg13g2_fill_2 FILLER_36_663 ();
 sg13g2_fill_2 FILLER_36_705 ();
 sg13g2_fill_2 FILLER_36_738 ();
 sg13g2_fill_1 FILLER_36_740 ();
 sg13g2_decap_4 FILLER_36_788 ();
 sg13g2_fill_1 FILLER_36_792 ();
 sg13g2_decap_4 FILLER_36_808 ();
 sg13g2_fill_2 FILLER_36_822 ();
 sg13g2_fill_1 FILLER_36_824 ();
 sg13g2_fill_2 FILLER_36_835 ();
 sg13g2_fill_2 FILLER_36_847 ();
 sg13g2_fill_2 FILLER_36_857 ();
 sg13g2_fill_1 FILLER_36_859 ();
 sg13g2_fill_2 FILLER_36_865 ();
 sg13g2_fill_1 FILLER_36_867 ();
 sg13g2_fill_1 FILLER_36_876 ();
 sg13g2_decap_8 FILLER_36_894 ();
 sg13g2_fill_2 FILLER_36_901 ();
 sg13g2_fill_2 FILLER_36_907 ();
 sg13g2_fill_1 FILLER_36_909 ();
 sg13g2_fill_1 FILLER_36_949 ();
 sg13g2_decap_4 FILLER_36_980 ();
 sg13g2_fill_1 FILLER_36_984 ();
 sg13g2_fill_2 FILLER_36_993 ();
 sg13g2_fill_1 FILLER_36_995 ();
 sg13g2_fill_2 FILLER_36_1005 ();
 sg13g2_fill_2 FILLER_36_1016 ();
 sg13g2_fill_1 FILLER_36_1018 ();
 sg13g2_decap_8 FILLER_36_1023 ();
 sg13g2_decap_4 FILLER_36_1030 ();
 sg13g2_fill_2 FILLER_36_1034 ();
 sg13g2_fill_2 FILLER_36_1055 ();
 sg13g2_fill_1 FILLER_36_1057 ();
 sg13g2_fill_2 FILLER_36_1062 ();
 sg13g2_fill_1 FILLER_36_1064 ();
 sg13g2_fill_1 FILLER_36_1087 ();
 sg13g2_fill_2 FILLER_36_1092 ();
 sg13g2_fill_1 FILLER_36_1094 ();
 sg13g2_fill_2 FILLER_36_1129 ();
 sg13g2_fill_1 FILLER_36_1131 ();
 sg13g2_fill_1 FILLER_36_1140 ();
 sg13g2_decap_4 FILLER_36_1146 ();
 sg13g2_fill_2 FILLER_36_1150 ();
 sg13g2_decap_4 FILLER_36_1162 ();
 sg13g2_decap_4 FILLER_36_1180 ();
 sg13g2_fill_1 FILLER_36_1184 ();
 sg13g2_decap_4 FILLER_36_1189 ();
 sg13g2_fill_2 FILLER_36_1193 ();
 sg13g2_fill_1 FILLER_36_1219 ();
 sg13g2_fill_1 FILLER_36_1224 ();
 sg13g2_fill_2 FILLER_36_1236 ();
 sg13g2_fill_1 FILLER_36_1238 ();
 sg13g2_decap_8 FILLER_36_1243 ();
 sg13g2_fill_1 FILLER_36_1259 ();
 sg13g2_fill_2 FILLER_36_1303 ();
 sg13g2_fill_2 FILLER_36_1323 ();
 sg13g2_fill_1 FILLER_36_1325 ();
 sg13g2_fill_1 FILLER_36_1376 ();
 sg13g2_fill_2 FILLER_36_1381 ();
 sg13g2_fill_1 FILLER_36_1383 ();
 sg13g2_decap_4 FILLER_36_1397 ();
 sg13g2_fill_2 FILLER_36_1405 ();
 sg13g2_fill_1 FILLER_36_1407 ();
 sg13g2_fill_2 FILLER_36_1422 ();
 sg13g2_decap_8 FILLER_36_1443 ();
 sg13g2_fill_1 FILLER_36_1450 ();
 sg13g2_fill_2 FILLER_36_1459 ();
 sg13g2_fill_2 FILLER_36_1466 ();
 sg13g2_fill_1 FILLER_36_1499 ();
 sg13g2_decap_8 FILLER_36_1506 ();
 sg13g2_fill_2 FILLER_36_1513 ();
 sg13g2_fill_1 FILLER_36_1520 ();
 sg13g2_fill_1 FILLER_36_1524 ();
 sg13g2_decap_8 FILLER_36_1530 ();
 sg13g2_decap_4 FILLER_36_1537 ();
 sg13g2_decap_4 FILLER_36_1554 ();
 sg13g2_fill_2 FILLER_36_1558 ();
 sg13g2_fill_2 FILLER_36_1565 ();
 sg13g2_fill_1 FILLER_36_1567 ();
 sg13g2_decap_4 FILLER_36_1573 ();
 sg13g2_fill_2 FILLER_36_1577 ();
 sg13g2_decap_4 FILLER_36_1584 ();
 sg13g2_decap_8 FILLER_36_1606 ();
 sg13g2_decap_8 FILLER_36_1613 ();
 sg13g2_decap_8 FILLER_36_1620 ();
 sg13g2_fill_2 FILLER_36_1627 ();
 sg13g2_fill_2 FILLER_36_1638 ();
 sg13g2_fill_1 FILLER_36_1640 ();
 sg13g2_fill_2 FILLER_36_1667 ();
 sg13g2_decap_8 FILLER_36_1673 ();
 sg13g2_decap_4 FILLER_36_1680 ();
 sg13g2_decap_8 FILLER_36_1689 ();
 sg13g2_decap_8 FILLER_36_1715 ();
 sg13g2_fill_2 FILLER_36_1722 ();
 sg13g2_fill_2 FILLER_36_1736 ();
 sg13g2_decap_4 FILLER_36_1747 ();
 sg13g2_fill_1 FILLER_36_1751 ();
 sg13g2_decap_4 FILLER_36_1763 ();
 sg13g2_fill_2 FILLER_36_1767 ();
 sg13g2_decap_4 FILLER_36_1774 ();
 sg13g2_fill_1 FILLER_36_1778 ();
 sg13g2_fill_1 FILLER_36_1791 ();
 sg13g2_decap_8 FILLER_36_1798 ();
 sg13g2_decap_4 FILLER_36_1805 ();
 sg13g2_fill_2 FILLER_36_1835 ();
 sg13g2_fill_1 FILLER_36_1896 ();
 sg13g2_fill_1 FILLER_36_1932 ();
 sg13g2_fill_1 FILLER_36_1945 ();
 sg13g2_fill_1 FILLER_36_1971 ();
 sg13g2_decap_8 FILLER_36_1976 ();
 sg13g2_fill_2 FILLER_36_1983 ();
 sg13g2_fill_1 FILLER_36_1985 ();
 sg13g2_decap_8 FILLER_36_1994 ();
 sg13g2_decap_4 FILLER_36_2001 ();
 sg13g2_fill_1 FILLER_36_2005 ();
 sg13g2_decap_8 FILLER_36_2025 ();
 sg13g2_fill_2 FILLER_36_2032 ();
 sg13g2_fill_1 FILLER_36_2034 ();
 sg13g2_decap_8 FILLER_36_2040 ();
 sg13g2_fill_2 FILLER_36_2047 ();
 sg13g2_decap_8 FILLER_36_2081 ();
 sg13g2_decap_8 FILLER_36_2088 ();
 sg13g2_decap_8 FILLER_36_2095 ();
 sg13g2_fill_2 FILLER_36_2102 ();
 sg13g2_fill_1 FILLER_36_2104 ();
 sg13g2_fill_1 FILLER_36_2113 ();
 sg13g2_fill_2 FILLER_36_2129 ();
 sg13g2_fill_2 FILLER_36_2158 ();
 sg13g2_decap_8 FILLER_36_2184 ();
 sg13g2_fill_2 FILLER_36_2191 ();
 sg13g2_fill_1 FILLER_36_2193 ();
 sg13g2_fill_2 FILLER_36_2207 ();
 sg13g2_decap_8 FILLER_36_2228 ();
 sg13g2_fill_2 FILLER_36_2235 ();
 sg13g2_fill_1 FILLER_36_2269 ();
 sg13g2_decap_4 FILLER_36_2287 ();
 sg13g2_fill_2 FILLER_36_2291 ();
 sg13g2_fill_2 FILLER_36_2298 ();
 sg13g2_fill_1 FILLER_36_2300 ();
 sg13g2_decap_4 FILLER_36_2319 ();
 sg13g2_fill_1 FILLER_36_2336 ();
 sg13g2_fill_2 FILLER_36_2348 ();
 sg13g2_fill_1 FILLER_36_2350 ();
 sg13g2_fill_2 FILLER_36_2369 ();
 sg13g2_decap_8 FILLER_36_2380 ();
 sg13g2_decap_8 FILLER_36_2387 ();
 sg13g2_fill_2 FILLER_36_2394 ();
 sg13g2_fill_1 FILLER_36_2405 ();
 sg13g2_decap_8 FILLER_36_2421 ();
 sg13g2_fill_2 FILLER_36_2428 ();
 sg13g2_fill_1 FILLER_36_2430 ();
 sg13g2_fill_1 FILLER_36_2445 ();
 sg13g2_fill_2 FILLER_36_2473 ();
 sg13g2_fill_1 FILLER_36_2475 ();
 sg13g2_decap_8 FILLER_36_2498 ();
 sg13g2_decap_8 FILLER_36_2505 ();
 sg13g2_decap_8 FILLER_36_2512 ();
 sg13g2_decap_4 FILLER_36_2519 ();
 sg13g2_fill_1 FILLER_36_2523 ();
 sg13g2_fill_2 FILLER_36_2532 ();
 sg13g2_decap_8 FILLER_36_2566 ();
 sg13g2_fill_2 FILLER_36_2573 ();
 sg13g2_fill_2 FILLER_36_2582 ();
 sg13g2_fill_1 FILLER_36_2645 ();
 sg13g2_decap_8 FILLER_36_2672 ();
 sg13g2_decap_8 FILLER_36_2679 ();
 sg13g2_decap_8 FILLER_36_2686 ();
 sg13g2_fill_2 FILLER_36_2693 ();
 sg13g2_fill_1 FILLER_36_2695 ();
 sg13g2_fill_2 FILLER_36_2714 ();
 sg13g2_fill_1 FILLER_36_2716 ();
 sg13g2_decap_8 FILLER_36_2756 ();
 sg13g2_fill_2 FILLER_36_2763 ();
 sg13g2_fill_1 FILLER_36_2765 ();
 sg13g2_decap_4 FILLER_36_2770 ();
 sg13g2_fill_2 FILLER_36_2774 ();
 sg13g2_fill_2 FILLER_36_2781 ();
 sg13g2_decap_8 FILLER_36_2798 ();
 sg13g2_decap_8 FILLER_36_2805 ();
 sg13g2_decap_8 FILLER_36_2812 ();
 sg13g2_decap_8 FILLER_36_2889 ();
 sg13g2_decap_4 FILLER_36_2896 ();
 sg13g2_fill_2 FILLER_36_2905 ();
 sg13g2_decap_8 FILLER_36_2915 ();
 sg13g2_fill_2 FILLER_36_2922 ();
 sg13g2_fill_1 FILLER_36_2924 ();
 sg13g2_fill_2 FILLER_36_2933 ();
 sg13g2_fill_1 FILLER_36_2953 ();
 sg13g2_fill_2 FILLER_36_2962 ();
 sg13g2_fill_1 FILLER_36_2964 ();
 sg13g2_decap_8 FILLER_36_2991 ();
 sg13g2_decap_8 FILLER_36_3011 ();
 sg13g2_decap_8 FILLER_36_3018 ();
 sg13g2_fill_1 FILLER_36_3025 ();
 sg13g2_fill_2 FILLER_36_3040 ();
 sg13g2_fill_1 FILLER_36_3042 ();
 sg13g2_decap_4 FILLER_36_3061 ();
 sg13g2_fill_1 FILLER_36_3065 ();
 sg13g2_decap_8 FILLER_36_3074 ();
 sg13g2_fill_2 FILLER_36_3081 ();
 sg13g2_fill_1 FILLER_36_3083 ();
 sg13g2_decap_4 FILLER_36_3089 ();
 sg13g2_fill_2 FILLER_36_3101 ();
 sg13g2_fill_2 FILLER_36_3129 ();
 sg13g2_decap_8 FILLER_36_3135 ();
 sg13g2_fill_2 FILLER_36_3142 ();
 sg13g2_fill_2 FILLER_36_3169 ();
 sg13g2_fill_1 FILLER_36_3171 ();
 sg13g2_decap_4 FILLER_36_3193 ();
 sg13g2_fill_2 FILLER_36_3223 ();
 sg13g2_fill_1 FILLER_36_3225 ();
 sg13g2_fill_2 FILLER_36_3235 ();
 sg13g2_decap_8 FILLER_36_3266 ();
 sg13g2_decap_8 FILLER_36_3273 ();
 sg13g2_decap_4 FILLER_36_3280 ();
 sg13g2_fill_2 FILLER_36_3284 ();
 sg13g2_decap_8 FILLER_36_3290 ();
 sg13g2_decap_4 FILLER_36_3297 ();
 sg13g2_decap_4 FILLER_36_3305 ();
 sg13g2_fill_2 FILLER_36_3309 ();
 sg13g2_decap_8 FILLER_36_3337 ();
 sg13g2_decap_4 FILLER_36_3344 ();
 sg13g2_fill_2 FILLER_36_3348 ();
 sg13g2_fill_1 FILLER_36_3355 ();
 sg13g2_fill_2 FILLER_36_3365 ();
 sg13g2_decap_8 FILLER_36_3384 ();
 sg13g2_decap_8 FILLER_36_3391 ();
 sg13g2_decap_8 FILLER_36_3428 ();
 sg13g2_decap_4 FILLER_36_3435 ();
 sg13g2_fill_2 FILLER_36_3439 ();
 sg13g2_decap_8 FILLER_36_3445 ();
 sg13g2_decap_8 FILLER_36_3452 ();
 sg13g2_decap_8 FILLER_36_3459 ();
 sg13g2_decap_8 FILLER_36_3466 ();
 sg13g2_fill_2 FILLER_36_3473 ();
 sg13g2_fill_1 FILLER_36_3475 ();
 sg13g2_decap_8 FILLER_36_3489 ();
 sg13g2_decap_8 FILLER_36_3496 ();
 sg13g2_decap_8 FILLER_36_3503 ();
 sg13g2_decap_8 FILLER_36_3510 ();
 sg13g2_decap_8 FILLER_36_3517 ();
 sg13g2_decap_8 FILLER_36_3524 ();
 sg13g2_decap_8 FILLER_36_3531 ();
 sg13g2_decap_8 FILLER_36_3538 ();
 sg13g2_decap_8 FILLER_36_3545 ();
 sg13g2_decap_8 FILLER_36_3552 ();
 sg13g2_decap_8 FILLER_36_3559 ();
 sg13g2_decap_8 FILLER_36_3566 ();
 sg13g2_decap_8 FILLER_36_3573 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_4 FILLER_37_7 ();
 sg13g2_fill_1 FILLER_37_15 ();
 sg13g2_decap_4 FILLER_37_85 ();
 sg13g2_fill_2 FILLER_37_89 ();
 sg13g2_fill_2 FILLER_37_117 ();
 sg13g2_fill_1 FILLER_37_119 ();
 sg13g2_fill_1 FILLER_37_158 ();
 sg13g2_fill_1 FILLER_37_165 ();
 sg13g2_fill_1 FILLER_37_170 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_4 FILLER_37_189 ();
 sg13g2_fill_1 FILLER_37_193 ();
 sg13g2_fill_2 FILLER_37_207 ();
 sg13g2_fill_1 FILLER_37_209 ();
 sg13g2_fill_2 FILLER_37_245 ();
 sg13g2_fill_2 FILLER_37_256 ();
 sg13g2_decap_4 FILLER_37_289 ();
 sg13g2_fill_2 FILLER_37_293 ();
 sg13g2_fill_2 FILLER_37_339 ();
 sg13g2_fill_1 FILLER_37_341 ();
 sg13g2_decap_8 FILLER_37_353 ();
 sg13g2_decap_4 FILLER_37_360 ();
 sg13g2_fill_1 FILLER_37_364 ();
 sg13g2_decap_4 FILLER_37_370 ();
 sg13g2_fill_1 FILLER_37_374 ();
 sg13g2_fill_2 FILLER_37_385 ();
 sg13g2_decap_4 FILLER_37_392 ();
 sg13g2_fill_2 FILLER_37_396 ();
 sg13g2_fill_2 FILLER_37_402 ();
 sg13g2_fill_1 FILLER_37_404 ();
 sg13g2_fill_2 FILLER_37_411 ();
 sg13g2_fill_2 FILLER_37_439 ();
 sg13g2_fill_2 FILLER_37_485 ();
 sg13g2_fill_1 FILLER_37_527 ();
 sg13g2_decap_8 FILLER_37_532 ();
 sg13g2_decap_4 FILLER_37_539 ();
 sg13g2_fill_2 FILLER_37_543 ();
 sg13g2_decap_4 FILLER_37_550 ();
 sg13g2_fill_1 FILLER_37_554 ();
 sg13g2_decap_4 FILLER_37_604 ();
 sg13g2_fill_2 FILLER_37_608 ();
 sg13g2_decap_8 FILLER_37_614 ();
 sg13g2_decap_8 FILLER_37_621 ();
 sg13g2_decap_8 FILLER_37_628 ();
 sg13g2_fill_1 FILLER_37_635 ();
 sg13g2_decap_4 FILLER_37_641 ();
 sg13g2_fill_1 FILLER_37_645 ();
 sg13g2_decap_8 FILLER_37_654 ();
 sg13g2_decap_8 FILLER_37_661 ();
 sg13g2_fill_2 FILLER_37_668 ();
 sg13g2_fill_2 FILLER_37_674 ();
 sg13g2_fill_1 FILLER_37_680 ();
 sg13g2_fill_1 FILLER_37_686 ();
 sg13g2_fill_1 FILLER_37_692 ();
 sg13g2_fill_1 FILLER_37_707 ();
 sg13g2_fill_2 FILLER_37_713 ();
 sg13g2_fill_1 FILLER_37_728 ();
 sg13g2_fill_2 FILLER_37_743 ();
 sg13g2_fill_1 FILLER_37_745 ();
 sg13g2_fill_2 FILLER_37_755 ();
 sg13g2_decap_4 FILLER_37_765 ();
 sg13g2_fill_1 FILLER_37_769 ();
 sg13g2_decap_4 FILLER_37_796 ();
 sg13g2_fill_2 FILLER_37_819 ();
 sg13g2_fill_1 FILLER_37_851 ();
 sg13g2_decap_8 FILLER_37_869 ();
 sg13g2_fill_2 FILLER_37_876 ();
 sg13g2_fill_1 FILLER_37_878 ();
 sg13g2_decap_8 FILLER_37_885 ();
 sg13g2_fill_2 FILLER_37_892 ();
 sg13g2_fill_1 FILLER_37_894 ();
 sg13g2_fill_2 FILLER_37_903 ();
 sg13g2_fill_1 FILLER_37_905 ();
 sg13g2_fill_1 FILLER_37_955 ();
 sg13g2_fill_1 FILLER_37_966 ();
 sg13g2_fill_1 FILLER_37_1007 ();
 sg13g2_decap_4 FILLER_37_1034 ();
 sg13g2_fill_1 FILLER_37_1042 ();
 sg13g2_fill_1 FILLER_37_1053 ();
 sg13g2_fill_2 FILLER_37_1080 ();
 sg13g2_fill_1 FILLER_37_1082 ();
 sg13g2_fill_2 FILLER_37_1092 ();
 sg13g2_fill_2 FILLER_37_1102 ();
 sg13g2_fill_1 FILLER_37_1104 ();
 sg13g2_decap_4 FILLER_37_1109 ();
 sg13g2_decap_4 FILLER_37_1121 ();
 sg13g2_fill_2 FILLER_37_1125 ();
 sg13g2_fill_1 FILLER_37_1181 ();
 sg13g2_fill_1 FILLER_37_1208 ();
 sg13g2_fill_2 FILLER_37_1244 ();
 sg13g2_fill_1 FILLER_37_1252 ();
 sg13g2_fill_1 FILLER_37_1281 ();
 sg13g2_decap_4 FILLER_37_1294 ();
 sg13g2_decap_4 FILLER_37_1302 ();
 sg13g2_fill_1 FILLER_37_1306 ();
 sg13g2_fill_2 FILLER_37_1310 ();
 sg13g2_decap_4 FILLER_37_1320 ();
 sg13g2_decap_4 FILLER_37_1343 ();
 sg13g2_fill_2 FILLER_37_1347 ();
 sg13g2_decap_8 FILLER_37_1362 ();
 sg13g2_decap_4 FILLER_37_1369 ();
 sg13g2_fill_2 FILLER_37_1394 ();
 sg13g2_fill_1 FILLER_37_1396 ();
 sg13g2_fill_1 FILLER_37_1436 ();
 sg13g2_fill_2 FILLER_37_1444 ();
 sg13g2_fill_1 FILLER_37_1446 ();
 sg13g2_fill_1 FILLER_37_1451 ();
 sg13g2_fill_1 FILLER_37_1457 ();
 sg13g2_decap_8 FILLER_37_1462 ();
 sg13g2_decap_8 FILLER_37_1469 ();
 sg13g2_fill_2 FILLER_37_1480 ();
 sg13g2_decap_8 FILLER_37_1495 ();
 sg13g2_fill_2 FILLER_37_1502 ();
 sg13g2_fill_1 FILLER_37_1504 ();
 sg13g2_decap_4 FILLER_37_1510 ();
 sg13g2_fill_1 FILLER_37_1514 ();
 sg13g2_decap_4 FILLER_37_1535 ();
 sg13g2_decap_4 FILLER_37_1556 ();
 sg13g2_fill_1 FILLER_37_1579 ();
 sg13g2_fill_1 FILLER_37_1588 ();
 sg13g2_fill_1 FILLER_37_1613 ();
 sg13g2_fill_1 FILLER_37_1624 ();
 sg13g2_decap_8 FILLER_37_1638 ();
 sg13g2_decap_8 FILLER_37_1645 ();
 sg13g2_fill_2 FILLER_37_1656 ();
 sg13g2_decap_4 FILLER_37_1698 ();
 sg13g2_fill_1 FILLER_37_1725 ();
 sg13g2_decap_4 FILLER_37_1747 ();
 sg13g2_fill_1 FILLER_37_1757 ();
 sg13g2_fill_1 FILLER_37_1773 ();
 sg13g2_fill_2 FILLER_37_1816 ();
 sg13g2_fill_2 FILLER_37_1831 ();
 sg13g2_fill_1 FILLER_37_1844 ();
 sg13g2_decap_8 FILLER_37_1853 ();
 sg13g2_decap_4 FILLER_37_1860 ();
 sg13g2_fill_1 FILLER_37_1864 ();
 sg13g2_fill_1 FILLER_37_1903 ();
 sg13g2_fill_2 FILLER_37_1935 ();
 sg13g2_decap_4 FILLER_37_1975 ();
 sg13g2_fill_2 FILLER_37_1979 ();
 sg13g2_decap_4 FILLER_37_1986 ();
 sg13g2_fill_2 FILLER_37_1995 ();
 sg13g2_decap_8 FILLER_37_2022 ();
 sg13g2_fill_2 FILLER_37_2029 ();
 sg13g2_fill_2 FILLER_37_2071 ();
 sg13g2_decap_8 FILLER_37_2081 ();
 sg13g2_decap_4 FILLER_37_2088 ();
 sg13g2_fill_2 FILLER_37_2116 ();
 sg13g2_decap_8 FILLER_37_2124 ();
 sg13g2_decap_8 FILLER_37_2131 ();
 sg13g2_fill_2 FILLER_37_2138 ();
 sg13g2_fill_1 FILLER_37_2140 ();
 sg13g2_fill_2 FILLER_37_2155 ();
 sg13g2_decap_4 FILLER_37_2171 ();
 sg13g2_fill_1 FILLER_37_2175 ();
 sg13g2_decap_8 FILLER_37_2198 ();
 sg13g2_decap_4 FILLER_37_2205 ();
 sg13g2_fill_1 FILLER_37_2209 ();
 sg13g2_fill_2 FILLER_37_2215 ();
 sg13g2_decap_8 FILLER_37_2222 ();
 sg13g2_decap_8 FILLER_37_2229 ();
 sg13g2_fill_1 FILLER_37_2236 ();
 sg13g2_decap_8 FILLER_37_2251 ();
 sg13g2_decap_4 FILLER_37_2258 ();
 sg13g2_fill_1 FILLER_37_2262 ();
 sg13g2_decap_8 FILLER_37_2268 ();
 sg13g2_fill_2 FILLER_37_2275 ();
 sg13g2_decap_4 FILLER_37_2285 ();
 sg13g2_fill_1 FILLER_37_2289 ();
 sg13g2_decap_8 FILLER_37_2310 ();
 sg13g2_decap_4 FILLER_37_2317 ();
 sg13g2_fill_1 FILLER_37_2331 ();
 sg13g2_fill_1 FILLER_37_2350 ();
 sg13g2_decap_8 FILLER_37_2356 ();
 sg13g2_fill_1 FILLER_37_2363 ();
 sg13g2_fill_2 FILLER_37_2368 ();
 sg13g2_fill_2 FILLER_37_2379 ();
 sg13g2_decap_8 FILLER_37_2391 ();
 sg13g2_fill_1 FILLER_37_2398 ();
 sg13g2_fill_1 FILLER_37_2408 ();
 sg13g2_decap_8 FILLER_37_2427 ();
 sg13g2_fill_1 FILLER_37_2439 ();
 sg13g2_fill_2 FILLER_37_2450 ();
 sg13g2_decap_8 FILLER_37_2539 ();
 sg13g2_decap_8 FILLER_37_2546 ();
 sg13g2_decap_8 FILLER_37_2557 ();
 sg13g2_fill_2 FILLER_37_2564 ();
 sg13g2_fill_1 FILLER_37_2566 ();
 sg13g2_decap_4 FILLER_37_2574 ();
 sg13g2_fill_2 FILLER_37_2582 ();
 sg13g2_fill_1 FILLER_37_2623 ();
 sg13g2_fill_2 FILLER_37_2631 ();
 sg13g2_fill_1 FILLER_37_2633 ();
 sg13g2_fill_2 FILLER_37_2638 ();
 sg13g2_decap_8 FILLER_37_2653 ();
 sg13g2_decap_8 FILLER_37_2716 ();
 sg13g2_fill_2 FILLER_37_2723 ();
 sg13g2_fill_1 FILLER_37_2725 ();
 sg13g2_decap_4 FILLER_37_2734 ();
 sg13g2_fill_1 FILLER_37_2738 ();
 sg13g2_fill_2 FILLER_37_2753 ();
 sg13g2_fill_1 FILLER_37_2755 ();
 sg13g2_fill_1 FILLER_37_2761 ();
 sg13g2_decap_4 FILLER_37_2766 ();
 sg13g2_fill_2 FILLER_37_2779 ();
 sg13g2_fill_1 FILLER_37_2807 ();
 sg13g2_decap_8 FILLER_37_2834 ();
 sg13g2_decap_8 FILLER_37_2841 ();
 sg13g2_decap_8 FILLER_37_2848 ();
 sg13g2_decap_8 FILLER_37_2855 ();
 sg13g2_fill_2 FILLER_37_2862 ();
 sg13g2_fill_2 FILLER_37_2892 ();
 sg13g2_decap_4 FILLER_37_2920 ();
 sg13g2_fill_1 FILLER_37_2924 ();
 sg13g2_decap_4 FILLER_37_2933 ();
 sg13g2_fill_1 FILLER_37_2937 ();
 sg13g2_fill_2 FILLER_37_2953 ();
 sg13g2_fill_1 FILLER_37_2955 ();
 sg13g2_fill_2 FILLER_37_2987 ();
 sg13g2_fill_1 FILLER_37_2989 ();
 sg13g2_decap_4 FILLER_37_3011 ();
 sg13g2_fill_2 FILLER_37_3024 ();
 sg13g2_fill_1 FILLER_37_3030 ();
 sg13g2_fill_1 FILLER_37_3040 ();
 sg13g2_fill_2 FILLER_37_3062 ();
 sg13g2_fill_1 FILLER_37_3064 ();
 sg13g2_decap_4 FILLER_37_3073 ();
 sg13g2_fill_2 FILLER_37_3081 ();
 sg13g2_fill_2 FILLER_37_3118 ();
 sg13g2_fill_1 FILLER_37_3120 ();
 sg13g2_fill_1 FILLER_37_3165 ();
 sg13g2_fill_1 FILLER_37_3171 ();
 sg13g2_decap_8 FILLER_37_3177 ();
 sg13g2_decap_4 FILLER_37_3184 ();
 sg13g2_fill_2 FILLER_37_3188 ();
 sg13g2_decap_8 FILLER_37_3198 ();
 sg13g2_decap_8 FILLER_37_3205 ();
 sg13g2_fill_2 FILLER_37_3212 ();
 sg13g2_decap_4 FILLER_37_3245 ();
 sg13g2_fill_1 FILLER_37_3249 ();
 sg13g2_decap_4 FILLER_37_3271 ();
 sg13g2_decap_8 FILLER_37_3288 ();
 sg13g2_fill_2 FILLER_37_3330 ();
 sg13g2_fill_2 FILLER_37_3350 ();
 sg13g2_decap_4 FILLER_37_3378 ();
 sg13g2_decap_8 FILLER_37_3390 ();
 sg13g2_decap_8 FILLER_37_3397 ();
 sg13g2_decap_8 FILLER_37_3404 ();
 sg13g2_fill_2 FILLER_37_3411 ();
 sg13g2_decap_8 FILLER_37_3426 ();
 sg13g2_decap_8 FILLER_37_3433 ();
 sg13g2_decap_8 FILLER_37_3440 ();
 sg13g2_decap_8 FILLER_37_3447 ();
 sg13g2_decap_8 FILLER_37_3454 ();
 sg13g2_decap_8 FILLER_37_3461 ();
 sg13g2_decap_8 FILLER_37_3468 ();
 sg13g2_decap_8 FILLER_37_3475 ();
 sg13g2_decap_8 FILLER_37_3482 ();
 sg13g2_decap_8 FILLER_37_3489 ();
 sg13g2_decap_8 FILLER_37_3496 ();
 sg13g2_decap_8 FILLER_37_3503 ();
 sg13g2_decap_8 FILLER_37_3510 ();
 sg13g2_decap_8 FILLER_37_3517 ();
 sg13g2_decap_8 FILLER_37_3524 ();
 sg13g2_decap_8 FILLER_37_3531 ();
 sg13g2_decap_8 FILLER_37_3538 ();
 sg13g2_decap_8 FILLER_37_3545 ();
 sg13g2_decap_8 FILLER_37_3552 ();
 sg13g2_decap_8 FILLER_37_3559 ();
 sg13g2_decap_8 FILLER_37_3566 ();
 sg13g2_decap_8 FILLER_37_3573 ();
 sg13g2_fill_1 FILLER_38_26 ();
 sg13g2_decap_8 FILLER_38_31 ();
 sg13g2_fill_2 FILLER_38_38 ();
 sg13g2_fill_1 FILLER_38_110 ();
 sg13g2_decap_4 FILLER_38_130 ();
 sg13g2_fill_2 FILLER_38_182 ();
 sg13g2_fill_1 FILLER_38_201 ();
 sg13g2_fill_2 FILLER_38_221 ();
 sg13g2_fill_1 FILLER_38_223 ();
 sg13g2_fill_2 FILLER_38_266 ();
 sg13g2_fill_1 FILLER_38_285 ();
 sg13g2_fill_2 FILLER_38_338 ();
 sg13g2_fill_1 FILLER_38_340 ();
 sg13g2_fill_2 FILLER_38_367 ();
 sg13g2_fill_1 FILLER_38_369 ();
 sg13g2_decap_4 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_410 ();
 sg13g2_decap_4 FILLER_38_416 ();
 sg13g2_decap_4 FILLER_38_424 ();
 sg13g2_fill_2 FILLER_38_428 ();
 sg13g2_fill_2 FILLER_38_455 ();
 sg13g2_fill_1 FILLER_38_457 ();
 sg13g2_fill_2 FILLER_38_486 ();
 sg13g2_fill_2 FILLER_38_496 ();
 sg13g2_fill_2 FILLER_38_511 ();
 sg13g2_fill_1 FILLER_38_513 ();
 sg13g2_fill_2 FILLER_38_532 ();
 sg13g2_decap_4 FILLER_38_542 ();
 sg13g2_fill_1 FILLER_38_570 ();
 sg13g2_fill_2 FILLER_38_588 ();
 sg13g2_decap_4 FILLER_38_616 ();
 sg13g2_decap_8 FILLER_38_646 ();
 sg13g2_fill_2 FILLER_38_653 ();
 sg13g2_fill_1 FILLER_38_655 ();
 sg13g2_fill_2 FILLER_38_660 ();
 sg13g2_fill_1 FILLER_38_718 ();
 sg13g2_fill_2 FILLER_38_724 ();
 sg13g2_fill_1 FILLER_38_726 ();
 sg13g2_fill_1 FILLER_38_749 ();
 sg13g2_fill_2 FILLER_38_755 ();
 sg13g2_fill_1 FILLER_38_757 ();
 sg13g2_decap_8 FILLER_38_771 ();
 sg13g2_decap_8 FILLER_38_778 ();
 sg13g2_fill_1 FILLER_38_785 ();
 sg13g2_decap_8 FILLER_38_808 ();
 sg13g2_fill_1 FILLER_38_815 ();
 sg13g2_fill_2 FILLER_38_820 ();
 sg13g2_fill_1 FILLER_38_822 ();
 sg13g2_fill_1 FILLER_38_839 ();
 sg13g2_fill_1 FILLER_38_858 ();
 sg13g2_fill_1 FILLER_38_871 ();
 sg13g2_decap_4 FILLER_38_893 ();
 sg13g2_fill_2 FILLER_38_897 ();
 sg13g2_decap_8 FILLER_38_965 ();
 sg13g2_fill_1 FILLER_38_972 ();
 sg13g2_fill_2 FILLER_38_986 ();
 sg13g2_fill_1 FILLER_38_988 ();
 sg13g2_fill_2 FILLER_38_1000 ();
 sg13g2_fill_2 FILLER_38_1028 ();
 sg13g2_fill_1 FILLER_38_1030 ();
 sg13g2_decap_4 FILLER_38_1040 ();
 sg13g2_fill_1 FILLER_38_1044 ();
 sg13g2_decap_8 FILLER_38_1053 ();
 sg13g2_fill_2 FILLER_38_1080 ();
 sg13g2_decap_4 FILLER_38_1088 ();
 sg13g2_decap_4 FILLER_38_1118 ();
 sg13g2_fill_1 FILLER_38_1122 ();
 sg13g2_fill_2 FILLER_38_1127 ();
 sg13g2_fill_1 FILLER_38_1129 ();
 sg13g2_decap_8 FILLER_38_1175 ();
 sg13g2_decap_4 FILLER_38_1182 ();
 sg13g2_fill_1 FILLER_38_1186 ();
 sg13g2_decap_8 FILLER_38_1208 ();
 sg13g2_decap_8 FILLER_38_1215 ();
 sg13g2_decap_8 FILLER_38_1222 ();
 sg13g2_decap_4 FILLER_38_1229 ();
 sg13g2_fill_2 FILLER_38_1268 ();
 sg13g2_fill_1 FILLER_38_1270 ();
 sg13g2_fill_1 FILLER_38_1284 ();
 sg13g2_fill_2 FILLER_38_1298 ();
 sg13g2_fill_2 FILLER_38_1309 ();
 sg13g2_decap_8 FILLER_38_1319 ();
 sg13g2_decap_8 FILLER_38_1352 ();
 sg13g2_decap_4 FILLER_38_1359 ();
 sg13g2_decap_8 FILLER_38_1398 ();
 sg13g2_fill_2 FILLER_38_1405 ();
 sg13g2_decap_4 FILLER_38_1416 ();
 sg13g2_fill_2 FILLER_38_1420 ();
 sg13g2_fill_2 FILLER_38_1431 ();
 sg13g2_fill_1 FILLER_38_1433 ();
 sg13g2_fill_2 FILLER_38_1450 ();
 sg13g2_fill_1 FILLER_38_1452 ();
 sg13g2_fill_2 FILLER_38_1458 ();
 sg13g2_decap_4 FILLER_38_1517 ();
 sg13g2_fill_2 FILLER_38_1542 ();
 sg13g2_decap_4 FILLER_38_1549 ();
 sg13g2_fill_1 FILLER_38_1558 ();
 sg13g2_decap_8 FILLER_38_1568 ();
 sg13g2_decap_8 FILLER_38_1575 ();
 sg13g2_fill_1 FILLER_38_1587 ();
 sg13g2_decap_8 FILLER_38_1602 ();
 sg13g2_decap_8 FILLER_38_1609 ();
 sg13g2_decap_8 FILLER_38_1629 ();
 sg13g2_decap_4 FILLER_38_1636 ();
 sg13g2_fill_1 FILLER_38_1640 ();
 sg13g2_fill_2 FILLER_38_1658 ();
 sg13g2_fill_1 FILLER_38_1692 ();
 sg13g2_fill_2 FILLER_38_1699 ();
 sg13g2_decap_8 FILLER_38_1713 ();
 sg13g2_decap_4 FILLER_38_1720 ();
 sg13g2_fill_1 FILLER_38_1732 ();
 sg13g2_decap_8 FILLER_38_1738 ();
 sg13g2_decap_8 FILLER_38_1745 ();
 sg13g2_fill_2 FILLER_38_1758 ();
 sg13g2_fill_1 FILLER_38_1760 ();
 sg13g2_decap_8 FILLER_38_1766 ();
 sg13g2_decap_4 FILLER_38_1773 ();
 sg13g2_fill_2 FILLER_38_1777 ();
 sg13g2_decap_8 FILLER_38_1787 ();
 sg13g2_fill_2 FILLER_38_1794 ();
 sg13g2_decap_8 FILLER_38_1801 ();
 sg13g2_decap_8 FILLER_38_1808 ();
 sg13g2_decap_8 FILLER_38_1815 ();
 sg13g2_fill_2 FILLER_38_1822 ();
 sg13g2_fill_1 FILLER_38_1850 ();
 sg13g2_fill_2 FILLER_38_1870 ();
 sg13g2_decap_4 FILLER_38_1885 ();
 sg13g2_fill_1 FILLER_38_1923 ();
 sg13g2_fill_1 FILLER_38_1959 ();
 sg13g2_decap_4 FILLER_38_1968 ();
 sg13g2_decap_8 FILLER_38_1997 ();
 sg13g2_decap_8 FILLER_38_2004 ();
 sg13g2_fill_1 FILLER_38_2011 ();
 sg13g2_decap_8 FILLER_38_2025 ();
 sg13g2_decap_8 FILLER_38_2032 ();
 sg13g2_decap_4 FILLER_38_2039 ();
 sg13g2_fill_1 FILLER_38_2043 ();
 sg13g2_fill_1 FILLER_38_2054 ();
 sg13g2_decap_4 FILLER_38_2076 ();
 sg13g2_fill_2 FILLER_38_2094 ();
 sg13g2_fill_1 FILLER_38_2096 ();
 sg13g2_decap_4 FILLER_38_2114 ();
 sg13g2_fill_2 FILLER_38_2118 ();
 sg13g2_decap_4 FILLER_38_2131 ();
 sg13g2_fill_1 FILLER_38_2140 ();
 sg13g2_decap_8 FILLER_38_2156 ();
 sg13g2_decap_8 FILLER_38_2163 ();
 sg13g2_decap_8 FILLER_38_2170 ();
 sg13g2_decap_8 FILLER_38_2177 ();
 sg13g2_fill_2 FILLER_38_2197 ();
 sg13g2_fill_2 FILLER_38_2207 ();
 sg13g2_fill_2 FILLER_38_2232 ();
 sg13g2_decap_4 FILLER_38_2258 ();
 sg13g2_fill_1 FILLER_38_2262 ();
 sg13g2_fill_1 FILLER_38_2272 ();
 sg13g2_fill_2 FILLER_38_2278 ();
 sg13g2_fill_2 FILLER_38_2294 ();
 sg13g2_fill_1 FILLER_38_2296 ();
 sg13g2_decap_4 FILLER_38_2302 ();
 sg13g2_fill_2 FILLER_38_2306 ();
 sg13g2_fill_1 FILLER_38_2341 ();
 sg13g2_decap_4 FILLER_38_2348 ();
 sg13g2_fill_1 FILLER_38_2352 ();
 sg13g2_fill_2 FILLER_38_2357 ();
 sg13g2_fill_1 FILLER_38_2359 ();
 sg13g2_decap_8 FILLER_38_2386 ();
 sg13g2_decap_4 FILLER_38_2393 ();
 sg13g2_fill_2 FILLER_38_2397 ();
 sg13g2_decap_4 FILLER_38_2426 ();
 sg13g2_fill_1 FILLER_38_2430 ();
 sg13g2_fill_1 FILLER_38_2445 ();
 sg13g2_decap_8 FILLER_38_2499 ();
 sg13g2_fill_1 FILLER_38_2506 ();
 sg13g2_decap_4 FILLER_38_2537 ();
 sg13g2_fill_1 FILLER_38_2541 ();
 sg13g2_fill_1 FILLER_38_2594 ();
 sg13g2_fill_2 FILLER_38_2599 ();
 sg13g2_decap_4 FILLER_38_2653 ();
 sg13g2_fill_1 FILLER_38_2657 ();
 sg13g2_decap_8 FILLER_38_2662 ();
 sg13g2_decap_8 FILLER_38_2669 ();
 sg13g2_decap_8 FILLER_38_2676 ();
 sg13g2_decap_8 FILLER_38_2683 ();
 sg13g2_fill_2 FILLER_38_2690 ();
 sg13g2_fill_1 FILLER_38_2692 ();
 sg13g2_fill_2 FILLER_38_2697 ();
 sg13g2_fill_1 FILLER_38_2699 ();
 sg13g2_fill_2 FILLER_38_2705 ();
 sg13g2_fill_1 FILLER_38_2707 ();
 sg13g2_fill_2 FILLER_38_2717 ();
 sg13g2_fill_1 FILLER_38_2719 ();
 sg13g2_fill_1 FILLER_38_2777 ();
 sg13g2_decap_8 FILLER_38_2798 ();
 sg13g2_decap_8 FILLER_38_2805 ();
 sg13g2_fill_2 FILLER_38_2812 ();
 sg13g2_fill_1 FILLER_38_2818 ();
 sg13g2_fill_1 FILLER_38_2848 ();
 sg13g2_fill_1 FILLER_38_2854 ();
 sg13g2_fill_2 FILLER_38_2863 ();
 sg13g2_fill_1 FILLER_38_2865 ();
 sg13g2_decap_8 FILLER_38_2891 ();
 sg13g2_fill_2 FILLER_38_2914 ();
 sg13g2_fill_1 FILLER_38_2916 ();
 sg13g2_decap_4 FILLER_38_2925 ();
 sg13g2_fill_2 FILLER_38_2929 ();
 sg13g2_decap_8 FILLER_38_2962 ();
 sg13g2_fill_2 FILLER_38_2969 ();
 sg13g2_fill_1 FILLER_38_2971 ();
 sg13g2_decap_4 FILLER_38_2976 ();
 sg13g2_fill_2 FILLER_38_2984 ();
 sg13g2_fill_1 FILLER_38_2986 ();
 sg13g2_fill_1 FILLER_38_2992 ();
 sg13g2_decap_4 FILLER_38_3010 ();
 sg13g2_fill_1 FILLER_38_3014 ();
 sg13g2_fill_2 FILLER_38_3045 ();
 sg13g2_decap_8 FILLER_38_3055 ();
 sg13g2_decap_8 FILLER_38_3062 ();
 sg13g2_fill_2 FILLER_38_3069 ();
 sg13g2_decap_4 FILLER_38_3106 ();
 sg13g2_fill_1 FILLER_38_3110 ();
 sg13g2_fill_2 FILLER_38_3125 ();
 sg13g2_fill_2 FILLER_38_3154 ();
 sg13g2_fill_1 FILLER_38_3156 ();
 sg13g2_fill_2 FILLER_38_3191 ();
 sg13g2_fill_2 FILLER_38_3214 ();
 sg13g2_decap_8 FILLER_38_3229 ();
 sg13g2_fill_2 FILLER_38_3236 ();
 sg13g2_fill_1 FILLER_38_3238 ();
 sg13g2_fill_1 FILLER_38_3309 ();
 sg13g2_decap_8 FILLER_38_3359 ();
 sg13g2_decap_8 FILLER_38_3366 ();
 sg13g2_decap_8 FILLER_38_3373 ();
 sg13g2_decap_8 FILLER_38_3380 ();
 sg13g2_decap_8 FILLER_38_3387 ();
 sg13g2_decap_8 FILLER_38_3394 ();
 sg13g2_decap_8 FILLER_38_3401 ();
 sg13g2_decap_8 FILLER_38_3408 ();
 sg13g2_decap_8 FILLER_38_3415 ();
 sg13g2_decap_8 FILLER_38_3422 ();
 sg13g2_decap_8 FILLER_38_3429 ();
 sg13g2_decap_8 FILLER_38_3436 ();
 sg13g2_decap_8 FILLER_38_3443 ();
 sg13g2_decap_8 FILLER_38_3450 ();
 sg13g2_decap_8 FILLER_38_3457 ();
 sg13g2_decap_8 FILLER_38_3464 ();
 sg13g2_decap_8 FILLER_38_3471 ();
 sg13g2_decap_8 FILLER_38_3478 ();
 sg13g2_decap_8 FILLER_38_3485 ();
 sg13g2_decap_8 FILLER_38_3492 ();
 sg13g2_decap_8 FILLER_38_3499 ();
 sg13g2_decap_8 FILLER_38_3506 ();
 sg13g2_decap_8 FILLER_38_3513 ();
 sg13g2_decap_8 FILLER_38_3520 ();
 sg13g2_decap_8 FILLER_38_3527 ();
 sg13g2_decap_8 FILLER_38_3534 ();
 sg13g2_decap_8 FILLER_38_3541 ();
 sg13g2_decap_8 FILLER_38_3548 ();
 sg13g2_decap_8 FILLER_38_3555 ();
 sg13g2_decap_8 FILLER_38_3562 ();
 sg13g2_decap_8 FILLER_38_3569 ();
 sg13g2_decap_4 FILLER_38_3576 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_39_7 ();
 sg13g2_fill_2 FILLER_39_35 ();
 sg13g2_fill_1 FILLER_39_37 ();
 sg13g2_fill_2 FILLER_39_47 ();
 sg13g2_fill_1 FILLER_39_49 ();
 sg13g2_fill_1 FILLER_39_59 ();
 sg13g2_fill_2 FILLER_39_63 ();
 sg13g2_fill_1 FILLER_39_65 ();
 sg13g2_decap_4 FILLER_39_78 ();
 sg13g2_decap_8 FILLER_39_86 ();
 sg13g2_decap_8 FILLER_39_93 ();
 sg13g2_fill_2 FILLER_39_100 ();
 sg13g2_fill_1 FILLER_39_102 ();
 sg13g2_decap_4 FILLER_39_107 ();
 sg13g2_decap_8 FILLER_39_118 ();
 sg13g2_fill_1 FILLER_39_125 ();
 sg13g2_fill_1 FILLER_39_160 ();
 sg13g2_decap_8 FILLER_39_166 ();
 sg13g2_decap_8 FILLER_39_173 ();
 sg13g2_decap_8 FILLER_39_184 ();
 sg13g2_fill_1 FILLER_39_191 ();
 sg13g2_fill_2 FILLER_39_202 ();
 sg13g2_fill_2 FILLER_39_238 ();
 sg13g2_fill_1 FILLER_39_240 ();
 sg13g2_decap_8 FILLER_39_253 ();
 sg13g2_decap_4 FILLER_39_260 ();
 sg13g2_decap_8 FILLER_39_282 ();
 sg13g2_decap_8 FILLER_39_289 ();
 sg13g2_fill_2 FILLER_39_296 ();
 sg13g2_fill_2 FILLER_39_302 ();
 sg13g2_fill_1 FILLER_39_304 ();
 sg13g2_decap_8 FILLER_39_310 ();
 sg13g2_decap_4 FILLER_39_317 ();
 sg13g2_fill_2 FILLER_39_321 ();
 sg13g2_decap_4 FILLER_39_336 ();
 sg13g2_fill_1 FILLER_39_340 ();
 sg13g2_decap_8 FILLER_39_364 ();
 sg13g2_fill_2 FILLER_39_371 ();
 sg13g2_fill_1 FILLER_39_373 ();
 sg13g2_fill_1 FILLER_39_379 ();
 sg13g2_fill_2 FILLER_39_384 ();
 sg13g2_fill_1 FILLER_39_386 ();
 sg13g2_decap_8 FILLER_39_396 ();
 sg13g2_decap_4 FILLER_39_403 ();
 sg13g2_fill_1 FILLER_39_407 ();
 sg13g2_decap_4 FILLER_39_416 ();
 sg13g2_decap_4 FILLER_39_432 ();
 sg13g2_fill_2 FILLER_39_455 ();
 sg13g2_fill_1 FILLER_39_457 ();
 sg13g2_decap_4 FILLER_39_502 ();
 sg13g2_fill_2 FILLER_39_518 ();
 sg13g2_decap_8 FILLER_39_553 ();
 sg13g2_fill_2 FILLER_39_568 ();
 sg13g2_decap_4 FILLER_39_580 ();
 sg13g2_decap_4 FILLER_39_598 ();
 sg13g2_decap_8 FILLER_39_620 ();
 sg13g2_decap_8 FILLER_39_637 ();
 sg13g2_fill_2 FILLER_39_644 ();
 sg13g2_fill_2 FILLER_39_672 ();
 sg13g2_fill_2 FILLER_39_683 ();
 sg13g2_fill_1 FILLER_39_685 ();
 sg13g2_fill_2 FILLER_39_694 ();
 sg13g2_decap_4 FILLER_39_714 ();
 sg13g2_fill_2 FILLER_39_718 ();
 sg13g2_fill_2 FILLER_39_724 ();
 sg13g2_fill_1 FILLER_39_726 ();
 sg13g2_fill_2 FILLER_39_741 ();
 sg13g2_fill_1 FILLER_39_743 ();
 sg13g2_decap_4 FILLER_39_754 ();
 sg13g2_fill_2 FILLER_39_815 ();
 sg13g2_fill_1 FILLER_39_817 ();
 sg13g2_fill_1 FILLER_39_823 ();
 sg13g2_fill_2 FILLER_39_845 ();
 sg13g2_fill_1 FILLER_39_857 ();
 sg13g2_fill_2 FILLER_39_861 ();
 sg13g2_fill_2 FILLER_39_871 ();
 sg13g2_decap_8 FILLER_39_888 ();
 sg13g2_decap_8 FILLER_39_895 ();
 sg13g2_decap_8 FILLER_39_902 ();
 sg13g2_fill_1 FILLER_39_909 ();
 sg13g2_fill_2 FILLER_39_924 ();
 sg13g2_fill_2 FILLER_39_970 ();
 sg13g2_fill_1 FILLER_39_1019 ();
 sg13g2_decap_4 FILLER_39_1072 ();
 sg13g2_decap_4 FILLER_39_1090 ();
 sg13g2_fill_2 FILLER_39_1094 ();
 sg13g2_fill_1 FILLER_39_1116 ();
 sg13g2_fill_1 FILLER_39_1126 ();
 sg13g2_fill_2 FILLER_39_1148 ();
 sg13g2_fill_1 FILLER_39_1150 ();
 sg13g2_decap_4 FILLER_39_1199 ();
 sg13g2_fill_2 FILLER_39_1203 ();
 sg13g2_decap_4 FILLER_39_1240 ();
 sg13g2_decap_4 FILLER_39_1248 ();
 sg13g2_fill_1 FILLER_39_1260 ();
 sg13g2_fill_2 FILLER_39_1266 ();
 sg13g2_fill_2 FILLER_39_1277 ();
 sg13g2_fill_1 FILLER_39_1279 ();
 sg13g2_fill_1 FILLER_39_1311 ();
 sg13g2_fill_2 FILLER_39_1327 ();
 sg13g2_fill_1 FILLER_39_1329 ();
 sg13g2_fill_1 FILLER_39_1334 ();
 sg13g2_decap_8 FILLER_39_1347 ();
 sg13g2_decap_8 FILLER_39_1372 ();
 sg13g2_decap_8 FILLER_39_1379 ();
 sg13g2_decap_8 FILLER_39_1386 ();
 sg13g2_fill_1 FILLER_39_1393 ();
 sg13g2_decap_8 FILLER_39_1403 ();
 sg13g2_decap_8 FILLER_39_1410 ();
 sg13g2_decap_4 FILLER_39_1417 ();
 sg13g2_fill_1 FILLER_39_1421 ();
 sg13g2_decap_4 FILLER_39_1430 ();
 sg13g2_fill_1 FILLER_39_1434 ();
 sg13g2_decap_8 FILLER_39_1440 ();
 sg13g2_decap_8 FILLER_39_1447 ();
 sg13g2_fill_1 FILLER_39_1459 ();
 sg13g2_decap_4 FILLER_39_1470 ();
 sg13g2_fill_2 FILLER_39_1474 ();
 sg13g2_fill_2 FILLER_39_1504 ();
 sg13g2_fill_1 FILLER_39_1506 ();
 sg13g2_decap_8 FILLER_39_1519 ();
 sg13g2_fill_1 FILLER_39_1526 ();
 sg13g2_decap_8 FILLER_39_1540 ();
 sg13g2_decap_8 FILLER_39_1547 ();
 sg13g2_fill_1 FILLER_39_1554 ();
 sg13g2_fill_2 FILLER_39_1573 ();
 sg13g2_fill_1 FILLER_39_1575 ();
 sg13g2_decap_4 FILLER_39_1580 ();
 sg13g2_fill_1 FILLER_39_1584 ();
 sg13g2_decap_8 FILLER_39_1588 ();
 sg13g2_decap_4 FILLER_39_1595 ();
 sg13g2_fill_1 FILLER_39_1599 ();
 sg13g2_decap_4 FILLER_39_1610 ();
 sg13g2_fill_2 FILLER_39_1654 ();
 sg13g2_fill_2 FILLER_39_1661 ();
 sg13g2_fill_1 FILLER_39_1663 ();
 sg13g2_fill_2 FILLER_39_1669 ();
 sg13g2_fill_1 FILLER_39_1671 ();
 sg13g2_decap_8 FILLER_39_1684 ();
 sg13g2_decap_4 FILLER_39_1691 ();
 sg13g2_fill_1 FILLER_39_1695 ();
 sg13g2_fill_1 FILLER_39_1700 ();
 sg13g2_decap_8 FILLER_39_1706 ();
 sg13g2_fill_2 FILLER_39_1713 ();
 sg13g2_fill_1 FILLER_39_1715 ();
 sg13g2_decap_8 FILLER_39_1739 ();
 sg13g2_fill_2 FILLER_39_1746 ();
 sg13g2_fill_1 FILLER_39_1748 ();
 sg13g2_decap_8 FILLER_39_1760 ();
 sg13g2_decap_8 FILLER_39_1767 ();
 sg13g2_decap_8 FILLER_39_1795 ();
 sg13g2_fill_2 FILLER_39_1816 ();
 sg13g2_fill_1 FILLER_39_1818 ();
 sg13g2_decap_8 FILLER_39_1854 ();
 sg13g2_decap_8 FILLER_39_1861 ();
 sg13g2_fill_2 FILLER_39_1874 ();
 sg13g2_decap_8 FILLER_39_1884 ();
 sg13g2_decap_8 FILLER_39_1896 ();
 sg13g2_fill_2 FILLER_39_1907 ();
 sg13g2_fill_1 FILLER_39_1909 ();
 sg13g2_fill_1 FILLER_39_1921 ();
 sg13g2_decap_4 FILLER_39_1933 ();
 sg13g2_decap_4 FILLER_39_1942 ();
 sg13g2_fill_2 FILLER_39_1946 ();
 sg13g2_decap_8 FILLER_39_1955 ();
 sg13g2_decap_4 FILLER_39_1962 ();
 sg13g2_fill_1 FILLER_39_1966 ();
 sg13g2_decap_4 FILLER_39_1987 ();
 sg13g2_fill_1 FILLER_39_1999 ();
 sg13g2_fill_1 FILLER_39_2032 ();
 sg13g2_fill_2 FILLER_39_2043 ();
 sg13g2_decap_4 FILLER_39_2068 ();
 sg13g2_fill_2 FILLER_39_2072 ();
 sg13g2_decap_8 FILLER_39_2082 ();
 sg13g2_fill_2 FILLER_39_2089 ();
 sg13g2_decap_8 FILLER_39_2096 ();
 sg13g2_fill_2 FILLER_39_2103 ();
 sg13g2_decap_4 FILLER_39_2163 ();
 sg13g2_fill_1 FILLER_39_2167 ();
 sg13g2_fill_1 FILLER_39_2176 ();
 sg13g2_fill_1 FILLER_39_2189 ();
 sg13g2_decap_8 FILLER_39_2203 ();
 sg13g2_decap_4 FILLER_39_2210 ();
 sg13g2_decap_4 FILLER_39_2224 ();
 sg13g2_fill_1 FILLER_39_2228 ();
 sg13g2_fill_2 FILLER_39_2238 ();
 sg13g2_fill_1 FILLER_39_2240 ();
 sg13g2_fill_2 FILLER_39_2246 ();
 sg13g2_decap_4 FILLER_39_2262 ();
 sg13g2_fill_1 FILLER_39_2266 ();
 sg13g2_decap_8 FILLER_39_2275 ();
 sg13g2_fill_2 FILLER_39_2282 ();
 sg13g2_fill_1 FILLER_39_2284 ();
 sg13g2_decap_8 FILLER_39_2290 ();
 sg13g2_decap_4 FILLER_39_2297 ();
 sg13g2_decap_8 FILLER_39_2309 ();
 sg13g2_fill_1 FILLER_39_2316 ();
 sg13g2_decap_8 FILLER_39_2331 ();
 sg13g2_fill_2 FILLER_39_2338 ();
 sg13g2_fill_1 FILLER_39_2340 ();
 sg13g2_fill_2 FILLER_39_2380 ();
 sg13g2_decap_8 FILLER_39_2387 ();
 sg13g2_fill_1 FILLER_39_2394 ();
 sg13g2_decap_4 FILLER_39_2421 ();
 sg13g2_fill_2 FILLER_39_2445 ();
 sg13g2_fill_1 FILLER_39_2447 ();
 sg13g2_fill_2 FILLER_39_2466 ();
 sg13g2_fill_1 FILLER_39_2468 ();
 sg13g2_decap_8 FILLER_39_2535 ();
 sg13g2_fill_2 FILLER_39_2542 ();
 sg13g2_fill_2 FILLER_39_2561 ();
 sg13g2_fill_1 FILLER_39_2563 ();
 sg13g2_fill_2 FILLER_39_2571 ();
 sg13g2_fill_2 FILLER_39_2600 ();
 sg13g2_fill_2 FILLER_39_2614 ();
 sg13g2_decap_8 FILLER_39_2633 ();
 sg13g2_decap_8 FILLER_39_2640 ();
 sg13g2_decap_4 FILLER_39_2673 ();
 sg13g2_fill_1 FILLER_39_2677 ();
 sg13g2_fill_2 FILLER_39_2735 ();
 sg13g2_decap_8 FILLER_39_2749 ();
 sg13g2_fill_2 FILLER_39_2756 ();
 sg13g2_fill_1 FILLER_39_2758 ();
 sg13g2_decap_8 FILLER_39_2763 ();
 sg13g2_decap_4 FILLER_39_2770 ();
 sg13g2_fill_2 FILLER_39_2774 ();
 sg13g2_decap_8 FILLER_39_2797 ();
 sg13g2_decap_4 FILLER_39_2804 ();
 sg13g2_decap_4 FILLER_39_2839 ();
 sg13g2_fill_1 FILLER_39_2843 ();
 sg13g2_decap_8 FILLER_39_2885 ();
 sg13g2_decap_4 FILLER_39_2892 ();
 sg13g2_fill_1 FILLER_39_2905 ();
 sg13g2_decap_8 FILLER_39_2932 ();
 sg13g2_decap_4 FILLER_39_2939 ();
 sg13g2_fill_1 FILLER_39_2943 ();
 sg13g2_decap_8 FILLER_39_2969 ();
 sg13g2_fill_2 FILLER_39_2976 ();
 sg13g2_fill_1 FILLER_39_2978 ();
 sg13g2_decap_4 FILLER_39_3023 ();
 sg13g2_fill_1 FILLER_39_3041 ();
 sg13g2_fill_1 FILLER_39_3056 ();
 sg13g2_fill_2 FILLER_39_3061 ();
 sg13g2_decap_4 FILLER_39_3071 ();
 sg13g2_fill_1 FILLER_39_3084 ();
 sg13g2_fill_2 FILLER_39_3107 ();
 sg13g2_decap_8 FILLER_39_3161 ();
 sg13g2_decap_4 FILLER_39_3168 ();
 sg13g2_decap_8 FILLER_39_3179 ();
 sg13g2_decap_4 FILLER_39_3186 ();
 sg13g2_decap_8 FILLER_39_3198 ();
 sg13g2_fill_2 FILLER_39_3205 ();
 sg13g2_fill_1 FILLER_39_3207 ();
 sg13g2_fill_2 FILLER_39_3253 ();
 sg13g2_fill_1 FILLER_39_3255 ();
 sg13g2_decap_4 FILLER_39_3274 ();
 sg13g2_fill_2 FILLER_39_3278 ();
 sg13g2_fill_1 FILLER_39_3289 ();
 sg13g2_decap_8 FILLER_39_3295 ();
 sg13g2_decap_4 FILLER_39_3302 ();
 sg13g2_fill_2 FILLER_39_3315 ();
 sg13g2_fill_1 FILLER_39_3317 ();
 sg13g2_decap_8 FILLER_39_3344 ();
 sg13g2_decap_8 FILLER_39_3351 ();
 sg13g2_decap_8 FILLER_39_3358 ();
 sg13g2_decap_8 FILLER_39_3365 ();
 sg13g2_decap_8 FILLER_39_3372 ();
 sg13g2_decap_8 FILLER_39_3379 ();
 sg13g2_decap_8 FILLER_39_3386 ();
 sg13g2_decap_8 FILLER_39_3393 ();
 sg13g2_decap_8 FILLER_39_3400 ();
 sg13g2_decap_8 FILLER_39_3407 ();
 sg13g2_decap_8 FILLER_39_3414 ();
 sg13g2_decap_8 FILLER_39_3421 ();
 sg13g2_decap_8 FILLER_39_3428 ();
 sg13g2_decap_8 FILLER_39_3435 ();
 sg13g2_decap_8 FILLER_39_3442 ();
 sg13g2_decap_8 FILLER_39_3449 ();
 sg13g2_decap_8 FILLER_39_3456 ();
 sg13g2_decap_8 FILLER_39_3463 ();
 sg13g2_decap_8 FILLER_39_3470 ();
 sg13g2_decap_8 FILLER_39_3477 ();
 sg13g2_decap_8 FILLER_39_3484 ();
 sg13g2_decap_8 FILLER_39_3491 ();
 sg13g2_decap_8 FILLER_39_3498 ();
 sg13g2_decap_8 FILLER_39_3505 ();
 sg13g2_decap_8 FILLER_39_3512 ();
 sg13g2_decap_8 FILLER_39_3519 ();
 sg13g2_decap_8 FILLER_39_3526 ();
 sg13g2_decap_8 FILLER_39_3533 ();
 sg13g2_decap_8 FILLER_39_3540 ();
 sg13g2_decap_8 FILLER_39_3547 ();
 sg13g2_decap_8 FILLER_39_3554 ();
 sg13g2_decap_8 FILLER_39_3561 ();
 sg13g2_decap_8 FILLER_39_3568 ();
 sg13g2_decap_4 FILLER_39_3575 ();
 sg13g2_fill_1 FILLER_39_3579 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_4 FILLER_40_7 ();
 sg13g2_fill_2 FILLER_40_15 ();
 sg13g2_fill_2 FILLER_40_44 ();
 sg13g2_fill_1 FILLER_40_46 ();
 sg13g2_decap_8 FILLER_40_79 ();
 sg13g2_decap_4 FILLER_40_86 ();
 sg13g2_fill_2 FILLER_40_90 ();
 sg13g2_fill_2 FILLER_40_118 ();
 sg13g2_fill_1 FILLER_40_165 ();
 sg13g2_decap_4 FILLER_40_228 ();
 sg13g2_fill_1 FILLER_40_241 ();
 sg13g2_fill_1 FILLER_40_246 ();
 sg13g2_fill_1 FILLER_40_256 ();
 sg13g2_decap_8 FILLER_40_267 ();
 sg13g2_decap_4 FILLER_40_274 ();
 sg13g2_fill_2 FILLER_40_294 ();
 sg13g2_fill_1 FILLER_40_296 ();
 sg13g2_fill_2 FILLER_40_321 ();
 sg13g2_decap_4 FILLER_40_349 ();
 sg13g2_fill_1 FILLER_40_353 ();
 sg13g2_fill_1 FILLER_40_362 ();
 sg13g2_decap_8 FILLER_40_369 ();
 sg13g2_fill_2 FILLER_40_376 ();
 sg13g2_fill_1 FILLER_40_378 ();
 sg13g2_fill_2 FILLER_40_383 ();
 sg13g2_fill_1 FILLER_40_385 ();
 sg13g2_decap_8 FILLER_40_402 ();
 sg13g2_fill_1 FILLER_40_409 ();
 sg13g2_decap_8 FILLER_40_447 ();
 sg13g2_decap_8 FILLER_40_454 ();
 sg13g2_decap_4 FILLER_40_461 ();
 sg13g2_fill_1 FILLER_40_465 ();
 sg13g2_fill_1 FILLER_40_480 ();
 sg13g2_decap_8 FILLER_40_490 ();
 sg13g2_decap_8 FILLER_40_497 ();
 sg13g2_decap_8 FILLER_40_504 ();
 sg13g2_decap_8 FILLER_40_511 ();
 sg13g2_decap_4 FILLER_40_518 ();
 sg13g2_decap_4 FILLER_40_538 ();
 sg13g2_decap_4 FILLER_40_586 ();
 sg13g2_fill_1 FILLER_40_594 ();
 sg13g2_fill_1 FILLER_40_613 ();
 sg13g2_decap_8 FILLER_40_619 ();
 sg13g2_decap_8 FILLER_40_630 ();
 sg13g2_decap_4 FILLER_40_642 ();
 sg13g2_decap_4 FILLER_40_669 ();
 sg13g2_decap_4 FILLER_40_703 ();
 sg13g2_fill_2 FILLER_40_707 ();
 sg13g2_decap_4 FILLER_40_745 ();
 sg13g2_fill_1 FILLER_40_749 ();
 sg13g2_fill_2 FILLER_40_760 ();
 sg13g2_fill_1 FILLER_40_762 ();
 sg13g2_decap_8 FILLER_40_769 ();
 sg13g2_decap_4 FILLER_40_780 ();
 sg13g2_fill_2 FILLER_40_788 ();
 sg13g2_fill_1 FILLER_40_790 ();
 sg13g2_decap_8 FILLER_40_795 ();
 sg13g2_fill_2 FILLER_40_802 ();
 sg13g2_fill_1 FILLER_40_804 ();
 sg13g2_fill_2 FILLER_40_813 ();
 sg13g2_fill_1 FILLER_40_823 ();
 sg13g2_fill_1 FILLER_40_834 ();
 sg13g2_fill_1 FILLER_40_874 ();
 sg13g2_decap_4 FILLER_40_894 ();
 sg13g2_fill_1 FILLER_40_898 ();
 sg13g2_fill_2 FILLER_40_938 ();
 sg13g2_fill_2 FILLER_40_967 ();
 sg13g2_fill_1 FILLER_40_969 ();
 sg13g2_decap_8 FILLER_40_1004 ();
 sg13g2_fill_2 FILLER_40_1011 ();
 sg13g2_fill_2 FILLER_40_1020 ();
 sg13g2_fill_1 FILLER_40_1022 ();
 sg13g2_decap_8 FILLER_40_1036 ();
 sg13g2_decap_8 FILLER_40_1043 ();
 sg13g2_fill_1 FILLER_40_1050 ();
 sg13g2_fill_2 FILLER_40_1055 ();
 sg13g2_fill_2 FILLER_40_1061 ();
 sg13g2_fill_2 FILLER_40_1072 ();
 sg13g2_decap_4 FILLER_40_1084 ();
 sg13g2_decap_8 FILLER_40_1093 ();
 sg13g2_fill_2 FILLER_40_1100 ();
 sg13g2_fill_1 FILLER_40_1102 ();
 sg13g2_fill_2 FILLER_40_1114 ();
 sg13g2_decap_8 FILLER_40_1126 ();
 sg13g2_decap_8 FILLER_40_1133 ();
 sg13g2_fill_2 FILLER_40_1140 ();
 sg13g2_fill_1 FILLER_40_1142 ();
 sg13g2_decap_8 FILLER_40_1149 ();
 sg13g2_fill_1 FILLER_40_1156 ();
 sg13g2_fill_2 FILLER_40_1171 ();
 sg13g2_fill_1 FILLER_40_1173 ();
 sg13g2_fill_1 FILLER_40_1182 ();
 sg13g2_fill_2 FILLER_40_1189 ();
 sg13g2_fill_2 FILLER_40_1208 ();
 sg13g2_fill_1 FILLER_40_1220 ();
 sg13g2_decap_4 FILLER_40_1284 ();
 sg13g2_fill_2 FILLER_40_1288 ();
 sg13g2_decap_4 FILLER_40_1298 ();
 sg13g2_decap_8 FILLER_40_1306 ();
 sg13g2_fill_2 FILLER_40_1313 ();
 sg13g2_fill_1 FILLER_40_1315 ();
 sg13g2_decap_4 FILLER_40_1348 ();
 sg13g2_fill_2 FILLER_40_1368 ();
 sg13g2_fill_1 FILLER_40_1370 ();
 sg13g2_fill_2 FILLER_40_1377 ();
 sg13g2_fill_1 FILLER_40_1389 ();
 sg13g2_fill_2 FILLER_40_1418 ();
 sg13g2_fill_1 FILLER_40_1420 ();
 sg13g2_fill_1 FILLER_40_1434 ();
 sg13g2_decap_4 FILLER_40_1445 ();
 sg13g2_fill_1 FILLER_40_1449 ();
 sg13g2_fill_2 FILLER_40_1485 ();
 sg13g2_fill_1 FILLER_40_1487 ();
 sg13g2_fill_2 FILLER_40_1498 ();
 sg13g2_fill_2 FILLER_40_1536 ();
 sg13g2_fill_1 FILLER_40_1551 ();
 sg13g2_fill_1 FILLER_40_1587 ();
 sg13g2_fill_1 FILLER_40_1632 ();
 sg13g2_fill_2 FILLER_40_1658 ();
 sg13g2_fill_1 FILLER_40_1660 ();
 sg13g2_fill_1 FILLER_40_1667 ();
 sg13g2_decap_4 FILLER_40_1676 ();
 sg13g2_fill_1 FILLER_40_1695 ();
 sg13g2_decap_8 FILLER_40_1716 ();
 sg13g2_fill_2 FILLER_40_1723 ();
 sg13g2_decap_8 FILLER_40_1737 ();
 sg13g2_fill_1 FILLER_40_1744 ();
 sg13g2_fill_1 FILLER_40_1767 ();
 sg13g2_fill_1 FILLER_40_1806 ();
 sg13g2_fill_1 FILLER_40_1815 ();
 sg13g2_fill_2 FILLER_40_1838 ();
 sg13g2_fill_1 FILLER_40_1851 ();
 sg13g2_fill_2 FILLER_40_1857 ();
 sg13g2_fill_1 FILLER_40_1862 ();
 sg13g2_fill_2 FILLER_40_1898 ();
 sg13g2_decap_8 FILLER_40_1926 ();
 sg13g2_fill_2 FILLER_40_1933 ();
 sg13g2_fill_1 FILLER_40_1935 ();
 sg13g2_fill_2 FILLER_40_1946 ();
 sg13g2_fill_1 FILLER_40_1948 ();
 sg13g2_decap_8 FILLER_40_1957 ();
 sg13g2_fill_2 FILLER_40_1964 ();
 sg13g2_fill_1 FILLER_40_1966 ();
 sg13g2_decap_8 FILLER_40_1982 ();
 sg13g2_decap_8 FILLER_40_1989 ();
 sg13g2_fill_2 FILLER_40_1996 ();
 sg13g2_fill_1 FILLER_40_1998 ();
 sg13g2_fill_2 FILLER_40_2019 ();
 sg13g2_decap_4 FILLER_40_2027 ();
 sg13g2_fill_1 FILLER_40_2039 ();
 sg13g2_decap_8 FILLER_40_2048 ();
 sg13g2_fill_2 FILLER_40_2055 ();
 sg13g2_decap_8 FILLER_40_2068 ();
 sg13g2_fill_1 FILLER_40_2075 ();
 sg13g2_fill_1 FILLER_40_2090 ();
 sg13g2_decap_8 FILLER_40_2102 ();
 sg13g2_decap_8 FILLER_40_2119 ();
 sg13g2_fill_2 FILLER_40_2126 ();
 sg13g2_decap_8 FILLER_40_2137 ();
 sg13g2_decap_4 FILLER_40_2144 ();
 sg13g2_fill_1 FILLER_40_2148 ();
 sg13g2_decap_8 FILLER_40_2157 ();
 sg13g2_fill_2 FILLER_40_2164 ();
 sg13g2_decap_8 FILLER_40_2174 ();
 sg13g2_fill_2 FILLER_40_2208 ();
 sg13g2_fill_1 FILLER_40_2210 ();
 sg13g2_decap_8 FILLER_40_2230 ();
 sg13g2_decap_4 FILLER_40_2237 ();
 sg13g2_decap_8 FILLER_40_2250 ();
 sg13g2_decap_4 FILLER_40_2257 ();
 sg13g2_fill_2 FILLER_40_2266 ();
 sg13g2_fill_1 FILLER_40_2268 ();
 sg13g2_decap_8 FILLER_40_2279 ();
 sg13g2_decap_4 FILLER_40_2286 ();
 sg13g2_fill_1 FILLER_40_2290 ();
 sg13g2_fill_2 FILLER_40_2322 ();
 sg13g2_decap_8 FILLER_40_2339 ();
 sg13g2_fill_2 FILLER_40_2346 ();
 sg13g2_fill_2 FILLER_40_2358 ();
 sg13g2_decap_8 FILLER_40_2409 ();
 sg13g2_decap_8 FILLER_40_2416 ();
 sg13g2_decap_8 FILLER_40_2423 ();
 sg13g2_fill_2 FILLER_40_2430 ();
 sg13g2_fill_1 FILLER_40_2432 ();
 sg13g2_fill_2 FILLER_40_2486 ();
 sg13g2_fill_1 FILLER_40_2488 ();
 sg13g2_fill_2 FILLER_40_2494 ();
 sg13g2_fill_1 FILLER_40_2496 ();
 sg13g2_fill_2 FILLER_40_2501 ();
 sg13g2_fill_1 FILLER_40_2503 ();
 sg13g2_decap_4 FILLER_40_2535 ();
 sg13g2_fill_2 FILLER_40_2544 ();
 sg13g2_fill_1 FILLER_40_2546 ();
 sg13g2_fill_2 FILLER_40_2559 ();
 sg13g2_fill_1 FILLER_40_2561 ();
 sg13g2_decap_8 FILLER_40_2665 ();
 sg13g2_decap_8 FILLER_40_2672 ();
 sg13g2_decap_8 FILLER_40_2679 ();
 sg13g2_fill_2 FILLER_40_2686 ();
 sg13g2_fill_2 FILLER_40_2701 ();
 sg13g2_decap_8 FILLER_40_2707 ();
 sg13g2_decap_8 FILLER_40_2718 ();
 sg13g2_decap_8 FILLER_40_2725 ();
 sg13g2_fill_1 FILLER_40_2732 ();
 sg13g2_fill_2 FILLER_40_2751 ();
 sg13g2_fill_1 FILLER_40_2753 ();
 sg13g2_decap_4 FILLER_40_2798 ();
 sg13g2_fill_2 FILLER_40_2802 ();
 sg13g2_decap_8 FILLER_40_2834 ();
 sg13g2_decap_8 FILLER_40_2841 ();
 sg13g2_fill_1 FILLER_40_2848 ();
 sg13g2_fill_2 FILLER_40_2854 ();
 sg13g2_decap_4 FILLER_40_2865 ();
 sg13g2_decap_4 FILLER_40_2887 ();
 sg13g2_decap_8 FILLER_40_2904 ();
 sg13g2_decap_4 FILLER_40_2911 ();
 sg13g2_decap_8 FILLER_40_2928 ();
 sg13g2_fill_1 FILLER_40_2935 ();
 sg13g2_decap_8 FILLER_40_2975 ();
 sg13g2_decap_4 FILLER_40_2982 ();
 sg13g2_fill_1 FILLER_40_2986 ();
 sg13g2_decap_4 FILLER_40_3013 ();
 sg13g2_fill_2 FILLER_40_3043 ();
 sg13g2_fill_1 FILLER_40_3045 ();
 sg13g2_fill_1 FILLER_40_3081 ();
 sg13g2_fill_2 FILLER_40_3117 ();
 sg13g2_fill_1 FILLER_40_3119 ();
 sg13g2_decap_8 FILLER_40_3124 ();
 sg13g2_decap_4 FILLER_40_3131 ();
 sg13g2_fill_2 FILLER_40_3135 ();
 sg13g2_fill_2 FILLER_40_3141 ();
 sg13g2_decap_4 FILLER_40_3147 ();
 sg13g2_fill_1 FILLER_40_3209 ();
 sg13g2_decap_8 FILLER_40_3228 ();
 sg13g2_decap_4 FILLER_40_3235 ();
 sg13g2_decap_4 FILLER_40_3326 ();
 sg13g2_fill_2 FILLER_40_3330 ();
 sg13g2_decap_8 FILLER_40_3340 ();
 sg13g2_decap_8 FILLER_40_3347 ();
 sg13g2_decap_8 FILLER_40_3354 ();
 sg13g2_decap_8 FILLER_40_3361 ();
 sg13g2_decap_8 FILLER_40_3368 ();
 sg13g2_decap_8 FILLER_40_3375 ();
 sg13g2_decap_8 FILLER_40_3382 ();
 sg13g2_decap_8 FILLER_40_3389 ();
 sg13g2_decap_8 FILLER_40_3396 ();
 sg13g2_decap_8 FILLER_40_3403 ();
 sg13g2_decap_8 FILLER_40_3410 ();
 sg13g2_decap_8 FILLER_40_3417 ();
 sg13g2_decap_8 FILLER_40_3424 ();
 sg13g2_decap_8 FILLER_40_3431 ();
 sg13g2_decap_8 FILLER_40_3438 ();
 sg13g2_decap_8 FILLER_40_3445 ();
 sg13g2_decap_8 FILLER_40_3452 ();
 sg13g2_decap_8 FILLER_40_3459 ();
 sg13g2_decap_8 FILLER_40_3466 ();
 sg13g2_decap_8 FILLER_40_3473 ();
 sg13g2_decap_8 FILLER_40_3480 ();
 sg13g2_decap_8 FILLER_40_3487 ();
 sg13g2_decap_8 FILLER_40_3494 ();
 sg13g2_decap_8 FILLER_40_3501 ();
 sg13g2_decap_8 FILLER_40_3508 ();
 sg13g2_decap_8 FILLER_40_3515 ();
 sg13g2_decap_8 FILLER_40_3522 ();
 sg13g2_decap_8 FILLER_40_3529 ();
 sg13g2_decap_8 FILLER_40_3536 ();
 sg13g2_decap_8 FILLER_40_3543 ();
 sg13g2_decap_8 FILLER_40_3550 ();
 sg13g2_decap_8 FILLER_40_3557 ();
 sg13g2_decap_8 FILLER_40_3564 ();
 sg13g2_decap_8 FILLER_40_3571 ();
 sg13g2_fill_2 FILLER_40_3578 ();
 sg13g2_fill_1 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_65 ();
 sg13g2_fill_1 FILLER_41_77 ();
 sg13g2_decap_4 FILLER_41_129 ();
 sg13g2_decap_8 FILLER_41_137 ();
 sg13g2_fill_2 FILLER_41_144 ();
 sg13g2_fill_2 FILLER_41_165 ();
 sg13g2_decap_8 FILLER_41_170 ();
 sg13g2_decap_8 FILLER_41_181 ();
 sg13g2_fill_1 FILLER_41_188 ();
 sg13g2_decap_4 FILLER_41_199 ();
 sg13g2_fill_1 FILLER_41_203 ();
 sg13g2_fill_2 FILLER_41_225 ();
 sg13g2_decap_4 FILLER_41_278 ();
 sg13g2_fill_1 FILLER_41_282 ();
 sg13g2_decap_4 FILLER_41_289 ();
 sg13g2_fill_1 FILLER_41_293 ();
 sg13g2_decap_4 FILLER_41_304 ();
 sg13g2_decap_4 FILLER_41_313 ();
 sg13g2_decap_8 FILLER_41_323 ();
 sg13g2_fill_2 FILLER_41_330 ();
 sg13g2_fill_1 FILLER_41_332 ();
 sg13g2_decap_8 FILLER_41_337 ();
 sg13g2_fill_1 FILLER_41_357 ();
 sg13g2_decap_4 FILLER_41_394 ();
 sg13g2_fill_1 FILLER_41_422 ();
 sg13g2_fill_2 FILLER_41_462 ();
 sg13g2_fill_1 FILLER_41_464 ();
 sg13g2_fill_2 FILLER_41_486 ();
 sg13g2_decap_8 FILLER_41_554 ();
 sg13g2_fill_2 FILLER_41_561 ();
 sg13g2_decap_8 FILLER_41_568 ();
 sg13g2_fill_1 FILLER_41_575 ();
 sg13g2_fill_2 FILLER_41_589 ();
 sg13g2_fill_1 FILLER_41_617 ();
 sg13g2_decap_4 FILLER_41_650 ();
 sg13g2_fill_1 FILLER_41_654 ();
 sg13g2_decap_8 FILLER_41_660 ();
 sg13g2_decap_4 FILLER_41_667 ();
 sg13g2_fill_1 FILLER_41_671 ();
 sg13g2_fill_2 FILLER_41_703 ();
 sg13g2_decap_8 FILLER_41_772 ();
 sg13g2_fill_1 FILLER_41_779 ();
 sg13g2_fill_1 FILLER_41_806 ();
 sg13g2_fill_1 FILLER_41_822 ();
 sg13g2_fill_2 FILLER_41_840 ();
 sg13g2_decap_4 FILLER_41_900 ();
 sg13g2_fill_2 FILLER_41_912 ();
 sg13g2_fill_1 FILLER_41_914 ();
 sg13g2_decap_8 FILLER_41_966 ();
 sg13g2_fill_1 FILLER_41_1002 ();
 sg13g2_decap_4 FILLER_41_1007 ();
 sg13g2_fill_2 FILLER_41_1011 ();
 sg13g2_fill_1 FILLER_41_1039 ();
 sg13g2_fill_2 FILLER_41_1066 ();
 sg13g2_fill_2 FILLER_41_1078 ();
 sg13g2_fill_1 FILLER_41_1080 ();
 sg13g2_fill_1 FILLER_41_1107 ();
 sg13g2_fill_2 FILLER_41_1165 ();
 sg13g2_fill_1 FILLER_41_1167 ();
 sg13g2_decap_4 FILLER_41_1184 ();
 sg13g2_fill_1 FILLER_41_1197 ();
 sg13g2_fill_1 FILLER_41_1212 ();
 sg13g2_fill_2 FILLER_41_1222 ();
 sg13g2_fill_2 FILLER_41_1234 ();
 sg13g2_fill_1 FILLER_41_1236 ();
 sg13g2_decap_4 FILLER_41_1277 ();
 sg13g2_fill_1 FILLER_41_1281 ();
 sg13g2_decap_8 FILLER_41_1313 ();
 sg13g2_fill_1 FILLER_41_1320 ();
 sg13g2_fill_1 FILLER_41_1326 ();
 sg13g2_decap_8 FILLER_41_1345 ();
 sg13g2_decap_4 FILLER_41_1352 ();
 sg13g2_fill_1 FILLER_41_1356 ();
 sg13g2_fill_1 FILLER_41_1372 ();
 sg13g2_decap_4 FILLER_41_1377 ();
 sg13g2_fill_2 FILLER_41_1381 ();
 sg13g2_fill_2 FILLER_41_1394 ();
 sg13g2_fill_1 FILLER_41_1396 ();
 sg13g2_fill_1 FILLER_41_1407 ();
 sg13g2_decap_4 FILLER_41_1418 ();
 sg13g2_fill_2 FILLER_41_1422 ();
 sg13g2_fill_1 FILLER_41_1434 ();
 sg13g2_fill_2 FILLER_41_1440 ();
 sg13g2_fill_1 FILLER_41_1442 ();
 sg13g2_decap_8 FILLER_41_1451 ();
 sg13g2_fill_1 FILLER_41_1458 ();
 sg13g2_decap_8 FILLER_41_1468 ();
 sg13g2_decap_8 FILLER_41_1475 ();
 sg13g2_fill_2 FILLER_41_1482 ();
 sg13g2_fill_1 FILLER_41_1484 ();
 sg13g2_decap_8 FILLER_41_1519 ();
 sg13g2_fill_1 FILLER_41_1526 ();
 sg13g2_decap_8 FILLER_41_1540 ();
 sg13g2_decap_8 FILLER_41_1547 ();
 sg13g2_fill_2 FILLER_41_1554 ();
 sg13g2_fill_2 FILLER_41_1559 ();
 sg13g2_decap_8 FILLER_41_1565 ();
 sg13g2_decap_4 FILLER_41_1572 ();
 sg13g2_fill_2 FILLER_41_1576 ();
 sg13g2_decap_4 FILLER_41_1596 ();
 sg13g2_decap_8 FILLER_41_1612 ();
 sg13g2_decap_8 FILLER_41_1619 ();
 sg13g2_decap_4 FILLER_41_1626 ();
 sg13g2_fill_2 FILLER_41_1663 ();
 sg13g2_fill_2 FILLER_41_1670 ();
 sg13g2_fill_1 FILLER_41_1672 ();
 sg13g2_decap_8 FILLER_41_1687 ();
 sg13g2_fill_1 FILLER_41_1694 ();
 sg13g2_fill_2 FILLER_41_1706 ();
 sg13g2_fill_2 FILLER_41_1725 ();
 sg13g2_fill_1 FILLER_41_1727 ();
 sg13g2_fill_2 FILLER_41_1752 ();
 sg13g2_fill_1 FILLER_41_1754 ();
 sg13g2_fill_2 FILLER_41_1760 ();
 sg13g2_fill_1 FILLER_41_1762 ();
 sg13g2_fill_1 FILLER_41_1767 ();
 sg13g2_decap_4 FILLER_41_1783 ();
 sg13g2_fill_2 FILLER_41_1787 ();
 sg13g2_fill_2 FILLER_41_1805 ();
 sg13g2_fill_2 FILLER_41_1825 ();
 sg13g2_fill_2 FILLER_41_1832 ();
 sg13g2_decap_8 FILLER_41_1847 ();
 sg13g2_decap_4 FILLER_41_1854 ();
 sg13g2_fill_1 FILLER_41_1858 ();
 sg13g2_fill_2 FILLER_41_1865 ();
 sg13g2_fill_2 FILLER_41_1872 ();
 sg13g2_decap_4 FILLER_41_1878 ();
 sg13g2_decap_4 FILLER_41_1904 ();
 sg13g2_decap_4 FILLER_41_1917 ();
 sg13g2_decap_4 FILLER_41_1959 ();
 sg13g2_fill_1 FILLER_41_1963 ();
 sg13g2_fill_2 FILLER_41_1974 ();
 sg13g2_decap_8 FILLER_41_1984 ();
 sg13g2_decap_8 FILLER_41_2004 ();
 sg13g2_decap_4 FILLER_41_2011 ();
 sg13g2_fill_2 FILLER_41_2015 ();
 sg13g2_decap_8 FILLER_41_2033 ();
 sg13g2_decap_4 FILLER_41_2040 ();
 sg13g2_fill_1 FILLER_41_2044 ();
 sg13g2_decap_8 FILLER_41_2099 ();
 sg13g2_decap_4 FILLER_41_2124 ();
 sg13g2_fill_2 FILLER_41_2142 ();
 sg13g2_fill_1 FILLER_41_2144 ();
 sg13g2_decap_4 FILLER_41_2150 ();
 sg13g2_fill_1 FILLER_41_2154 ();
 sg13g2_decap_8 FILLER_41_2176 ();
 sg13g2_decap_8 FILLER_41_2183 ();
 sg13g2_fill_2 FILLER_41_2190 ();
 sg13g2_fill_1 FILLER_41_2192 ();
 sg13g2_fill_2 FILLER_41_2197 ();
 sg13g2_fill_1 FILLER_41_2199 ();
 sg13g2_decap_8 FILLER_41_2205 ();
 sg13g2_fill_2 FILLER_41_2212 ();
 sg13g2_fill_2 FILLER_41_2235 ();
 sg13g2_fill_1 FILLER_41_2237 ();
 sg13g2_fill_1 FILLER_41_2243 ();
 sg13g2_fill_2 FILLER_41_2254 ();
 sg13g2_decap_8 FILLER_41_2282 ();
 sg13g2_decap_8 FILLER_41_2289 ();
 sg13g2_fill_2 FILLER_41_2296 ();
 sg13g2_fill_1 FILLER_41_2298 ();
 sg13g2_decap_8 FILLER_41_2311 ();
 sg13g2_fill_2 FILLER_41_2318 ();
 sg13g2_fill_1 FILLER_41_2325 ();
 sg13g2_decap_8 FILLER_41_2330 ();
 sg13g2_decap_8 FILLER_41_2337 ();
 sg13g2_fill_1 FILLER_41_2344 ();
 sg13g2_decap_4 FILLER_41_2355 ();
 sg13g2_fill_2 FILLER_41_2381 ();
 sg13g2_fill_1 FILLER_41_2383 ();
 sg13g2_decap_8 FILLER_41_2410 ();
 sg13g2_decap_4 FILLER_41_2427 ();
 sg13g2_fill_2 FILLER_41_2431 ();
 sg13g2_fill_1 FILLER_41_2443 ();
 sg13g2_fill_1 FILLER_41_2448 ();
 sg13g2_fill_1 FILLER_41_2482 ();
 sg13g2_fill_2 FILLER_41_2503 ();
 sg13g2_fill_2 FILLER_41_2510 ();
 sg13g2_fill_2 FILLER_41_2517 ();
 sg13g2_fill_1 FILLER_41_2519 ();
 sg13g2_decap_8 FILLER_41_2524 ();
 sg13g2_decap_8 FILLER_41_2531 ();
 sg13g2_decap_8 FILLER_41_2538 ();
 sg13g2_fill_2 FILLER_41_2549 ();
 sg13g2_fill_1 FILLER_41_2551 ();
 sg13g2_decap_8 FILLER_41_2557 ();
 sg13g2_decap_8 FILLER_41_2564 ();
 sg13g2_fill_2 FILLER_41_2571 ();
 sg13g2_decap_8 FILLER_41_2577 ();
 sg13g2_fill_2 FILLER_41_2584 ();
 sg13g2_fill_1 FILLER_41_2586 ();
 sg13g2_decap_4 FILLER_41_2594 ();
 sg13g2_fill_2 FILLER_41_2598 ();
 sg13g2_fill_1 FILLER_41_2605 ();
 sg13g2_fill_2 FILLER_41_2668 ();
 sg13g2_fill_1 FILLER_41_2670 ();
 sg13g2_decap_8 FILLER_41_2705 ();
 sg13g2_decap_8 FILLER_41_2712 ();
 sg13g2_fill_2 FILLER_41_2762 ();
 sg13g2_fill_1 FILLER_41_2764 ();
 sg13g2_fill_1 FILLER_41_2769 ();
 sg13g2_fill_1 FILLER_41_2775 ();
 sg13g2_fill_2 FILLER_41_2780 ();
 sg13g2_fill_1 FILLER_41_2782 ();
 sg13g2_decap_8 FILLER_41_2792 ();
 sg13g2_fill_1 FILLER_41_2799 ();
 sg13g2_fill_2 FILLER_41_2805 ();
 sg13g2_fill_1 FILLER_41_2807 ();
 sg13g2_decap_4 FILLER_41_2812 ();
 sg13g2_fill_1 FILLER_41_2816 ();
 sg13g2_fill_2 FILLER_41_2848 ();
 sg13g2_decap_4 FILLER_41_2876 ();
 sg13g2_fill_2 FILLER_41_2919 ();
 sg13g2_decap_8 FILLER_41_2930 ();
 sg13g2_decap_8 FILLER_41_2937 ();
 sg13g2_decap_8 FILLER_41_2984 ();
 sg13g2_decap_4 FILLER_41_2991 ();
 sg13g2_fill_2 FILLER_41_2995 ();
 sg13g2_decap_4 FILLER_41_3010 ();
 sg13g2_decap_4 FILLER_41_3028 ();
 sg13g2_fill_1 FILLER_41_3032 ();
 sg13g2_decap_4 FILLER_41_3045 ();
 sg13g2_fill_2 FILLER_41_3058 ();
 sg13g2_fill_1 FILLER_41_3060 ();
 sg13g2_decap_8 FILLER_41_3083 ();
 sg13g2_fill_2 FILLER_41_3090 ();
 sg13g2_fill_1 FILLER_41_3092 ();
 sg13g2_decap_4 FILLER_41_3097 ();
 sg13g2_fill_2 FILLER_41_3101 ();
 sg13g2_fill_2 FILLER_41_3108 ();
 sg13g2_decap_8 FILLER_41_3114 ();
 sg13g2_decap_8 FILLER_41_3121 ();
 sg13g2_decap_4 FILLER_41_3128 ();
 sg13g2_decap_8 FILLER_41_3163 ();
 sg13g2_decap_4 FILLER_41_3170 ();
 sg13g2_fill_2 FILLER_41_3174 ();
 sg13g2_decap_8 FILLER_41_3180 ();
 sg13g2_decap_8 FILLER_41_3187 ();
 sg13g2_fill_1 FILLER_41_3220 ();
 sg13g2_decap_8 FILLER_41_3252 ();
 sg13g2_decap_8 FILLER_41_3259 ();
 sg13g2_decap_8 FILLER_41_3266 ();
 sg13g2_fill_2 FILLER_41_3273 ();
 sg13g2_decap_8 FILLER_41_3279 ();
 sg13g2_decap_4 FILLER_41_3286 ();
 sg13g2_fill_2 FILLER_41_3290 ();
 sg13g2_decap_4 FILLER_41_3296 ();
 sg13g2_fill_1 FILLER_41_3300 ();
 sg13g2_fill_2 FILLER_41_3319 ();
 sg13g2_decap_8 FILLER_41_3347 ();
 sg13g2_decap_8 FILLER_41_3354 ();
 sg13g2_decap_8 FILLER_41_3361 ();
 sg13g2_decap_8 FILLER_41_3368 ();
 sg13g2_decap_8 FILLER_41_3375 ();
 sg13g2_decap_8 FILLER_41_3382 ();
 sg13g2_decap_8 FILLER_41_3389 ();
 sg13g2_decap_8 FILLER_41_3396 ();
 sg13g2_decap_8 FILLER_41_3403 ();
 sg13g2_decap_8 FILLER_41_3410 ();
 sg13g2_decap_8 FILLER_41_3417 ();
 sg13g2_decap_8 FILLER_41_3424 ();
 sg13g2_decap_8 FILLER_41_3431 ();
 sg13g2_decap_8 FILLER_41_3438 ();
 sg13g2_decap_8 FILLER_41_3445 ();
 sg13g2_decap_8 FILLER_41_3452 ();
 sg13g2_decap_8 FILLER_41_3459 ();
 sg13g2_decap_8 FILLER_41_3466 ();
 sg13g2_decap_8 FILLER_41_3473 ();
 sg13g2_decap_8 FILLER_41_3480 ();
 sg13g2_decap_8 FILLER_41_3487 ();
 sg13g2_decap_8 FILLER_41_3494 ();
 sg13g2_decap_8 FILLER_41_3501 ();
 sg13g2_decap_8 FILLER_41_3508 ();
 sg13g2_decap_8 FILLER_41_3515 ();
 sg13g2_decap_8 FILLER_41_3522 ();
 sg13g2_decap_8 FILLER_41_3529 ();
 sg13g2_decap_8 FILLER_41_3536 ();
 sg13g2_decap_8 FILLER_41_3543 ();
 sg13g2_decap_8 FILLER_41_3550 ();
 sg13g2_decap_8 FILLER_41_3557 ();
 sg13g2_decap_8 FILLER_41_3564 ();
 sg13g2_decap_8 FILLER_41_3571 ();
 sg13g2_fill_2 FILLER_41_3578 ();
 sg13g2_decap_4 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_4 ();
 sg13g2_fill_1 FILLER_42_40 ();
 sg13g2_fill_1 FILLER_42_50 ();
 sg13g2_fill_2 FILLER_42_76 ();
 sg13g2_fill_1 FILLER_42_88 ();
 sg13g2_fill_2 FILLER_42_93 ();
 sg13g2_fill_1 FILLER_42_108 ();
 sg13g2_fill_2 FILLER_42_153 ();
 sg13g2_decap_4 FILLER_42_181 ();
 sg13g2_fill_1 FILLER_42_185 ();
 sg13g2_fill_2 FILLER_42_191 ();
 sg13g2_decap_8 FILLER_42_198 ();
 sg13g2_decap_8 FILLER_42_205 ();
 sg13g2_decap_4 FILLER_42_212 ();
 sg13g2_fill_1 FILLER_42_216 ();
 sg13g2_fill_1 FILLER_42_225 ();
 sg13g2_decap_8 FILLER_42_230 ();
 sg13g2_decap_8 FILLER_42_237 ();
 sg13g2_decap_8 FILLER_42_244 ();
 sg13g2_decap_8 FILLER_42_251 ();
 sg13g2_decap_4 FILLER_42_258 ();
 sg13g2_fill_2 FILLER_42_280 ();
 sg13g2_fill_1 FILLER_42_304 ();
 sg13g2_decap_8 FILLER_42_341 ();
 sg13g2_decap_8 FILLER_42_348 ();
 sg13g2_decap_4 FILLER_42_355 ();
 sg13g2_fill_1 FILLER_42_375 ();
 sg13g2_fill_2 FILLER_42_389 ();
 sg13g2_fill_1 FILLER_42_449 ();
 sg13g2_fill_2 FILLER_42_460 ();
 sg13g2_fill_1 FILLER_42_462 ();
 sg13g2_fill_2 FILLER_42_468 ();
 sg13g2_decap_8 FILLER_42_484 ();
 sg13g2_fill_1 FILLER_42_491 ();
 sg13g2_fill_2 FILLER_42_501 ();
 sg13g2_decap_4 FILLER_42_516 ();
 sg13g2_fill_2 FILLER_42_530 ();
 sg13g2_decap_8 FILLER_42_535 ();
 sg13g2_fill_2 FILLER_42_542 ();
 sg13g2_fill_2 FILLER_42_557 ();
 sg13g2_fill_1 FILLER_42_563 ();
 sg13g2_decap_4 FILLER_42_573 ();
 sg13g2_fill_1 FILLER_42_577 ();
 sg13g2_fill_2 FILLER_42_604 ();
 sg13g2_decap_8 FILLER_42_611 ();
 sg13g2_decap_8 FILLER_42_618 ();
 sg13g2_decap_8 FILLER_42_625 ();
 sg13g2_decap_8 FILLER_42_637 ();
 sg13g2_decap_8 FILLER_42_644 ();
 sg13g2_decap_4 FILLER_42_651 ();
 sg13g2_fill_2 FILLER_42_678 ();
 sg13g2_decap_4 FILLER_42_686 ();
 sg13g2_decap_4 FILLER_42_695 ();
 sg13g2_fill_1 FILLER_42_699 ();
 sg13g2_fill_2 FILLER_42_726 ();
 sg13g2_decap_4 FILLER_42_760 ();
 sg13g2_fill_2 FILLER_42_764 ();
 sg13g2_fill_2 FILLER_42_796 ();
 sg13g2_fill_1 FILLER_42_798 ();
 sg13g2_decap_8 FILLER_42_873 ();
 sg13g2_fill_1 FILLER_42_880 ();
 sg13g2_fill_1 FILLER_42_896 ();
 sg13g2_decap_8 FILLER_42_905 ();
 sg13g2_fill_2 FILLER_42_916 ();
 sg13g2_decap_4 FILLER_42_922 ();
 sg13g2_decap_4 FILLER_42_930 ();
 sg13g2_fill_1 FILLER_42_940 ();
 sg13g2_fill_1 FILLER_42_959 ();
 sg13g2_decap_4 FILLER_42_1018 ();
 sg13g2_fill_2 FILLER_42_1022 ();
 sg13g2_fill_1 FILLER_42_1028 ();
 sg13g2_decap_8 FILLER_42_1033 ();
 sg13g2_fill_2 FILLER_42_1040 ();
 sg13g2_fill_1 FILLER_42_1042 ();
 sg13g2_decap_8 FILLER_42_1048 ();
 sg13g2_decap_4 FILLER_42_1055 ();
 sg13g2_fill_2 FILLER_42_1068 ();
 sg13g2_fill_1 FILLER_42_1070 ();
 sg13g2_fill_1 FILLER_42_1080 ();
 sg13g2_fill_1 FILLER_42_1091 ();
 sg13g2_fill_2 FILLER_42_1096 ();
 sg13g2_fill_1 FILLER_42_1098 ();
 sg13g2_decap_8 FILLER_42_1107 ();
 sg13g2_fill_1 FILLER_42_1114 ();
 sg13g2_fill_2 FILLER_42_1137 ();
 sg13g2_decap_4 FILLER_42_1179 ();
 sg13g2_fill_1 FILLER_42_1183 ();
 sg13g2_fill_1 FILLER_42_1220 ();
 sg13g2_fill_1 FILLER_42_1232 ();
 sg13g2_fill_2 FILLER_42_1245 ();
 sg13g2_fill_1 FILLER_42_1247 ();
 sg13g2_fill_2 FILLER_42_1267 ();
 sg13g2_fill_1 FILLER_42_1278 ();
 sg13g2_decap_8 FILLER_42_1303 ();
 sg13g2_decap_8 FILLER_42_1310 ();
 sg13g2_decap_8 FILLER_42_1321 ();
 sg13g2_fill_2 FILLER_42_1328 ();
 sg13g2_fill_1 FILLER_42_1343 ();
 sg13g2_decap_4 FILLER_42_1377 ();
 sg13g2_decap_4 FILLER_42_1386 ();
 sg13g2_fill_1 FILLER_42_1390 ();
 sg13g2_fill_2 FILLER_42_1395 ();
 sg13g2_fill_1 FILLER_42_1397 ();
 sg13g2_fill_2 FILLER_42_1402 ();
 sg13g2_fill_2 FILLER_42_1408 ();
 sg13g2_fill_1 FILLER_42_1410 ();
 sg13g2_decap_8 FILLER_42_1421 ();
 sg13g2_decap_4 FILLER_42_1428 ();
 sg13g2_decap_8 FILLER_42_1455 ();
 sg13g2_decap_4 FILLER_42_1462 ();
 sg13g2_fill_2 FILLER_42_1466 ();
 sg13g2_fill_1 FILLER_42_1480 ();
 sg13g2_decap_8 FILLER_42_1491 ();
 sg13g2_decap_4 FILLER_42_1498 ();
 sg13g2_fill_1 FILLER_42_1502 ();
 sg13g2_fill_2 FILLER_42_1515 ();
 sg13g2_fill_2 FILLER_42_1526 ();
 sg13g2_fill_1 FILLER_42_1528 ();
 sg13g2_fill_2 FILLER_42_1533 ();
 sg13g2_fill_1 FILLER_42_1543 ();
 sg13g2_decap_4 FILLER_42_1576 ();
 sg13g2_fill_1 FILLER_42_1580 ();
 sg13g2_decap_8 FILLER_42_1586 ();
 sg13g2_decap_8 FILLER_42_1593 ();
 sg13g2_fill_1 FILLER_42_1600 ();
 sg13g2_fill_1 FILLER_42_1610 ();
 sg13g2_fill_1 FILLER_42_1616 ();
 sg13g2_decap_4 FILLER_42_1621 ();
 sg13g2_fill_2 FILLER_42_1625 ();
 sg13g2_decap_8 FILLER_42_1632 ();
 sg13g2_fill_2 FILLER_42_1663 ();
 sg13g2_fill_1 FILLER_42_1665 ();
 sg13g2_fill_1 FILLER_42_1677 ();
 sg13g2_fill_2 FILLER_42_1694 ();
 sg13g2_fill_1 FILLER_42_1696 ();
 sg13g2_fill_1 FILLER_42_1700 ();
 sg13g2_decap_4 FILLER_42_1716 ();
 sg13g2_fill_1 FILLER_42_1720 ();
 sg13g2_decap_4 FILLER_42_1739 ();
 sg13g2_fill_2 FILLER_42_1743 ();
 sg13g2_fill_1 FILLER_42_1771 ();
 sg13g2_fill_1 FILLER_42_1784 ();
 sg13g2_fill_2 FILLER_42_1803 ();
 sg13g2_fill_1 FILLER_42_1819 ();
 sg13g2_decap_8 FILLER_42_1895 ();
 sg13g2_fill_2 FILLER_42_1902 ();
 sg13g2_fill_1 FILLER_42_1904 ();
 sg13g2_fill_2 FILLER_42_1908 ();
 sg13g2_fill_1 FILLER_42_1910 ();
 sg13g2_decap_8 FILLER_42_1921 ();
 sg13g2_decap_8 FILLER_42_1928 ();
 sg13g2_decap_8 FILLER_42_1940 ();
 sg13g2_fill_1 FILLER_42_1947 ();
 sg13g2_decap_8 FILLER_42_1953 ();
 sg13g2_decap_8 FILLER_42_1960 ();
 sg13g2_decap_4 FILLER_42_1979 ();
 sg13g2_fill_2 FILLER_42_1983 ();
 sg13g2_decap_4 FILLER_42_1990 ();
 sg13g2_decap_8 FILLER_42_1999 ();
 sg13g2_decap_4 FILLER_42_2006 ();
 sg13g2_fill_1 FILLER_42_2010 ();
 sg13g2_decap_8 FILLER_42_2034 ();
 sg13g2_decap_4 FILLER_42_2041 ();
 sg13g2_fill_2 FILLER_42_2045 ();
 sg13g2_decap_8 FILLER_42_2053 ();
 sg13g2_decap_8 FILLER_42_2060 ();
 sg13g2_decap_8 FILLER_42_2067 ();
 sg13g2_fill_2 FILLER_42_2074 ();
 sg13g2_decap_8 FILLER_42_2089 ();
 sg13g2_decap_8 FILLER_42_2096 ();
 sg13g2_decap_8 FILLER_42_2103 ();
 sg13g2_fill_1 FILLER_42_2110 ();
 sg13g2_decap_8 FILLER_42_2124 ();
 sg13g2_fill_1 FILLER_42_2131 ();
 sg13g2_decap_4 FILLER_42_2145 ();
 sg13g2_fill_1 FILLER_42_2155 ();
 sg13g2_fill_2 FILLER_42_2161 ();
 sg13g2_decap_4 FILLER_42_2171 ();
 sg13g2_fill_1 FILLER_42_2175 ();
 sg13g2_fill_2 FILLER_42_2189 ();
 sg13g2_fill_1 FILLER_42_2191 ();
 sg13g2_decap_8 FILLER_42_2197 ();
 sg13g2_fill_1 FILLER_42_2204 ();
 sg13g2_fill_2 FILLER_42_2209 ();
 sg13g2_decap_8 FILLER_42_2216 ();
 sg13g2_decap_4 FILLER_42_2227 ();
 sg13g2_fill_2 FILLER_42_2256 ();
 sg13g2_fill_1 FILLER_42_2258 ();
 sg13g2_decap_4 FILLER_42_2263 ();
 sg13g2_fill_2 FILLER_42_2267 ();
 sg13g2_fill_2 FILLER_42_2273 ();
 sg13g2_fill_1 FILLER_42_2275 ();
 sg13g2_decap_8 FILLER_42_2281 ();
 sg13g2_fill_2 FILLER_42_2304 ();
 sg13g2_fill_1 FILLER_42_2311 ();
 sg13g2_decap_4 FILLER_42_2339 ();
 sg13g2_fill_1 FILLER_42_2343 ();
 sg13g2_fill_2 FILLER_42_2369 ();
 sg13g2_fill_1 FILLER_42_2371 ();
 sg13g2_decap_4 FILLER_42_2377 ();
 sg13g2_fill_2 FILLER_42_2381 ();
 sg13g2_fill_2 FILLER_42_2387 ();
 sg13g2_fill_2 FILLER_42_2407 ();
 sg13g2_fill_2 FILLER_42_2435 ();
 sg13g2_fill_2 FILLER_42_2441 ();
 sg13g2_fill_2 FILLER_42_2456 ();
 sg13g2_fill_1 FILLER_42_2458 ();
 sg13g2_fill_2 FILLER_42_2467 ();
 sg13g2_fill_1 FILLER_42_2469 ();
 sg13g2_fill_2 FILLER_42_2483 ();
 sg13g2_decap_4 FILLER_42_2490 ();
 sg13g2_fill_1 FILLER_42_2494 ();
 sg13g2_decap_8 FILLER_42_2504 ();
 sg13g2_fill_1 FILLER_42_2511 ();
 sg13g2_decap_4 FILLER_42_2520 ();
 sg13g2_fill_1 FILLER_42_2524 ();
 sg13g2_fill_1 FILLER_42_2549 ();
 sg13g2_fill_2 FILLER_42_2583 ();
 sg13g2_fill_1 FILLER_42_2625 ();
 sg13g2_fill_2 FILLER_42_2651 ();
 sg13g2_fill_2 FILLER_42_2657 ();
 sg13g2_decap_8 FILLER_42_2663 ();
 sg13g2_decap_8 FILLER_42_2670 ();
 sg13g2_decap_8 FILLER_42_2677 ();
 sg13g2_fill_1 FILLER_42_2684 ();
 sg13g2_decap_8 FILLER_42_2689 ();
 sg13g2_decap_8 FILLER_42_2696 ();
 sg13g2_decap_8 FILLER_42_2703 ();
 sg13g2_decap_8 FILLER_42_2710 ();
 sg13g2_decap_8 FILLER_42_2717 ();
 sg13g2_decap_8 FILLER_42_2724 ();
 sg13g2_decap_8 FILLER_42_2731 ();
 sg13g2_decap_8 FILLER_42_2738 ();
 sg13g2_decap_8 FILLER_42_2745 ();
 sg13g2_decap_8 FILLER_42_2752 ();
 sg13g2_decap_4 FILLER_42_2759 ();
 sg13g2_fill_2 FILLER_42_2789 ();
 sg13g2_fill_1 FILLER_42_2791 ();
 sg13g2_decap_8 FILLER_42_2849 ();
 sg13g2_decap_4 FILLER_42_2856 ();
 sg13g2_fill_1 FILLER_42_2860 ();
 sg13g2_decap_4 FILLER_42_2874 ();
 sg13g2_fill_2 FILLER_42_2887 ();
 sg13g2_decap_4 FILLER_42_2898 ();
 sg13g2_fill_2 FILLER_42_2902 ();
 sg13g2_fill_2 FILLER_42_2966 ();
 sg13g2_decap_8 FILLER_42_2985 ();
 sg13g2_decap_8 FILLER_42_2992 ();
 sg13g2_decap_4 FILLER_42_3025 ();
 sg13g2_fill_1 FILLER_42_3029 ();
 sg13g2_fill_2 FILLER_42_3056 ();
 sg13g2_decap_8 FILLER_42_3084 ();
 sg13g2_decap_8 FILLER_42_3091 ();
 sg13g2_fill_1 FILLER_42_3098 ();
 sg13g2_fill_2 FILLER_42_3139 ();
 sg13g2_fill_1 FILLER_42_3158 ();
 sg13g2_fill_1 FILLER_42_3164 ();
 sg13g2_decap_4 FILLER_42_3169 ();
 sg13g2_fill_2 FILLER_42_3173 ();
 sg13g2_fill_2 FILLER_42_3198 ();
 sg13g2_fill_1 FILLER_42_3200 ();
 sg13g2_decap_8 FILLER_42_3214 ();
 sg13g2_decap_4 FILLER_42_3221 ();
 sg13g2_fill_2 FILLER_42_3225 ();
 sg13g2_decap_4 FILLER_42_3231 ();
 sg13g2_fill_1 FILLER_42_3235 ();
 sg13g2_decap_8 FILLER_42_3249 ();
 sg13g2_decap_8 FILLER_42_3256 ();
 sg13g2_decap_8 FILLER_42_3263 ();
 sg13g2_decap_8 FILLER_42_3270 ();
 sg13g2_decap_8 FILLER_42_3277 ();
 sg13g2_decap_8 FILLER_42_3284 ();
 sg13g2_decap_8 FILLER_42_3291 ();
 sg13g2_decap_8 FILLER_42_3298 ();
 sg13g2_decap_4 FILLER_42_3305 ();
 sg13g2_fill_1 FILLER_42_3309 ();
 sg13g2_decap_8 FILLER_42_3314 ();
 sg13g2_decap_8 FILLER_42_3321 ();
 sg13g2_fill_1 FILLER_42_3328 ();
 sg13g2_decap_8 FILLER_42_3338 ();
 sg13g2_decap_8 FILLER_42_3345 ();
 sg13g2_decap_8 FILLER_42_3352 ();
 sg13g2_decap_8 FILLER_42_3359 ();
 sg13g2_decap_8 FILLER_42_3366 ();
 sg13g2_decap_8 FILLER_42_3373 ();
 sg13g2_decap_8 FILLER_42_3380 ();
 sg13g2_decap_8 FILLER_42_3387 ();
 sg13g2_decap_8 FILLER_42_3394 ();
 sg13g2_decap_8 FILLER_42_3401 ();
 sg13g2_decap_8 FILLER_42_3408 ();
 sg13g2_decap_8 FILLER_42_3415 ();
 sg13g2_decap_8 FILLER_42_3422 ();
 sg13g2_decap_8 FILLER_42_3429 ();
 sg13g2_decap_8 FILLER_42_3436 ();
 sg13g2_decap_8 FILLER_42_3443 ();
 sg13g2_decap_8 FILLER_42_3450 ();
 sg13g2_decap_8 FILLER_42_3457 ();
 sg13g2_decap_8 FILLER_42_3464 ();
 sg13g2_decap_8 FILLER_42_3471 ();
 sg13g2_decap_8 FILLER_42_3478 ();
 sg13g2_decap_8 FILLER_42_3485 ();
 sg13g2_decap_8 FILLER_42_3492 ();
 sg13g2_decap_8 FILLER_42_3499 ();
 sg13g2_decap_8 FILLER_42_3506 ();
 sg13g2_decap_8 FILLER_42_3513 ();
 sg13g2_decap_8 FILLER_42_3520 ();
 sg13g2_decap_8 FILLER_42_3527 ();
 sg13g2_decap_8 FILLER_42_3534 ();
 sg13g2_decap_8 FILLER_42_3541 ();
 sg13g2_decap_8 FILLER_42_3548 ();
 sg13g2_decap_8 FILLER_42_3555 ();
 sg13g2_decap_8 FILLER_42_3562 ();
 sg13g2_decap_8 FILLER_42_3569 ();
 sg13g2_decap_4 FILLER_42_3576 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_4 FILLER_43_7 ();
 sg13g2_fill_1 FILLER_43_24 ();
 sg13g2_fill_2 FILLER_43_39 ();
 sg13g2_decap_8 FILLER_43_61 ();
 sg13g2_fill_1 FILLER_43_68 ();
 sg13g2_fill_2 FILLER_43_114 ();
 sg13g2_decap_8 FILLER_43_134 ();
 sg13g2_fill_2 FILLER_43_173 ();
 sg13g2_fill_1 FILLER_43_175 ();
 sg13g2_decap_4 FILLER_43_206 ();
 sg13g2_fill_2 FILLER_43_241 ();
 sg13g2_fill_2 FILLER_43_258 ();
 sg13g2_fill_1 FILLER_43_260 ();
 sg13g2_decap_8 FILLER_43_266 ();
 sg13g2_fill_2 FILLER_43_273 ();
 sg13g2_decap_8 FILLER_43_287 ();
 sg13g2_decap_8 FILLER_43_294 ();
 sg13g2_decap_4 FILLER_43_301 ();
 sg13g2_fill_1 FILLER_43_305 ();
 sg13g2_fill_1 FILLER_43_339 ();
 sg13g2_fill_2 FILLER_43_344 ();
 sg13g2_decap_4 FILLER_43_352 ();
 sg13g2_fill_2 FILLER_43_361 ();
 sg13g2_fill_1 FILLER_43_363 ();
 sg13g2_decap_8 FILLER_43_390 ();
 sg13g2_fill_2 FILLER_43_397 ();
 sg13g2_decap_8 FILLER_43_403 ();
 sg13g2_fill_2 FILLER_43_410 ();
 sg13g2_fill_2 FILLER_43_416 ();
 sg13g2_fill_1 FILLER_43_418 ();
 sg13g2_fill_1 FILLER_43_424 ();
 sg13g2_fill_1 FILLER_43_434 ();
 sg13g2_decap_8 FILLER_43_467 ();
 sg13g2_decap_8 FILLER_43_474 ();
 sg13g2_fill_2 FILLER_43_494 ();
 sg13g2_decap_8 FILLER_43_509 ();
 sg13g2_fill_2 FILLER_43_516 ();
 sg13g2_fill_1 FILLER_43_518 ();
 sg13g2_fill_2 FILLER_43_527 ();
 sg13g2_decap_8 FILLER_43_578 ();
 sg13g2_fill_2 FILLER_43_598 ();
 sg13g2_fill_2 FILLER_43_609 ();
 sg13g2_fill_1 FILLER_43_616 ();
 sg13g2_fill_1 FILLER_43_634 ();
 sg13g2_decap_4 FILLER_43_639 ();
 sg13g2_fill_1 FILLER_43_643 ();
 sg13g2_decap_8 FILLER_43_648 ();
 sg13g2_fill_2 FILLER_43_655 ();
 sg13g2_decap_8 FILLER_43_665 ();
 sg13g2_decap_4 FILLER_43_672 ();
 sg13g2_fill_2 FILLER_43_690 ();
 sg13g2_fill_2 FILLER_43_700 ();
 sg13g2_fill_1 FILLER_43_702 ();
 sg13g2_fill_1 FILLER_43_724 ();
 sg13g2_fill_1 FILLER_43_734 ();
 sg13g2_fill_1 FILLER_43_741 ();
 sg13g2_decap_4 FILLER_43_768 ();
 sg13g2_fill_1 FILLER_43_772 ();
 sg13g2_decap_4 FILLER_43_804 ();
 sg13g2_fill_2 FILLER_43_808 ();
 sg13g2_fill_1 FILLER_43_849 ();
 sg13g2_fill_2 FILLER_43_864 ();
 sg13g2_fill_1 FILLER_43_866 ();
 sg13g2_fill_1 FILLER_43_889 ();
 sg13g2_fill_2 FILLER_43_901 ();
 sg13g2_fill_1 FILLER_43_940 ();
 sg13g2_fill_1 FILLER_43_973 ();
 sg13g2_decap_8 FILLER_43_1006 ();
 sg13g2_fill_1 FILLER_43_1013 ();
 sg13g2_fill_2 FILLER_43_1097 ();
 sg13g2_fill_1 FILLER_43_1099 ();
 sg13g2_fill_2 FILLER_43_1140 ();
 sg13g2_fill_1 FILLER_43_1142 ();
 sg13g2_decap_8 FILLER_43_1160 ();
 sg13g2_fill_2 FILLER_43_1167 ();
 sg13g2_fill_1 FILLER_43_1169 ();
 sg13g2_decap_8 FILLER_43_1184 ();
 sg13g2_fill_2 FILLER_43_1191 ();
 sg13g2_fill_1 FILLER_43_1193 ();
 sg13g2_decap_4 FILLER_43_1198 ();
 sg13g2_fill_1 FILLER_43_1202 ();
 sg13g2_fill_2 FILLER_43_1208 ();
 sg13g2_decap_4 FILLER_43_1214 ();
 sg13g2_fill_2 FILLER_43_1218 ();
 sg13g2_fill_1 FILLER_43_1224 ();
 sg13g2_fill_1 FILLER_43_1246 ();
 sg13g2_fill_2 FILLER_43_1255 ();
 sg13g2_fill_1 FILLER_43_1257 ();
 sg13g2_fill_1 FILLER_43_1264 ();
 sg13g2_decap_8 FILLER_43_1291 ();
 sg13g2_decap_8 FILLER_43_1298 ();
 sg13g2_fill_1 FILLER_43_1305 ();
 sg13g2_decap_8 FILLER_43_1348 ();
 sg13g2_fill_1 FILLER_43_1355 ();
 sg13g2_fill_2 FILLER_43_1377 ();
 sg13g2_fill_1 FILLER_43_1379 ();
 sg13g2_fill_2 FILLER_43_1390 ();
 sg13g2_fill_1 FILLER_43_1392 ();
 sg13g2_fill_2 FILLER_43_1398 ();
 sg13g2_decap_4 FILLER_43_1421 ();
 sg13g2_fill_2 FILLER_43_1425 ();
 sg13g2_decap_8 FILLER_43_1446 ();
 sg13g2_fill_2 FILLER_43_1453 ();
 sg13g2_fill_1 FILLER_43_1455 ();
 sg13g2_fill_1 FILLER_43_1461 ();
 sg13g2_decap_8 FILLER_43_1475 ();
 sg13g2_decap_8 FILLER_43_1482 ();
 sg13g2_fill_2 FILLER_43_1515 ();
 sg13g2_fill_1 FILLER_43_1517 ();
 sg13g2_fill_2 FILLER_43_1573 ();
 sg13g2_fill_1 FILLER_43_1575 ();
 sg13g2_decap_4 FILLER_43_1602 ();
 sg13g2_fill_1 FILLER_43_1649 ();
 sg13g2_decap_8 FILLER_43_1666 ();
 sg13g2_decap_4 FILLER_43_1673 ();
 sg13g2_fill_1 FILLER_43_1677 ();
 sg13g2_decap_8 FILLER_43_1684 ();
 sg13g2_fill_2 FILLER_43_1691 ();
 sg13g2_fill_2 FILLER_43_1703 ();
 sg13g2_decap_8 FILLER_43_1736 ();
 sg13g2_decap_4 FILLER_43_1751 ();
 sg13g2_fill_1 FILLER_43_1755 ();
 sg13g2_fill_1 FILLER_43_1760 ();
 sg13g2_decap_8 FILLER_43_1788 ();
 sg13g2_decap_4 FILLER_43_1795 ();
 sg13g2_fill_2 FILLER_43_1816 ();
 sg13g2_fill_1 FILLER_43_1818 ();
 sg13g2_decap_4 FILLER_43_1827 ();
 sg13g2_fill_2 FILLER_43_1835 ();
 sg13g2_decap_8 FILLER_43_1842 ();
 sg13g2_decap_8 FILLER_43_1849 ();
 sg13g2_fill_2 FILLER_43_1856 ();
 sg13g2_decap_4 FILLER_43_1867 ();
 sg13g2_fill_2 FILLER_43_1871 ();
 sg13g2_fill_2 FILLER_43_1884 ();
 sg13g2_fill_1 FILLER_43_1886 ();
 sg13g2_decap_8 FILLER_43_1932 ();
 sg13g2_fill_1 FILLER_43_1939 ();
 sg13g2_fill_2 FILLER_43_1959 ();
 sg13g2_fill_1 FILLER_43_1961 ();
 sg13g2_decap_8 FILLER_43_1976 ();
 sg13g2_fill_2 FILLER_43_1983 ();
 sg13g2_fill_1 FILLER_43_1985 ();
 sg13g2_decap_8 FILLER_43_2009 ();
 sg13g2_decap_4 FILLER_43_2016 ();
 sg13g2_fill_1 FILLER_43_2039 ();
 sg13g2_fill_2 FILLER_43_2059 ();
 sg13g2_fill_2 FILLER_43_2067 ();
 sg13g2_fill_1 FILLER_43_2069 ();
 sg13g2_decap_4 FILLER_43_2078 ();
 sg13g2_fill_1 FILLER_43_2082 ();
 sg13g2_decap_8 FILLER_43_2091 ();
 sg13g2_decap_4 FILLER_43_2098 ();
 sg13g2_decap_4 FILLER_43_2121 ();
 sg13g2_fill_1 FILLER_43_2125 ();
 sg13g2_decap_8 FILLER_43_2134 ();
 sg13g2_decap_4 FILLER_43_2141 ();
 sg13g2_fill_1 FILLER_43_2145 ();
 sg13g2_fill_2 FILLER_43_2151 ();
 sg13g2_decap_8 FILLER_43_2166 ();
 sg13g2_fill_2 FILLER_43_2173 ();
 sg13g2_fill_2 FILLER_43_2203 ();
 sg13g2_decap_8 FILLER_43_2223 ();
 sg13g2_decap_8 FILLER_43_2230 ();
 sg13g2_decap_4 FILLER_43_2237 ();
 sg13g2_fill_2 FILLER_43_2250 ();
 sg13g2_fill_1 FILLER_43_2252 ();
 sg13g2_fill_2 FILLER_43_2271 ();
 sg13g2_decap_8 FILLER_43_2292 ();
 sg13g2_decap_4 FILLER_43_2308 ();
 sg13g2_fill_2 FILLER_43_2312 ();
 sg13g2_decap_4 FILLER_43_2319 ();
 sg13g2_fill_2 FILLER_43_2329 ();
 sg13g2_decap_8 FILLER_43_2344 ();
 sg13g2_decap_8 FILLER_43_2359 ();
 sg13g2_fill_2 FILLER_43_2375 ();
 sg13g2_fill_2 FILLER_43_2438 ();
 sg13g2_fill_1 FILLER_43_2440 ();
 sg13g2_decap_4 FILLER_43_2461 ();
 sg13g2_fill_1 FILLER_43_2465 ();
 sg13g2_fill_2 FILLER_43_2475 ();
 sg13g2_fill_1 FILLER_43_2477 ();
 sg13g2_fill_2 FILLER_43_2491 ();
 sg13g2_fill_1 FILLER_43_2493 ();
 sg13g2_fill_2 FILLER_43_2504 ();
 sg13g2_fill_1 FILLER_43_2514 ();
 sg13g2_decap_8 FILLER_43_2519 ();
 sg13g2_decap_4 FILLER_43_2526 ();
 sg13g2_fill_2 FILLER_43_2534 ();
 sg13g2_fill_1 FILLER_43_2536 ();
 sg13g2_decap_4 FILLER_43_2547 ();
 sg13g2_fill_1 FILLER_43_2551 ();
 sg13g2_decap_4 FILLER_43_2556 ();
 sg13g2_fill_1 FILLER_43_2560 ();
 sg13g2_fill_2 FILLER_43_2565 ();
 sg13g2_fill_1 FILLER_43_2567 ();
 sg13g2_fill_2 FILLER_43_2593 ();
 sg13g2_fill_1 FILLER_43_2595 ();
 sg13g2_fill_1 FILLER_43_2600 ();
 sg13g2_decap_4 FILLER_43_2634 ();
 sg13g2_fill_2 FILLER_43_2638 ();
 sg13g2_fill_2 FILLER_43_2647 ();
 sg13g2_decap_8 FILLER_43_2727 ();
 sg13g2_decap_8 FILLER_43_2734 ();
 sg13g2_decap_8 FILLER_43_2741 ();
 sg13g2_decap_8 FILLER_43_2748 ();
 sg13g2_decap_8 FILLER_43_2755 ();
 sg13g2_fill_2 FILLER_43_2762 ();
 sg13g2_fill_1 FILLER_43_2764 ();
 sg13g2_decap_8 FILLER_43_2795 ();
 sg13g2_decap_4 FILLER_43_2802 ();
 sg13g2_fill_2 FILLER_43_2806 ();
 sg13g2_fill_1 FILLER_43_2812 ();
 sg13g2_decap_8 FILLER_43_2843 ();
 sg13g2_decap_8 FILLER_43_2850 ();
 sg13g2_fill_1 FILLER_43_2857 ();
 sg13g2_decap_4 FILLER_43_2884 ();
 sg13g2_fill_1 FILLER_43_2888 ();
 sg13g2_decap_8 FILLER_43_2915 ();
 sg13g2_decap_8 FILLER_43_2922 ();
 sg13g2_decap_8 FILLER_43_2929 ();
 sg13g2_fill_2 FILLER_43_2936 ();
 sg13g2_decap_8 FILLER_43_2942 ();
 sg13g2_decap_8 FILLER_43_2949 ();
 sg13g2_decap_4 FILLER_43_2956 ();
 sg13g2_decap_8 FILLER_43_2986 ();
 sg13g2_decap_8 FILLER_43_2993 ();
 sg13g2_decap_8 FILLER_43_3000 ();
 sg13g2_fill_2 FILLER_43_3007 ();
 sg13g2_fill_1 FILLER_43_3009 ();
 sg13g2_decap_8 FILLER_43_3014 ();
 sg13g2_decap_8 FILLER_43_3021 ();
 sg13g2_decap_4 FILLER_43_3028 ();
 sg13g2_fill_1 FILLER_43_3032 ();
 sg13g2_fill_2 FILLER_43_3038 ();
 sg13g2_fill_1 FILLER_43_3040 ();
 sg13g2_decap_8 FILLER_43_3045 ();
 sg13g2_decap_8 FILLER_43_3052 ();
 sg13g2_decap_8 FILLER_43_3059 ();
 sg13g2_fill_2 FILLER_43_3066 ();
 sg13g2_fill_1 FILLER_43_3068 ();
 sg13g2_decap_8 FILLER_43_3074 ();
 sg13g2_decap_8 FILLER_43_3081 ();
 sg13g2_decap_8 FILLER_43_3088 ();
 sg13g2_decap_8 FILLER_43_3095 ();
 sg13g2_decap_8 FILLER_43_3102 ();
 sg13g2_fill_1 FILLER_43_3109 ();
 sg13g2_decap_8 FILLER_43_3114 ();
 sg13g2_fill_2 FILLER_43_3121 ();
 sg13g2_decap_8 FILLER_43_3149 ();
 sg13g2_fill_1 FILLER_43_3156 ();
 sg13g2_fill_2 FILLER_43_3183 ();
 sg13g2_decap_8 FILLER_43_3211 ();
 sg13g2_decap_8 FILLER_43_3218 ();
 sg13g2_decap_8 FILLER_43_3225 ();
 sg13g2_decap_8 FILLER_43_3232 ();
 sg13g2_decap_8 FILLER_43_3239 ();
 sg13g2_decap_8 FILLER_43_3246 ();
 sg13g2_decap_8 FILLER_43_3253 ();
 sg13g2_decap_8 FILLER_43_3260 ();
 sg13g2_decap_8 FILLER_43_3267 ();
 sg13g2_decap_8 FILLER_43_3274 ();
 sg13g2_decap_8 FILLER_43_3281 ();
 sg13g2_decap_8 FILLER_43_3288 ();
 sg13g2_decap_8 FILLER_43_3295 ();
 sg13g2_decap_8 FILLER_43_3302 ();
 sg13g2_decap_8 FILLER_43_3309 ();
 sg13g2_decap_8 FILLER_43_3316 ();
 sg13g2_decap_8 FILLER_43_3323 ();
 sg13g2_decap_8 FILLER_43_3330 ();
 sg13g2_decap_8 FILLER_43_3337 ();
 sg13g2_decap_8 FILLER_43_3344 ();
 sg13g2_decap_8 FILLER_43_3351 ();
 sg13g2_decap_8 FILLER_43_3358 ();
 sg13g2_decap_8 FILLER_43_3365 ();
 sg13g2_decap_8 FILLER_43_3372 ();
 sg13g2_decap_8 FILLER_43_3379 ();
 sg13g2_decap_8 FILLER_43_3386 ();
 sg13g2_decap_8 FILLER_43_3393 ();
 sg13g2_decap_8 FILLER_43_3400 ();
 sg13g2_decap_8 FILLER_43_3407 ();
 sg13g2_decap_8 FILLER_43_3414 ();
 sg13g2_decap_8 FILLER_43_3421 ();
 sg13g2_decap_8 FILLER_43_3428 ();
 sg13g2_decap_8 FILLER_43_3435 ();
 sg13g2_decap_8 FILLER_43_3442 ();
 sg13g2_decap_8 FILLER_43_3449 ();
 sg13g2_decap_8 FILLER_43_3456 ();
 sg13g2_decap_8 FILLER_43_3463 ();
 sg13g2_decap_8 FILLER_43_3470 ();
 sg13g2_decap_8 FILLER_43_3477 ();
 sg13g2_decap_8 FILLER_43_3484 ();
 sg13g2_decap_8 FILLER_43_3491 ();
 sg13g2_decap_8 FILLER_43_3498 ();
 sg13g2_decap_8 FILLER_43_3505 ();
 sg13g2_decap_8 FILLER_43_3512 ();
 sg13g2_decap_8 FILLER_43_3519 ();
 sg13g2_decap_8 FILLER_43_3526 ();
 sg13g2_decap_8 FILLER_43_3533 ();
 sg13g2_decap_8 FILLER_43_3540 ();
 sg13g2_decap_8 FILLER_43_3547 ();
 sg13g2_decap_8 FILLER_43_3554 ();
 sg13g2_decap_8 FILLER_43_3561 ();
 sg13g2_decap_8 FILLER_43_3568 ();
 sg13g2_decap_4 FILLER_43_3575 ();
 sg13g2_fill_1 FILLER_43_3579 ();
 sg13g2_fill_2 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_28 ();
 sg13g2_fill_1 FILLER_44_30 ();
 sg13g2_fill_2 FILLER_44_41 ();
 sg13g2_decap_8 FILLER_44_86 ();
 sg13g2_decap_4 FILLER_44_93 ();
 sg13g2_fill_2 FILLER_44_97 ();
 sg13g2_fill_1 FILLER_44_103 ();
 sg13g2_fill_2 FILLER_44_109 ();
 sg13g2_fill_1 FILLER_44_111 ();
 sg13g2_fill_1 FILLER_44_138 ();
 sg13g2_decap_8 FILLER_44_156 ();
 sg13g2_decap_8 FILLER_44_163 ();
 sg13g2_fill_1 FILLER_44_170 ();
 sg13g2_decap_8 FILLER_44_176 ();
 sg13g2_fill_1 FILLER_44_183 ();
 sg13g2_decap_4 FILLER_44_189 ();
 sg13g2_decap_8 FILLER_44_216 ();
 sg13g2_fill_2 FILLER_44_223 ();
 sg13g2_decap_4 FILLER_44_239 ();
 sg13g2_fill_1 FILLER_44_243 ();
 sg13g2_decap_8 FILLER_44_256 ();
 sg13g2_decap_4 FILLER_44_263 ();
 sg13g2_fill_1 FILLER_44_267 ();
 sg13g2_fill_2 FILLER_44_281 ();
 sg13g2_fill_1 FILLER_44_283 ();
 sg13g2_fill_2 FILLER_44_293 ();
 sg13g2_fill_1 FILLER_44_295 ();
 sg13g2_decap_8 FILLER_44_300 ();
 sg13g2_decap_4 FILLER_44_307 ();
 sg13g2_decap_8 FILLER_44_353 ();
 sg13g2_fill_2 FILLER_44_360 ();
 sg13g2_fill_1 FILLER_44_362 ();
 sg13g2_fill_2 FILLER_44_415 ();
 sg13g2_fill_1 FILLER_44_417 ();
 sg13g2_fill_1 FILLER_44_423 ();
 sg13g2_fill_1 FILLER_44_448 ();
 sg13g2_decap_8 FILLER_44_469 ();
 sg13g2_decap_4 FILLER_44_476 ();
 sg13g2_fill_1 FILLER_44_480 ();
 sg13g2_decap_4 FILLER_44_512 ();
 sg13g2_fill_1 FILLER_44_516 ();
 sg13g2_decap_4 FILLER_44_522 ();
 sg13g2_fill_1 FILLER_44_526 ();
 sg13g2_fill_2 FILLER_44_561 ();
 sg13g2_fill_1 FILLER_44_563 ();
 sg13g2_decap_4 FILLER_44_573 ();
 sg13g2_decap_8 FILLER_44_581 ();
 sg13g2_decap_8 FILLER_44_588 ();
 sg13g2_fill_2 FILLER_44_595 ();
 sg13g2_fill_1 FILLER_44_597 ();
 sg13g2_fill_1 FILLER_44_608 ();
 sg13g2_fill_2 FILLER_44_633 ();
 sg13g2_fill_1 FILLER_44_665 ();
 sg13g2_fill_1 FILLER_44_692 ();
 sg13g2_fill_1 FILLER_44_711 ();
 sg13g2_fill_2 FILLER_44_727 ();
 sg13g2_fill_1 FILLER_44_748 ();
 sg13g2_decap_8 FILLER_44_768 ();
 sg13g2_decap_4 FILLER_44_775 ();
 sg13g2_fill_1 FILLER_44_794 ();
 sg13g2_decap_8 FILLER_44_806 ();
 sg13g2_decap_8 FILLER_44_813 ();
 sg13g2_fill_1 FILLER_44_820 ();
 sg13g2_fill_2 FILLER_44_825 ();
 sg13g2_fill_2 FILLER_44_830 ();
 sg13g2_fill_1 FILLER_44_842 ();
 sg13g2_decap_8 FILLER_44_874 ();
 sg13g2_fill_1 FILLER_44_901 ();
 sg13g2_fill_2 FILLER_44_915 ();
 sg13g2_decap_4 FILLER_44_953 ();
 sg13g2_fill_1 FILLER_44_957 ();
 sg13g2_fill_2 FILLER_44_962 ();
 sg13g2_fill_1 FILLER_44_976 ();
 sg13g2_decap_4 FILLER_44_1029 ();
 sg13g2_decap_8 FILLER_44_1052 ();
 sg13g2_fill_2 FILLER_44_1059 ();
 sg13g2_fill_2 FILLER_44_1071 ();
 sg13g2_fill_2 FILLER_44_1108 ();
 sg13g2_decap_4 FILLER_44_1138 ();
 sg13g2_fill_2 FILLER_44_1154 ();
 sg13g2_fill_1 FILLER_44_1156 ();
 sg13g2_decap_4 FILLER_44_1188 ();
 sg13g2_fill_1 FILLER_44_1192 ();
 sg13g2_decap_8 FILLER_44_1211 ();
 sg13g2_fill_2 FILLER_44_1218 ();
 sg13g2_fill_1 FILLER_44_1246 ();
 sg13g2_fill_1 FILLER_44_1260 ();
 sg13g2_decap_8 FILLER_44_1265 ();
 sg13g2_fill_1 FILLER_44_1272 ();
 sg13g2_fill_2 FILLER_44_1286 ();
 sg13g2_decap_4 FILLER_44_1301 ();
 sg13g2_fill_1 FILLER_44_1305 ();
 sg13g2_decap_8 FILLER_44_1311 ();
 sg13g2_fill_1 FILLER_44_1318 ();
 sg13g2_decap_4 FILLER_44_1356 ();
 sg13g2_fill_2 FILLER_44_1360 ();
 sg13g2_fill_2 FILLER_44_1375 ();
 sg13g2_fill_2 FILLER_44_1388 ();
 sg13g2_fill_1 FILLER_44_1390 ();
 sg13g2_fill_2 FILLER_44_1399 ();
 sg13g2_fill_2 FILLER_44_1405 ();
 sg13g2_decap_4 FILLER_44_1427 ();
 sg13g2_fill_2 FILLER_44_1431 ();
 sg13g2_decap_8 FILLER_44_1438 ();
 sg13g2_fill_1 FILLER_44_1445 ();
 sg13g2_decap_4 FILLER_44_1454 ();
 sg13g2_fill_2 FILLER_44_1471 ();
 sg13g2_fill_1 FILLER_44_1473 ();
 sg13g2_decap_8 FILLER_44_1492 ();
 sg13g2_fill_1 FILLER_44_1499 ();
 sg13g2_decap_4 FILLER_44_1518 ();
 sg13g2_fill_2 FILLER_44_1522 ();
 sg13g2_decap_8 FILLER_44_1569 ();
 sg13g2_decap_8 FILLER_44_1579 ();
 sg13g2_fill_1 FILLER_44_1586 ();
 sg13g2_decap_8 FILLER_44_1615 ();
 sg13g2_decap_8 FILLER_44_1622 ();
 sg13g2_decap_8 FILLER_44_1629 ();
 sg13g2_decap_8 FILLER_44_1636 ();
 sg13g2_fill_2 FILLER_44_1654 ();
 sg13g2_decap_4 FILLER_44_1662 ();
 sg13g2_fill_2 FILLER_44_1666 ();
 sg13g2_fill_1 FILLER_44_1672 ();
 sg13g2_decap_4 FILLER_44_1685 ();
 sg13g2_fill_1 FILLER_44_1689 ();
 sg13g2_decap_8 FILLER_44_1701 ();
 sg13g2_decap_8 FILLER_44_1708 ();
 sg13g2_fill_1 FILLER_44_1715 ();
 sg13g2_decap_8 FILLER_44_1720 ();
 sg13g2_decap_4 FILLER_44_1727 ();
 sg13g2_fill_2 FILLER_44_1747 ();
 sg13g2_fill_2 FILLER_44_1761 ();
 sg13g2_fill_1 FILLER_44_1763 ();
 sg13g2_decap_8 FILLER_44_1769 ();
 sg13g2_fill_1 FILLER_44_1776 ();
 sg13g2_decap_4 FILLER_44_1786 ();
 sg13g2_fill_2 FILLER_44_1790 ();
 sg13g2_fill_2 FILLER_44_1826 ();
 sg13g2_fill_1 FILLER_44_1828 ();
 sg13g2_decap_4 FILLER_44_1852 ();
 sg13g2_fill_2 FILLER_44_1856 ();
 sg13g2_fill_1 FILLER_44_1861 ();
 sg13g2_fill_1 FILLER_44_1867 ();
 sg13g2_fill_2 FILLER_44_1887 ();
 sg13g2_decap_8 FILLER_44_1894 ();
 sg13g2_fill_2 FILLER_44_1901 ();
 sg13g2_decap_4 FILLER_44_1959 ();
 sg13g2_fill_1 FILLER_44_1963 ();
 sg13g2_decap_8 FILLER_44_1988 ();
 sg13g2_fill_1 FILLER_44_1995 ();
 sg13g2_fill_1 FILLER_44_2005 ();
 sg13g2_decap_8 FILLER_44_2019 ();
 sg13g2_decap_4 FILLER_44_2026 ();
 sg13g2_fill_1 FILLER_44_2067 ();
 sg13g2_fill_2 FILLER_44_2073 ();
 sg13g2_fill_1 FILLER_44_2083 ();
 sg13g2_fill_2 FILLER_44_2108 ();
 sg13g2_fill_2 FILLER_44_2116 ();
 sg13g2_fill_2 FILLER_44_2126 ();
 sg13g2_fill_2 FILLER_44_2141 ();
 sg13g2_fill_1 FILLER_44_2143 ();
 sg13g2_decap_8 FILLER_44_2171 ();
 sg13g2_fill_2 FILLER_44_2178 ();
 sg13g2_decap_4 FILLER_44_2184 ();
 sg13g2_fill_1 FILLER_44_2188 ();
 sg13g2_fill_1 FILLER_44_2208 ();
 sg13g2_fill_1 FILLER_44_2238 ();
 sg13g2_decap_8 FILLER_44_2249 ();
 sg13g2_fill_2 FILLER_44_2256 ();
 sg13g2_decap_4 FILLER_44_2262 ();
 sg13g2_fill_2 FILLER_44_2266 ();
 sg13g2_fill_2 FILLER_44_2273 ();
 sg13g2_decap_8 FILLER_44_2284 ();
 sg13g2_fill_2 FILLER_44_2291 ();
 sg13g2_decap_4 FILLER_44_2298 ();
 sg13g2_fill_1 FILLER_44_2314 ();
 sg13g2_fill_1 FILLER_44_2344 ();
 sg13g2_decap_8 FILLER_44_2376 ();
 sg13g2_decap_4 FILLER_44_2383 ();
 sg13g2_fill_1 FILLER_44_2387 ();
 sg13g2_decap_8 FILLER_44_2396 ();
 sg13g2_decap_4 FILLER_44_2403 ();
 sg13g2_fill_2 FILLER_44_2420 ();
 sg13g2_decap_4 FILLER_44_2427 ();
 sg13g2_fill_2 FILLER_44_2431 ();
 sg13g2_decap_8 FILLER_44_2437 ();
 sg13g2_decap_4 FILLER_44_2444 ();
 sg13g2_decap_8 FILLER_44_2463 ();
 sg13g2_decap_4 FILLER_44_2470 ();
 sg13g2_fill_2 FILLER_44_2479 ();
 sg13g2_decap_8 FILLER_44_2486 ();
 sg13g2_decap_8 FILLER_44_2493 ();
 sg13g2_fill_1 FILLER_44_2508 ();
 sg13g2_fill_1 FILLER_44_2533 ();
 sg13g2_decap_4 FILLER_44_2565 ();
 sg13g2_fill_1 FILLER_44_2595 ();
 sg13g2_decap_8 FILLER_44_2600 ();
 sg13g2_fill_2 FILLER_44_2607 ();
 sg13g2_fill_2 FILLER_44_2627 ();
 sg13g2_decap_8 FILLER_44_2666 ();
 sg13g2_fill_2 FILLER_44_2673 ();
 sg13g2_fill_1 FILLER_44_2675 ();
 sg13g2_decap_8 FILLER_44_2689 ();
 sg13g2_decap_8 FILLER_44_2696 ();
 sg13g2_fill_2 FILLER_44_2703 ();
 sg13g2_decap_8 FILLER_44_2709 ();
 sg13g2_decap_8 FILLER_44_2727 ();
 sg13g2_decap_8 FILLER_44_2734 ();
 sg13g2_decap_8 FILLER_44_2741 ();
 sg13g2_decap_4 FILLER_44_2748 ();
 sg13g2_decap_8 FILLER_44_2755 ();
 sg13g2_decap_8 FILLER_44_2762 ();
 sg13g2_decap_4 FILLER_44_2769 ();
 sg13g2_fill_1 FILLER_44_2773 ();
 sg13g2_fill_2 FILLER_44_2778 ();
 sg13g2_decap_8 FILLER_44_2801 ();
 sg13g2_fill_1 FILLER_44_2808 ();
 sg13g2_decap_8 FILLER_44_2813 ();
 sg13g2_decap_8 FILLER_44_2820 ();
 sg13g2_fill_1 FILLER_44_2827 ();
 sg13g2_decap_8 FILLER_44_2841 ();
 sg13g2_decap_8 FILLER_44_2848 ();
 sg13g2_decap_8 FILLER_44_2855 ();
 sg13g2_decap_8 FILLER_44_2862 ();
 sg13g2_decap_8 FILLER_44_2873 ();
 sg13g2_decap_8 FILLER_44_2880 ();
 sg13g2_decap_8 FILLER_44_2887 ();
 sg13g2_decap_4 FILLER_44_2894 ();
 sg13g2_fill_2 FILLER_44_2898 ();
 sg13g2_fill_1 FILLER_44_2904 ();
 sg13g2_decap_8 FILLER_44_2914 ();
 sg13g2_decap_8 FILLER_44_2921 ();
 sg13g2_decap_8 FILLER_44_2928 ();
 sg13g2_decap_8 FILLER_44_2935 ();
 sg13g2_decap_8 FILLER_44_2942 ();
 sg13g2_decap_8 FILLER_44_2949 ();
 sg13g2_decap_8 FILLER_44_2956 ();
 sg13g2_decap_8 FILLER_44_2963 ();
 sg13g2_fill_1 FILLER_44_2970 ();
 sg13g2_decap_8 FILLER_44_2975 ();
 sg13g2_decap_8 FILLER_44_2982 ();
 sg13g2_decap_8 FILLER_44_2989 ();
 sg13g2_fill_1 FILLER_44_2996 ();
 sg13g2_decap_8 FILLER_44_3003 ();
 sg13g2_decap_8 FILLER_44_3010 ();
 sg13g2_decap_8 FILLER_44_3017 ();
 sg13g2_decap_8 FILLER_44_3024 ();
 sg13g2_decap_8 FILLER_44_3031 ();
 sg13g2_decap_8 FILLER_44_3038 ();
 sg13g2_decap_8 FILLER_44_3045 ();
 sg13g2_decap_8 FILLER_44_3052 ();
 sg13g2_decap_8 FILLER_44_3059 ();
 sg13g2_decap_8 FILLER_44_3066 ();
 sg13g2_decap_8 FILLER_44_3073 ();
 sg13g2_decap_8 FILLER_44_3080 ();
 sg13g2_decap_8 FILLER_44_3087 ();
 sg13g2_decap_8 FILLER_44_3094 ();
 sg13g2_decap_8 FILLER_44_3101 ();
 sg13g2_decap_8 FILLER_44_3108 ();
 sg13g2_decap_8 FILLER_44_3115 ();
 sg13g2_decap_8 FILLER_44_3122 ();
 sg13g2_decap_4 FILLER_44_3129 ();
 sg13g2_decap_8 FILLER_44_3137 ();
 sg13g2_decap_8 FILLER_44_3144 ();
 sg13g2_decap_8 FILLER_44_3151 ();
 sg13g2_decap_8 FILLER_44_3158 ();
 sg13g2_fill_2 FILLER_44_3165 ();
 sg13g2_fill_1 FILLER_44_3167 ();
 sg13g2_decap_8 FILLER_44_3172 ();
 sg13g2_decap_8 FILLER_44_3179 ();
 sg13g2_decap_8 FILLER_44_3186 ();
 sg13g2_decap_8 FILLER_44_3193 ();
 sg13g2_decap_8 FILLER_44_3200 ();
 sg13g2_decap_8 FILLER_44_3207 ();
 sg13g2_decap_8 FILLER_44_3214 ();
 sg13g2_decap_8 FILLER_44_3221 ();
 sg13g2_decap_8 FILLER_44_3228 ();
 sg13g2_decap_8 FILLER_44_3235 ();
 sg13g2_decap_8 FILLER_44_3242 ();
 sg13g2_decap_8 FILLER_44_3249 ();
 sg13g2_decap_8 FILLER_44_3256 ();
 sg13g2_decap_8 FILLER_44_3263 ();
 sg13g2_decap_8 FILLER_44_3270 ();
 sg13g2_decap_8 FILLER_44_3277 ();
 sg13g2_decap_8 FILLER_44_3284 ();
 sg13g2_decap_8 FILLER_44_3291 ();
 sg13g2_decap_8 FILLER_44_3298 ();
 sg13g2_decap_8 FILLER_44_3305 ();
 sg13g2_decap_8 FILLER_44_3312 ();
 sg13g2_decap_8 FILLER_44_3319 ();
 sg13g2_decap_8 FILLER_44_3326 ();
 sg13g2_decap_8 FILLER_44_3333 ();
 sg13g2_decap_8 FILLER_44_3340 ();
 sg13g2_decap_8 FILLER_44_3347 ();
 sg13g2_decap_8 FILLER_44_3354 ();
 sg13g2_decap_8 FILLER_44_3361 ();
 sg13g2_decap_8 FILLER_44_3368 ();
 sg13g2_decap_8 FILLER_44_3375 ();
 sg13g2_decap_8 FILLER_44_3382 ();
 sg13g2_decap_8 FILLER_44_3389 ();
 sg13g2_decap_8 FILLER_44_3396 ();
 sg13g2_decap_8 FILLER_44_3403 ();
 sg13g2_decap_8 FILLER_44_3410 ();
 sg13g2_decap_8 FILLER_44_3417 ();
 sg13g2_decap_8 FILLER_44_3424 ();
 sg13g2_decap_8 FILLER_44_3431 ();
 sg13g2_decap_8 FILLER_44_3438 ();
 sg13g2_decap_8 FILLER_44_3445 ();
 sg13g2_decap_8 FILLER_44_3452 ();
 sg13g2_decap_8 FILLER_44_3459 ();
 sg13g2_decap_8 FILLER_44_3466 ();
 sg13g2_decap_8 FILLER_44_3473 ();
 sg13g2_decap_8 FILLER_44_3480 ();
 sg13g2_decap_8 FILLER_44_3487 ();
 sg13g2_decap_8 FILLER_44_3494 ();
 sg13g2_decap_8 FILLER_44_3501 ();
 sg13g2_decap_8 FILLER_44_3508 ();
 sg13g2_decap_8 FILLER_44_3515 ();
 sg13g2_decap_8 FILLER_44_3522 ();
 sg13g2_decap_8 FILLER_44_3529 ();
 sg13g2_decap_8 FILLER_44_3536 ();
 sg13g2_decap_8 FILLER_44_3543 ();
 sg13g2_decap_8 FILLER_44_3550 ();
 sg13g2_decap_8 FILLER_44_3557 ();
 sg13g2_decap_8 FILLER_44_3564 ();
 sg13g2_decap_8 FILLER_44_3571 ();
 sg13g2_fill_2 FILLER_44_3578 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_4 FILLER_45_7 ();
 sg13g2_fill_2 FILLER_45_11 ();
 sg13g2_decap_8 FILLER_45_17 ();
 sg13g2_fill_1 FILLER_45_24 ();
 sg13g2_fill_1 FILLER_45_65 ();
 sg13g2_decap_4 FILLER_45_85 ();
 sg13g2_fill_2 FILLER_45_89 ();
 sg13g2_decap_4 FILLER_45_117 ();
 sg13g2_fill_1 FILLER_45_121 ();
 sg13g2_fill_1 FILLER_45_200 ();
 sg13g2_fill_1 FILLER_45_221 ();
 sg13g2_fill_2 FILLER_45_283 ();
 sg13g2_fill_1 FILLER_45_311 ();
 sg13g2_decap_4 FILLER_45_328 ();
 sg13g2_fill_2 FILLER_45_357 ();
 sg13g2_fill_1 FILLER_45_359 ();
 sg13g2_fill_1 FILLER_45_391 ();
 sg13g2_fill_1 FILLER_45_424 ();
 sg13g2_fill_2 FILLER_45_452 ();
 sg13g2_decap_4 FILLER_45_480 ();
 sg13g2_fill_1 FILLER_45_484 ();
 sg13g2_fill_2 FILLER_45_564 ();
 sg13g2_decap_4 FILLER_45_592 ();
 sg13g2_fill_1 FILLER_45_596 ();
 sg13g2_decap_4 FILLER_45_607 ();
 sg13g2_fill_1 FILLER_45_611 ();
 sg13g2_decap_4 FILLER_45_627 ();
 sg13g2_fill_2 FILLER_45_631 ();
 sg13g2_fill_2 FILLER_45_654 ();
 sg13g2_fill_2 FILLER_45_669 ();
 sg13g2_fill_1 FILLER_45_697 ();
 sg13g2_fill_2 FILLER_45_711 ();
 sg13g2_fill_1 FILLER_45_713 ();
 sg13g2_fill_2 FILLER_45_740 ();
 sg13g2_fill_1 FILLER_45_742 ();
 sg13g2_fill_1 FILLER_45_773 ();
 sg13g2_fill_2 FILLER_45_802 ();
 sg13g2_fill_1 FILLER_45_817 ();
 sg13g2_fill_2 FILLER_45_826 ();
 sg13g2_fill_1 FILLER_45_834 ();
 sg13g2_fill_1 FILLER_45_840 ();
 sg13g2_decap_8 FILLER_45_846 ();
 sg13g2_fill_1 FILLER_45_853 ();
 sg13g2_decap_8 FILLER_45_858 ();
 sg13g2_decap_8 FILLER_45_865 ();
 sg13g2_fill_1 FILLER_45_872 ();
 sg13g2_fill_2 FILLER_45_912 ();
 sg13g2_fill_1 FILLER_45_942 ();
 sg13g2_decap_4 FILLER_45_961 ();
 sg13g2_decap_4 FILLER_45_969 ();
 sg13g2_fill_2 FILLER_45_973 ();
 sg13g2_fill_1 FILLER_45_979 ();
 sg13g2_fill_1 FILLER_45_984 ();
 sg13g2_decap_4 FILLER_45_995 ();
 sg13g2_fill_2 FILLER_45_999 ();
 sg13g2_fill_2 FILLER_45_1005 ();
 sg13g2_fill_1 FILLER_45_1007 ();
 sg13g2_decap_8 FILLER_45_1012 ();
 sg13g2_decap_8 FILLER_45_1019 ();
 sg13g2_decap_4 FILLER_45_1026 ();
 sg13g2_fill_2 FILLER_45_1067 ();
 sg13g2_decap_8 FILLER_45_1095 ();
 sg13g2_decap_8 FILLER_45_1112 ();
 sg13g2_decap_8 FILLER_45_1119 ();
 sg13g2_decap_8 FILLER_45_1126 ();
 sg13g2_decap_8 FILLER_45_1133 ();
 sg13g2_decap_8 FILLER_45_1144 ();
 sg13g2_fill_2 FILLER_45_1151 ();
 sg13g2_fill_2 FILLER_45_1168 ();
 sg13g2_fill_1 FILLER_45_1178 ();
 sg13g2_fill_2 FILLER_45_1187 ();
 sg13g2_fill_1 FILLER_45_1189 ();
 sg13g2_decap_8 FILLER_45_1237 ();
 sg13g2_decap_8 FILLER_45_1244 ();
 sg13g2_fill_2 FILLER_45_1251 ();
 sg13g2_fill_2 FILLER_45_1270 ();
 sg13g2_fill_1 FILLER_45_1272 ();
 sg13g2_fill_2 FILLER_45_1277 ();
 sg13g2_fill_1 FILLER_45_1279 ();
 sg13g2_fill_2 FILLER_45_1352 ();
 sg13g2_fill_1 FILLER_45_1376 ();
 sg13g2_fill_1 FILLER_45_1383 ();
 sg13g2_fill_2 FILLER_45_1389 ();
 sg13g2_fill_2 FILLER_45_1395 ();
 sg13g2_fill_1 FILLER_45_1407 ();
 sg13g2_fill_1 FILLER_45_1413 ();
 sg13g2_decap_8 FILLER_45_1418 ();
 sg13g2_decap_8 FILLER_45_1425 ();
 sg13g2_decap_4 FILLER_45_1432 ();
 sg13g2_decap_4 FILLER_45_1446 ();
 sg13g2_fill_1 FILLER_45_1450 ();
 sg13g2_decap_4 FILLER_45_1459 ();
 sg13g2_fill_1 FILLER_45_1463 ();
 sg13g2_decap_4 FILLER_45_1470 ();
 sg13g2_fill_2 FILLER_45_1518 ();
 sg13g2_fill_1 FILLER_45_1550 ();
 sg13g2_fill_1 FILLER_45_1557 ();
 sg13g2_fill_2 FILLER_45_1605 ();
 sg13g2_fill_1 FILLER_45_1607 ();
 sg13g2_fill_2 FILLER_45_1648 ();
 sg13g2_decap_8 FILLER_45_1659 ();
 sg13g2_fill_2 FILLER_45_1666 ();
 sg13g2_fill_1 FILLER_45_1668 ();
 sg13g2_fill_1 FILLER_45_1680 ();
 sg13g2_fill_2 FILLER_45_1689 ();
 sg13g2_fill_2 FILLER_45_1711 ();
 sg13g2_fill_2 FILLER_45_1718 ();
 sg13g2_decap_4 FILLER_45_1738 ();
 sg13g2_fill_2 FILLER_45_1742 ();
 sg13g2_decap_8 FILLER_45_1758 ();
 sg13g2_decap_4 FILLER_45_1765 ();
 sg13g2_fill_2 FILLER_45_1791 ();
 sg13g2_decap_8 FILLER_45_1825 ();
 sg13g2_decap_4 FILLER_45_1832 ();
 sg13g2_fill_1 FILLER_45_1849 ();
 sg13g2_fill_2 FILLER_45_1881 ();
 sg13g2_decap_8 FILLER_45_1902 ();
 sg13g2_decap_8 FILLER_45_1909 ();
 sg13g2_fill_1 FILLER_45_1916 ();
 sg13g2_fill_2 FILLER_45_1931 ();
 sg13g2_fill_2 FILLER_45_1942 ();
 sg13g2_fill_1 FILLER_45_1944 ();
 sg13g2_decap_4 FILLER_45_1959 ();
 sg13g2_fill_2 FILLER_45_1977 ();
 sg13g2_decap_4 FILLER_45_1986 ();
 sg13g2_fill_1 FILLER_45_1990 ();
 sg13g2_decap_8 FILLER_45_2022 ();
 sg13g2_fill_2 FILLER_45_2039 ();
 sg13g2_fill_1 FILLER_45_2041 ();
 sg13g2_decap_8 FILLER_45_2057 ();
 sg13g2_fill_2 FILLER_45_2064 ();
 sg13g2_fill_1 FILLER_45_2066 ();
 sg13g2_fill_1 FILLER_45_2080 ();
 sg13g2_fill_2 FILLER_45_2087 ();
 sg13g2_decap_4 FILLER_45_2099 ();
 sg13g2_fill_2 FILLER_45_2103 ();
 sg13g2_fill_1 FILLER_45_2109 ();
 sg13g2_decap_8 FILLER_45_2115 ();
 sg13g2_fill_2 FILLER_45_2122 ();
 sg13g2_decap_4 FILLER_45_2128 ();
 sg13g2_fill_1 FILLER_45_2132 ();
 sg13g2_decap_8 FILLER_45_2137 ();
 sg13g2_decap_8 FILLER_45_2160 ();
 sg13g2_fill_2 FILLER_45_2167 ();
 sg13g2_fill_2 FILLER_45_2209 ();
 sg13g2_fill_1 FILLER_45_2217 ();
 sg13g2_decap_8 FILLER_45_2223 ();
 sg13g2_decap_8 FILLER_45_2230 ();
 sg13g2_decap_4 FILLER_45_2237 ();
 sg13g2_fill_1 FILLER_45_2241 ();
 sg13g2_decap_8 FILLER_45_2257 ();
 sg13g2_fill_1 FILLER_45_2264 ();
 sg13g2_fill_1 FILLER_45_2270 ();
 sg13g2_fill_2 FILLER_45_2291 ();
 sg13g2_fill_1 FILLER_45_2293 ();
 sg13g2_decap_8 FILLER_45_2299 ();
 sg13g2_decap_4 FILLER_45_2306 ();
 sg13g2_fill_1 FILLER_45_2310 ();
 sg13g2_decap_8 FILLER_45_2316 ();
 sg13g2_decap_4 FILLER_45_2323 ();
 sg13g2_fill_2 FILLER_45_2327 ();
 sg13g2_decap_4 FILLER_45_2333 ();
 sg13g2_fill_1 FILLER_45_2337 ();
 sg13g2_decap_8 FILLER_45_2346 ();
 sg13g2_fill_2 FILLER_45_2358 ();
 sg13g2_decap_4 FILLER_45_2364 ();
 sg13g2_fill_1 FILLER_45_2368 ();
 sg13g2_decap_8 FILLER_45_2385 ();
 sg13g2_decap_4 FILLER_45_2392 ();
 sg13g2_fill_2 FILLER_45_2396 ();
 sg13g2_fill_2 FILLER_45_2419 ();
 sg13g2_fill_1 FILLER_45_2421 ();
 sg13g2_decap_4 FILLER_45_2455 ();
 sg13g2_fill_2 FILLER_45_2477 ();
 sg13g2_fill_2 FILLER_45_2493 ();
 sg13g2_decap_4 FILLER_45_2500 ();
 sg13g2_fill_2 FILLER_45_2508 ();
 sg13g2_decap_8 FILLER_45_2526 ();
 sg13g2_decap_8 FILLER_45_2533 ();
 sg13g2_decap_4 FILLER_45_2540 ();
 sg13g2_fill_1 FILLER_45_2549 ();
 sg13g2_decap_8 FILLER_45_2554 ();
 sg13g2_fill_2 FILLER_45_2561 ();
 sg13g2_fill_1 FILLER_45_2563 ();
 sg13g2_fill_2 FILLER_45_2576 ();
 sg13g2_fill_1 FILLER_45_2621 ();
 sg13g2_decap_4 FILLER_45_2638 ();
 sg13g2_fill_1 FILLER_45_2642 ();
 sg13g2_decap_4 FILLER_45_2659 ();
 sg13g2_fill_1 FILLER_45_2663 ();
 sg13g2_fill_2 FILLER_45_2716 ();
 sg13g2_fill_2 FILLER_45_2755 ();
 sg13g2_decap_8 FILLER_45_2821 ();
 sg13g2_decap_8 FILLER_45_2828 ();
 sg13g2_fill_1 FILLER_45_2835 ();
 sg13g2_decap_8 FILLER_45_2840 ();
 sg13g2_fill_2 FILLER_45_2847 ();
 sg13g2_decap_8 FILLER_45_2862 ();
 sg13g2_fill_2 FILLER_45_2869 ();
 sg13g2_decap_8 FILLER_45_2897 ();
 sg13g2_decap_8 FILLER_45_2904 ();
 sg13g2_decap_8 FILLER_45_2911 ();
 sg13g2_decap_8 FILLER_45_2918 ();
 sg13g2_decap_8 FILLER_45_2925 ();
 sg13g2_decap_8 FILLER_45_2932 ();
 sg13g2_decap_8 FILLER_45_2939 ();
 sg13g2_decap_8 FILLER_45_2946 ();
 sg13g2_decap_8 FILLER_45_2953 ();
 sg13g2_decap_8 FILLER_45_2960 ();
 sg13g2_decap_8 FILLER_45_2967 ();
 sg13g2_decap_8 FILLER_45_2974 ();
 sg13g2_decap_8 FILLER_45_2981 ();
 sg13g2_decap_4 FILLER_45_2988 ();
 sg13g2_fill_2 FILLER_45_2992 ();
 sg13g2_decap_8 FILLER_45_3004 ();
 sg13g2_decap_8 FILLER_45_3011 ();
 sg13g2_decap_8 FILLER_45_3018 ();
 sg13g2_decap_8 FILLER_45_3025 ();
 sg13g2_decap_8 FILLER_45_3032 ();
 sg13g2_decap_8 FILLER_45_3039 ();
 sg13g2_decap_8 FILLER_45_3046 ();
 sg13g2_decap_8 FILLER_45_3053 ();
 sg13g2_decap_8 FILLER_45_3060 ();
 sg13g2_decap_8 FILLER_45_3067 ();
 sg13g2_decap_8 FILLER_45_3074 ();
 sg13g2_decap_8 FILLER_45_3081 ();
 sg13g2_decap_8 FILLER_45_3088 ();
 sg13g2_decap_8 FILLER_45_3095 ();
 sg13g2_decap_8 FILLER_45_3102 ();
 sg13g2_decap_8 FILLER_45_3109 ();
 sg13g2_decap_8 FILLER_45_3116 ();
 sg13g2_decap_8 FILLER_45_3123 ();
 sg13g2_decap_8 FILLER_45_3130 ();
 sg13g2_decap_8 FILLER_45_3137 ();
 sg13g2_decap_8 FILLER_45_3144 ();
 sg13g2_decap_8 FILLER_45_3151 ();
 sg13g2_decap_8 FILLER_45_3158 ();
 sg13g2_decap_8 FILLER_45_3165 ();
 sg13g2_decap_8 FILLER_45_3172 ();
 sg13g2_decap_8 FILLER_45_3179 ();
 sg13g2_decap_8 FILLER_45_3186 ();
 sg13g2_decap_8 FILLER_45_3193 ();
 sg13g2_decap_8 FILLER_45_3200 ();
 sg13g2_decap_8 FILLER_45_3207 ();
 sg13g2_decap_8 FILLER_45_3214 ();
 sg13g2_decap_8 FILLER_45_3221 ();
 sg13g2_decap_8 FILLER_45_3228 ();
 sg13g2_decap_8 FILLER_45_3235 ();
 sg13g2_decap_8 FILLER_45_3242 ();
 sg13g2_decap_8 FILLER_45_3249 ();
 sg13g2_decap_8 FILLER_45_3256 ();
 sg13g2_decap_8 FILLER_45_3263 ();
 sg13g2_decap_8 FILLER_45_3270 ();
 sg13g2_decap_8 FILLER_45_3277 ();
 sg13g2_decap_8 FILLER_45_3284 ();
 sg13g2_decap_8 FILLER_45_3291 ();
 sg13g2_decap_8 FILLER_45_3298 ();
 sg13g2_decap_8 FILLER_45_3305 ();
 sg13g2_decap_8 FILLER_45_3312 ();
 sg13g2_decap_8 FILLER_45_3319 ();
 sg13g2_decap_8 FILLER_45_3326 ();
 sg13g2_decap_8 FILLER_45_3333 ();
 sg13g2_decap_8 FILLER_45_3340 ();
 sg13g2_decap_8 FILLER_45_3347 ();
 sg13g2_decap_8 FILLER_45_3354 ();
 sg13g2_decap_8 FILLER_45_3361 ();
 sg13g2_decap_8 FILLER_45_3368 ();
 sg13g2_decap_8 FILLER_45_3375 ();
 sg13g2_decap_8 FILLER_45_3382 ();
 sg13g2_decap_8 FILLER_45_3389 ();
 sg13g2_decap_8 FILLER_45_3396 ();
 sg13g2_decap_8 FILLER_45_3403 ();
 sg13g2_decap_8 FILLER_45_3410 ();
 sg13g2_decap_8 FILLER_45_3417 ();
 sg13g2_decap_8 FILLER_45_3424 ();
 sg13g2_decap_8 FILLER_45_3431 ();
 sg13g2_decap_8 FILLER_45_3438 ();
 sg13g2_decap_8 FILLER_45_3445 ();
 sg13g2_decap_8 FILLER_45_3452 ();
 sg13g2_decap_8 FILLER_45_3459 ();
 sg13g2_decap_8 FILLER_45_3466 ();
 sg13g2_decap_8 FILLER_45_3473 ();
 sg13g2_decap_8 FILLER_45_3480 ();
 sg13g2_decap_8 FILLER_45_3487 ();
 sg13g2_decap_8 FILLER_45_3494 ();
 sg13g2_decap_8 FILLER_45_3501 ();
 sg13g2_decap_8 FILLER_45_3508 ();
 sg13g2_decap_8 FILLER_45_3515 ();
 sg13g2_decap_8 FILLER_45_3522 ();
 sg13g2_decap_8 FILLER_45_3529 ();
 sg13g2_decap_8 FILLER_45_3536 ();
 sg13g2_decap_8 FILLER_45_3543 ();
 sg13g2_decap_8 FILLER_45_3550 ();
 sg13g2_decap_8 FILLER_45_3557 ();
 sg13g2_decap_8 FILLER_45_3564 ();
 sg13g2_decap_8 FILLER_45_3571 ();
 sg13g2_fill_2 FILLER_45_3578 ();
 sg13g2_fill_2 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_28 ();
 sg13g2_fill_1 FILLER_46_43 ();
 sg13g2_decap_8 FILLER_46_66 ();
 sg13g2_decap_8 FILLER_46_78 ();
 sg13g2_decap_8 FILLER_46_85 ();
 sg13g2_fill_2 FILLER_46_92 ();
 sg13g2_fill_2 FILLER_46_99 ();
 sg13g2_fill_1 FILLER_46_101 ();
 sg13g2_decap_8 FILLER_46_106 ();
 sg13g2_fill_1 FILLER_46_113 ();
 sg13g2_decap_4 FILLER_46_129 ();
 sg13g2_fill_2 FILLER_46_146 ();
 sg13g2_fill_1 FILLER_46_148 ();
 sg13g2_fill_2 FILLER_46_172 ();
 sg13g2_fill_1 FILLER_46_174 ();
 sg13g2_fill_2 FILLER_46_178 ();
 sg13g2_decap_4 FILLER_46_223 ();
 sg13g2_fill_2 FILLER_46_236 ();
 sg13g2_fill_1 FILLER_46_242 ();
 sg13g2_decap_4 FILLER_46_248 ();
 sg13g2_fill_2 FILLER_46_252 ();
 sg13g2_fill_1 FILLER_46_263 ();
 sg13g2_fill_2 FILLER_46_271 ();
 sg13g2_fill_2 FILLER_46_310 ();
 sg13g2_fill_1 FILLER_46_312 ();
 sg13g2_fill_2 FILLER_46_322 ();
 sg13g2_fill_1 FILLER_46_324 ();
 sg13g2_decap_8 FILLER_46_328 ();
 sg13g2_decap_8 FILLER_46_335 ();
 sg13g2_fill_2 FILLER_46_369 ();
 sg13g2_fill_1 FILLER_46_380 ();
 sg13g2_fill_2 FILLER_46_404 ();
 sg13g2_decap_8 FILLER_46_415 ();
 sg13g2_fill_2 FILLER_46_422 ();
 sg13g2_fill_1 FILLER_46_424 ();
 sg13g2_fill_2 FILLER_46_475 ();
 sg13g2_fill_1 FILLER_46_507 ();
 sg13g2_decap_8 FILLER_46_529 ();
 sg13g2_decap_4 FILLER_46_536 ();
 sg13g2_fill_2 FILLER_46_548 ();
 sg13g2_decap_8 FILLER_46_554 ();
 sg13g2_fill_1 FILLER_46_566 ();
 sg13g2_decap_4 FILLER_46_571 ();
 sg13g2_fill_1 FILLER_46_575 ();
 sg13g2_fill_2 FILLER_46_593 ();
 sg13g2_fill_1 FILLER_46_595 ();
 sg13g2_fill_2 FILLER_46_601 ();
 sg13g2_decap_4 FILLER_46_611 ();
 sg13g2_fill_1 FILLER_46_615 ();
 sg13g2_fill_2 FILLER_46_628 ();
 sg13g2_fill_1 FILLER_46_656 ();
 sg13g2_fill_2 FILLER_46_671 ();
 sg13g2_fill_1 FILLER_46_673 ();
 sg13g2_fill_2 FILLER_46_696 ();
 sg13g2_fill_2 FILLER_46_712 ();
 sg13g2_fill_1 FILLER_46_714 ();
 sg13g2_fill_2 FILLER_46_725 ();
 sg13g2_fill_1 FILLER_46_727 ();
 sg13g2_fill_2 FILLER_46_737 ();
 sg13g2_fill_2 FILLER_46_757 ();
 sg13g2_fill_2 FILLER_46_768 ();
 sg13g2_fill_1 FILLER_46_770 ();
 sg13g2_decap_4 FILLER_46_776 ();
 sg13g2_fill_1 FILLER_46_806 ();
 sg13g2_fill_1 FILLER_46_815 ();
 sg13g2_fill_1 FILLER_46_833 ();
 sg13g2_fill_2 FILLER_46_852 ();
 sg13g2_fill_1 FILLER_46_854 ();
 sg13g2_decap_4 FILLER_46_860 ();
 sg13g2_fill_1 FILLER_46_864 ();
 sg13g2_decap_4 FILLER_46_873 ();
 sg13g2_decap_4 FILLER_46_898 ();
 sg13g2_fill_2 FILLER_46_902 ();
 sg13g2_fill_1 FILLER_46_929 ();
 sg13g2_decap_8 FILLER_46_941 ();
 sg13g2_fill_1 FILLER_46_953 ();
 sg13g2_fill_1 FILLER_46_980 ();
 sg13g2_fill_1 FILLER_46_996 ();
 sg13g2_fill_2 FILLER_46_1028 ();
 sg13g2_fill_1 FILLER_46_1030 ();
 sg13g2_fill_1 FILLER_46_1079 ();
 sg13g2_decap_4 FILLER_46_1084 ();
 sg13g2_fill_1 FILLER_46_1088 ();
 sg13g2_fill_1 FILLER_46_1094 ();
 sg13g2_decap_8 FILLER_46_1121 ();
 sg13g2_fill_1 FILLER_46_1128 ();
 sg13g2_decap_4 FILLER_46_1155 ();
 sg13g2_decap_4 FILLER_46_1172 ();
 sg13g2_fill_1 FILLER_46_1176 ();
 sg13g2_decap_8 FILLER_46_1190 ();
 sg13g2_fill_2 FILLER_46_1197 ();
 sg13g2_fill_1 FILLER_46_1199 ();
 sg13g2_fill_2 FILLER_46_1204 ();
 sg13g2_decap_8 FILLER_46_1214 ();
 sg13g2_fill_2 FILLER_46_1221 ();
 sg13g2_fill_1 FILLER_46_1223 ();
 sg13g2_decap_8 FILLER_46_1229 ();
 sg13g2_decap_4 FILLER_46_1236 ();
 sg13g2_fill_2 FILLER_46_1240 ();
 sg13g2_fill_1 FILLER_46_1282 ();
 sg13g2_decap_8 FILLER_46_1291 ();
 sg13g2_decap_8 FILLER_46_1298 ();
 sg13g2_fill_2 FILLER_46_1305 ();
 sg13g2_decap_4 FILLER_46_1311 ();
 sg13g2_fill_1 FILLER_46_1324 ();
 sg13g2_fill_1 FILLER_46_1357 ();
 sg13g2_fill_2 FILLER_46_1371 ();
 sg13g2_decap_8 FILLER_46_1377 ();
 sg13g2_fill_2 FILLER_46_1387 ();
 sg13g2_fill_2 FILLER_46_1402 ();
 sg13g2_decap_4 FILLER_46_1424 ();
 sg13g2_fill_1 FILLER_46_1428 ();
 sg13g2_decap_4 FILLER_46_1455 ();
 sg13g2_fill_1 FILLER_46_1459 ();
 sg13g2_fill_1 FILLER_46_1464 ();
 sg13g2_decap_8 FILLER_46_1479 ();
 sg13g2_decap_8 FILLER_46_1486 ();
 sg13g2_decap_8 FILLER_46_1493 ();
 sg13g2_fill_1 FILLER_46_1500 ();
 sg13g2_decap_4 FILLER_46_1513 ();
 sg13g2_fill_1 FILLER_46_1517 ();
 sg13g2_fill_2 FILLER_46_1534 ();
 sg13g2_fill_2 FILLER_46_1540 ();
 sg13g2_fill_2 FILLER_46_1551 ();
 sg13g2_decap_4 FILLER_46_1563 ();
 sg13g2_fill_2 FILLER_46_1567 ();
 sg13g2_fill_2 FILLER_46_1574 ();
 sg13g2_decap_8 FILLER_46_1579 ();
 sg13g2_decap_4 FILLER_46_1586 ();
 sg13g2_decap_4 FILLER_46_1594 ();
 sg13g2_fill_1 FILLER_46_1598 ();
 sg13g2_decap_8 FILLER_46_1612 ();
 sg13g2_decap_8 FILLER_46_1623 ();
 sg13g2_decap_4 FILLER_46_1630 ();
 sg13g2_fill_2 FILLER_46_1643 ();
 sg13g2_decap_8 FILLER_46_1657 ();
 sg13g2_decap_8 FILLER_46_1664 ();
 sg13g2_fill_1 FILLER_46_1671 ();
 sg13g2_fill_2 FILLER_46_1686 ();
 sg13g2_fill_2 FILLER_46_1713 ();
 sg13g2_decap_4 FILLER_46_1718 ();
 sg13g2_fill_2 FILLER_46_1722 ();
 sg13g2_decap_8 FILLER_46_1737 ();
 sg13g2_fill_1 FILLER_46_1744 ();
 sg13g2_decap_8 FILLER_46_1769 ();
 sg13g2_decap_8 FILLER_46_1787 ();
 sg13g2_fill_1 FILLER_46_1794 ();
 sg13g2_decap_4 FILLER_46_1819 ();
 sg13g2_decap_4 FILLER_46_1833 ();
 sg13g2_fill_2 FILLER_46_1837 ();
 sg13g2_decap_8 FILLER_46_1844 ();
 sg13g2_fill_2 FILLER_46_1851 ();
 sg13g2_fill_1 FILLER_46_1853 ();
 sg13g2_fill_2 FILLER_46_1858 ();
 sg13g2_fill_2 FILLER_46_1869 ();
 sg13g2_fill_1 FILLER_46_1882 ();
 sg13g2_fill_1 FILLER_46_1898 ();
 sg13g2_decap_4 FILLER_46_1912 ();
 sg13g2_fill_2 FILLER_46_1916 ();
 sg13g2_fill_2 FILLER_46_1966 ();
 sg13g2_fill_1 FILLER_46_1986 ();
 sg13g2_decap_8 FILLER_46_1995 ();
 sg13g2_decap_4 FILLER_46_2002 ();
 sg13g2_decap_8 FILLER_46_2014 ();
 sg13g2_fill_2 FILLER_46_2021 ();
 sg13g2_fill_1 FILLER_46_2031 ();
 sg13g2_fill_2 FILLER_46_2042 ();
 sg13g2_fill_1 FILLER_46_2044 ();
 sg13g2_fill_2 FILLER_46_2055 ();
 sg13g2_fill_1 FILLER_46_2057 ();
 sg13g2_fill_2 FILLER_46_2072 ();
 sg13g2_fill_2 FILLER_46_2079 ();
 sg13g2_fill_1 FILLER_46_2081 ();
 sg13g2_fill_2 FILLER_46_2088 ();
 sg13g2_fill_1 FILLER_46_2090 ();
 sg13g2_fill_2 FILLER_46_2100 ();
 sg13g2_fill_1 FILLER_46_2107 ();
 sg13g2_fill_1 FILLER_46_2113 ();
 sg13g2_decap_8 FILLER_46_2123 ();
 sg13g2_fill_2 FILLER_46_2130 ();
 sg13g2_decap_4 FILLER_46_2136 ();
 sg13g2_decap_4 FILLER_46_2145 ();
 sg13g2_fill_1 FILLER_46_2149 ();
 sg13g2_decap_4 FILLER_46_2155 ();
 sg13g2_fill_2 FILLER_46_2159 ();
 sg13g2_fill_2 FILLER_46_2165 ();
 sg13g2_fill_1 FILLER_46_2167 ();
 sg13g2_decap_8 FILLER_46_2173 ();
 sg13g2_decap_8 FILLER_46_2180 ();
 sg13g2_fill_2 FILLER_46_2187 ();
 sg13g2_fill_1 FILLER_46_2189 ();
 sg13g2_decap_4 FILLER_46_2198 ();
 sg13g2_fill_1 FILLER_46_2202 ();
 sg13g2_decap_8 FILLER_46_2207 ();
 sg13g2_decap_4 FILLER_46_2214 ();
 sg13g2_fill_1 FILLER_46_2245 ();
 sg13g2_fill_1 FILLER_46_2260 ();
 sg13g2_fill_2 FILLER_46_2270 ();
 sg13g2_fill_1 FILLER_46_2272 ();
 sg13g2_decap_8 FILLER_46_2286 ();
 sg13g2_fill_2 FILLER_46_2293 ();
 sg13g2_fill_1 FILLER_46_2295 ();
 sg13g2_fill_2 FILLER_46_2301 ();
 sg13g2_decap_4 FILLER_46_2311 ();
 sg13g2_fill_2 FILLER_46_2315 ();
 sg13g2_fill_2 FILLER_46_2326 ();
 sg13g2_fill_1 FILLER_46_2328 ();
 sg13g2_fill_2 FILLER_46_2338 ();
 sg13g2_fill_1 FILLER_46_2340 ();
 sg13g2_fill_1 FILLER_46_2345 ();
 sg13g2_decap_8 FILLER_46_2355 ();
 sg13g2_fill_1 FILLER_46_2362 ();
 sg13g2_fill_1 FILLER_46_2397 ();
 sg13g2_decap_4 FILLER_46_2415 ();
 sg13g2_fill_1 FILLER_46_2419 ();
 sg13g2_decap_8 FILLER_46_2429 ();
 sg13g2_fill_1 FILLER_46_2436 ();
 sg13g2_fill_2 FILLER_46_2446 ();
 sg13g2_fill_1 FILLER_46_2448 ();
 sg13g2_decap_4 FILLER_46_2484 ();
 sg13g2_fill_2 FILLER_46_2488 ();
 sg13g2_fill_2 FILLER_46_2525 ();
 sg13g2_decap_8 FILLER_46_2531 ();
 sg13g2_decap_4 FILLER_46_2538 ();
 sg13g2_fill_2 FILLER_46_2542 ();
 sg13g2_decap_8 FILLER_46_2584 ();
 sg13g2_decap_4 FILLER_46_2591 ();
 sg13g2_fill_2 FILLER_46_2595 ();
 sg13g2_fill_2 FILLER_46_2601 ();
 sg13g2_decap_4 FILLER_46_2631 ();
 sg13g2_decap_8 FILLER_46_2661 ();
 sg13g2_decap_8 FILLER_46_2668 ();
 sg13g2_fill_2 FILLER_46_2679 ();
 sg13g2_fill_1 FILLER_46_2681 ();
 sg13g2_fill_2 FILLER_46_2687 ();
 sg13g2_fill_1 FILLER_46_2689 ();
 sg13g2_fill_2 FILLER_46_2714 ();
 sg13g2_fill_2 FILLER_46_2729 ();
 sg13g2_fill_1 FILLER_46_2731 ();
 sg13g2_fill_2 FILLER_46_2750 ();
 sg13g2_decap_8 FILLER_46_2755 ();
 sg13g2_fill_1 FILLER_46_2762 ();
 sg13g2_fill_2 FILLER_46_2822 ();
 sg13g2_fill_1 FILLER_46_2824 ();
 sg13g2_fill_2 FILLER_46_2851 ();
 sg13g2_decap_4 FILLER_46_2866 ();
 sg13g2_fill_1 FILLER_46_2870 ();
 sg13g2_fill_1 FILLER_46_2884 ();
 sg13g2_decap_8 FILLER_46_2893 ();
 sg13g2_decap_8 FILLER_46_2900 ();
 sg13g2_decap_8 FILLER_46_2907 ();
 sg13g2_fill_1 FILLER_46_2914 ();
 sg13g2_decap_8 FILLER_46_2919 ();
 sg13g2_fill_2 FILLER_46_2926 ();
 sg13g2_decap_8 FILLER_46_2933 ();
 sg13g2_decap_8 FILLER_46_2940 ();
 sg13g2_decap_8 FILLER_46_2947 ();
 sg13g2_decap_8 FILLER_46_2954 ();
 sg13g2_decap_8 FILLER_46_2961 ();
 sg13g2_decap_8 FILLER_46_2968 ();
 sg13g2_decap_8 FILLER_46_2975 ();
 sg13g2_decap_8 FILLER_46_2982 ();
 sg13g2_decap_8 FILLER_46_2989 ();
 sg13g2_decap_8 FILLER_46_2996 ();
 sg13g2_decap_8 FILLER_46_3003 ();
 sg13g2_decap_8 FILLER_46_3010 ();
 sg13g2_decap_8 FILLER_46_3017 ();
 sg13g2_decap_8 FILLER_46_3024 ();
 sg13g2_decap_8 FILLER_46_3031 ();
 sg13g2_decap_8 FILLER_46_3038 ();
 sg13g2_decap_8 FILLER_46_3045 ();
 sg13g2_decap_8 FILLER_46_3052 ();
 sg13g2_decap_8 FILLER_46_3059 ();
 sg13g2_decap_8 FILLER_46_3066 ();
 sg13g2_decap_8 FILLER_46_3073 ();
 sg13g2_decap_8 FILLER_46_3080 ();
 sg13g2_decap_8 FILLER_46_3087 ();
 sg13g2_decap_8 FILLER_46_3094 ();
 sg13g2_decap_8 FILLER_46_3101 ();
 sg13g2_decap_8 FILLER_46_3108 ();
 sg13g2_decap_8 FILLER_46_3115 ();
 sg13g2_decap_8 FILLER_46_3122 ();
 sg13g2_decap_8 FILLER_46_3129 ();
 sg13g2_decap_8 FILLER_46_3136 ();
 sg13g2_decap_8 FILLER_46_3143 ();
 sg13g2_decap_8 FILLER_46_3150 ();
 sg13g2_decap_8 FILLER_46_3157 ();
 sg13g2_decap_8 FILLER_46_3164 ();
 sg13g2_decap_8 FILLER_46_3171 ();
 sg13g2_decap_8 FILLER_46_3178 ();
 sg13g2_decap_8 FILLER_46_3185 ();
 sg13g2_decap_8 FILLER_46_3192 ();
 sg13g2_decap_8 FILLER_46_3199 ();
 sg13g2_decap_8 FILLER_46_3206 ();
 sg13g2_decap_8 FILLER_46_3213 ();
 sg13g2_decap_8 FILLER_46_3220 ();
 sg13g2_decap_8 FILLER_46_3227 ();
 sg13g2_decap_8 FILLER_46_3234 ();
 sg13g2_decap_8 FILLER_46_3241 ();
 sg13g2_decap_8 FILLER_46_3248 ();
 sg13g2_decap_8 FILLER_46_3255 ();
 sg13g2_decap_8 FILLER_46_3262 ();
 sg13g2_decap_8 FILLER_46_3269 ();
 sg13g2_decap_8 FILLER_46_3276 ();
 sg13g2_decap_8 FILLER_46_3283 ();
 sg13g2_decap_8 FILLER_46_3290 ();
 sg13g2_decap_8 FILLER_46_3297 ();
 sg13g2_decap_8 FILLER_46_3304 ();
 sg13g2_decap_8 FILLER_46_3311 ();
 sg13g2_decap_8 FILLER_46_3318 ();
 sg13g2_decap_8 FILLER_46_3325 ();
 sg13g2_decap_8 FILLER_46_3332 ();
 sg13g2_decap_8 FILLER_46_3339 ();
 sg13g2_decap_8 FILLER_46_3346 ();
 sg13g2_decap_8 FILLER_46_3353 ();
 sg13g2_decap_8 FILLER_46_3360 ();
 sg13g2_decap_8 FILLER_46_3367 ();
 sg13g2_decap_8 FILLER_46_3374 ();
 sg13g2_decap_8 FILLER_46_3381 ();
 sg13g2_decap_8 FILLER_46_3388 ();
 sg13g2_decap_8 FILLER_46_3395 ();
 sg13g2_decap_8 FILLER_46_3402 ();
 sg13g2_decap_8 FILLER_46_3409 ();
 sg13g2_decap_8 FILLER_46_3416 ();
 sg13g2_decap_8 FILLER_46_3423 ();
 sg13g2_decap_8 FILLER_46_3430 ();
 sg13g2_decap_8 FILLER_46_3437 ();
 sg13g2_decap_8 FILLER_46_3444 ();
 sg13g2_decap_8 FILLER_46_3451 ();
 sg13g2_decap_8 FILLER_46_3458 ();
 sg13g2_decap_8 FILLER_46_3465 ();
 sg13g2_decap_8 FILLER_46_3472 ();
 sg13g2_decap_8 FILLER_46_3479 ();
 sg13g2_decap_8 FILLER_46_3486 ();
 sg13g2_decap_8 FILLER_46_3493 ();
 sg13g2_decap_8 FILLER_46_3500 ();
 sg13g2_decap_8 FILLER_46_3507 ();
 sg13g2_decap_8 FILLER_46_3514 ();
 sg13g2_decap_8 FILLER_46_3521 ();
 sg13g2_decap_8 FILLER_46_3528 ();
 sg13g2_decap_8 FILLER_46_3535 ();
 sg13g2_decap_8 FILLER_46_3542 ();
 sg13g2_decap_8 FILLER_46_3549 ();
 sg13g2_decap_8 FILLER_46_3556 ();
 sg13g2_decap_8 FILLER_46_3563 ();
 sg13g2_decap_8 FILLER_46_3570 ();
 sg13g2_fill_2 FILLER_46_3577 ();
 sg13g2_fill_1 FILLER_46_3579 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_4 FILLER_47_7 ();
 sg13g2_fill_2 FILLER_47_11 ();
 sg13g2_decap_4 FILLER_47_17 ();
 sg13g2_fill_1 FILLER_47_21 ();
 sg13g2_fill_1 FILLER_47_43 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_fill_1 FILLER_47_91 ();
 sg13g2_fill_2 FILLER_47_141 ();
 sg13g2_decap_8 FILLER_47_215 ();
 sg13g2_decap_8 FILLER_47_222 ();
 sg13g2_decap_4 FILLER_47_229 ();
 sg13g2_fill_1 FILLER_47_233 ();
 sg13g2_fill_1 FILLER_47_239 ();
 sg13g2_decap_8 FILLER_47_252 ();
 sg13g2_fill_2 FILLER_47_259 ();
 sg13g2_fill_1 FILLER_47_261 ();
 sg13g2_fill_1 FILLER_47_272 ();
 sg13g2_fill_2 FILLER_47_281 ();
 sg13g2_decap_4 FILLER_47_288 ();
 sg13g2_fill_1 FILLER_47_292 ();
 sg13g2_fill_2 FILLER_47_329 ();
 sg13g2_fill_1 FILLER_47_339 ();
 sg13g2_fill_2 FILLER_47_343 ();
 sg13g2_fill_1 FILLER_47_345 ();
 sg13g2_fill_2 FILLER_47_355 ();
 sg13g2_fill_1 FILLER_47_366 ();
 sg13g2_fill_1 FILLER_47_471 ();
 sg13g2_decap_8 FILLER_47_480 ();
 sg13g2_decap_8 FILLER_47_496 ();
 sg13g2_decap_4 FILLER_47_503 ();
 sg13g2_fill_2 FILLER_47_528 ();
 sg13g2_fill_1 FILLER_47_530 ();
 sg13g2_fill_1 FILLER_47_567 ();
 sg13g2_fill_1 FILLER_47_573 ();
 sg13g2_decap_4 FILLER_47_603 ();
 sg13g2_fill_2 FILLER_47_620 ();
 sg13g2_decap_4 FILLER_47_626 ();
 sg13g2_fill_1 FILLER_47_630 ();
 sg13g2_fill_2 FILLER_47_714 ();
 sg13g2_fill_2 FILLER_47_735 ();
 sg13g2_fill_1 FILLER_47_737 ();
 sg13g2_fill_1 FILLER_47_751 ();
 sg13g2_fill_1 FILLER_47_757 ();
 sg13g2_fill_1 FILLER_47_762 ();
 sg13g2_fill_1 FILLER_47_773 ();
 sg13g2_decap_8 FILLER_47_784 ();
 sg13g2_fill_2 FILLER_47_791 ();
 sg13g2_fill_1 FILLER_47_793 ();
 sg13g2_fill_2 FILLER_47_820 ();
 sg13g2_decap_4 FILLER_47_847 ();
 sg13g2_decap_4 FILLER_47_867 ();
 sg13g2_fill_1 FILLER_47_871 ();
 sg13g2_fill_1 FILLER_47_884 ();
 sg13g2_fill_2 FILLER_47_907 ();
 sg13g2_decap_4 FILLER_47_953 ();
 sg13g2_fill_2 FILLER_47_957 ();
 sg13g2_fill_1 FILLER_47_976 ();
 sg13g2_fill_1 FILLER_47_991 ();
 sg13g2_fill_2 FILLER_47_1006 ();
 sg13g2_fill_1 FILLER_47_1008 ();
 sg13g2_decap_8 FILLER_47_1083 ();
 sg13g2_fill_1 FILLER_47_1090 ();
 sg13g2_decap_4 FILLER_47_1101 ();
 sg13g2_fill_1 FILLER_47_1105 ();
 sg13g2_decap_4 FILLER_47_1121 ();
 sg13g2_fill_1 FILLER_47_1125 ();
 sg13g2_decap_4 FILLER_47_1156 ();
 sg13g2_fill_2 FILLER_47_1160 ();
 sg13g2_fill_1 FILLER_47_1214 ();
 sg13g2_fill_1 FILLER_47_1229 ();
 sg13g2_fill_2 FILLER_47_1238 ();
 sg13g2_fill_1 FILLER_47_1240 ();
 sg13g2_decap_8 FILLER_47_1246 ();
 sg13g2_decap_8 FILLER_47_1261 ();
 sg13g2_decap_8 FILLER_47_1268 ();
 sg13g2_fill_2 FILLER_47_1275 ();
 sg13g2_fill_1 FILLER_47_1277 ();
 sg13g2_fill_2 FILLER_47_1282 ();
 sg13g2_fill_2 FILLER_47_1333 ();
 sg13g2_fill_1 FILLER_47_1335 ();
 sg13g2_fill_2 FILLER_47_1351 ();
 sg13g2_fill_1 FILLER_47_1384 ();
 sg13g2_decap_8 FILLER_47_1389 ();
 sg13g2_decap_8 FILLER_47_1396 ();
 sg13g2_decap_4 FILLER_47_1403 ();
 sg13g2_fill_2 FILLER_47_1412 ();
 sg13g2_fill_1 FILLER_47_1414 ();
 sg13g2_decap_4 FILLER_47_1420 ();
 sg13g2_decap_8 FILLER_47_1429 ();
 sg13g2_decap_8 FILLER_47_1436 ();
 sg13g2_fill_2 FILLER_47_1448 ();
 sg13g2_fill_1 FILLER_47_1460 ();
 sg13g2_fill_2 FILLER_47_1501 ();
 sg13g2_decap_8 FILLER_47_1511 ();
 sg13g2_fill_2 FILLER_47_1530 ();
 sg13g2_decap_8 FILLER_47_1567 ();
 sg13g2_fill_2 FILLER_47_1574 ();
 sg13g2_decap_4 FILLER_47_1621 ();
 sg13g2_fill_1 FILLER_47_1635 ();
 sg13g2_fill_2 FILLER_47_1646 ();
 sg13g2_fill_1 FILLER_47_1654 ();
 sg13g2_decap_4 FILLER_47_1664 ();
 sg13g2_fill_2 FILLER_47_1668 ();
 sg13g2_fill_2 FILLER_47_1685 ();
 sg13g2_fill_1 FILLER_47_1687 ();
 sg13g2_decap_4 FILLER_47_1691 ();
 sg13g2_fill_1 FILLER_47_1695 ();
 sg13g2_fill_1 FILLER_47_1706 ();
 sg13g2_fill_1 FILLER_47_1726 ();
 sg13g2_fill_2 FILLER_47_1745 ();
 sg13g2_decap_4 FILLER_47_1764 ();
 sg13g2_decap_8 FILLER_47_1778 ();
 sg13g2_decap_8 FILLER_47_1785 ();
 sg13g2_decap_4 FILLER_47_1792 ();
 sg13g2_fill_1 FILLER_47_1796 ();
 sg13g2_fill_1 FILLER_47_1805 ();
 sg13g2_decap_4 FILLER_47_1815 ();
 sg13g2_fill_2 FILLER_47_1819 ();
 sg13g2_fill_2 FILLER_47_1866 ();
 sg13g2_fill_1 FILLER_47_1868 ();
 sg13g2_fill_2 FILLER_47_1895 ();
 sg13g2_fill_1 FILLER_47_1897 ();
 sg13g2_decap_4 FILLER_47_1919 ();
 sg13g2_decap_4 FILLER_47_1956 ();
 sg13g2_fill_2 FILLER_47_1960 ();
 sg13g2_fill_2 FILLER_47_1973 ();
 sg13g2_decap_4 FILLER_47_1978 ();
 sg13g2_fill_1 FILLER_47_1982 ();
 sg13g2_decap_4 FILLER_47_1988 ();
 sg13g2_decap_8 FILLER_47_2000 ();
 sg13g2_decap_4 FILLER_47_2007 ();
 sg13g2_fill_1 FILLER_47_2011 ();
 sg13g2_fill_1 FILLER_47_2020 ();
 sg13g2_fill_2 FILLER_47_2026 ();
 sg13g2_fill_1 FILLER_47_2028 ();
 sg13g2_fill_1 FILLER_47_2042 ();
 sg13g2_decap_4 FILLER_47_2053 ();
 sg13g2_fill_1 FILLER_47_2057 ();
 sg13g2_decap_4 FILLER_47_2070 ();
 sg13g2_fill_1 FILLER_47_2074 ();
 sg13g2_fill_2 FILLER_47_2083 ();
 sg13g2_fill_1 FILLER_47_2085 ();
 sg13g2_fill_2 FILLER_47_2094 ();
 sg13g2_fill_2 FILLER_47_2100 ();
 sg13g2_fill_1 FILLER_47_2102 ();
 sg13g2_fill_2 FILLER_47_2118 ();
 sg13g2_fill_2 FILLER_47_2163 ();
 sg13g2_decap_4 FILLER_47_2179 ();
 sg13g2_fill_1 FILLER_47_2202 ();
 sg13g2_decap_8 FILLER_47_2226 ();
 sg13g2_decap_8 FILLER_47_2237 ();
 sg13g2_decap_4 FILLER_47_2256 ();
 sg13g2_fill_1 FILLER_47_2260 ();
 sg13g2_decap_4 FILLER_47_2281 ();
 sg13g2_fill_2 FILLER_47_2285 ();
 sg13g2_decap_8 FILLER_47_2292 ();
 sg13g2_fill_2 FILLER_47_2299 ();
 sg13g2_decap_4 FILLER_47_2316 ();
 sg13g2_fill_2 FILLER_47_2328 ();
 sg13g2_fill_1 FILLER_47_2330 ();
 sg13g2_fill_1 FILLER_47_2357 ();
 sg13g2_fill_1 FILLER_47_2379 ();
 sg13g2_fill_2 FILLER_47_2396 ();
 sg13g2_decap_8 FILLER_47_2413 ();
 sg13g2_decap_4 FILLER_47_2420 ();
 sg13g2_fill_2 FILLER_47_2424 ();
 sg13g2_decap_4 FILLER_47_2431 ();
 sg13g2_fill_1 FILLER_47_2435 ();
 sg13g2_decap_8 FILLER_47_2461 ();
 sg13g2_fill_2 FILLER_47_2468 ();
 sg13g2_decap_8 FILLER_47_2500 ();
 sg13g2_fill_1 FILLER_47_2515 ();
 sg13g2_fill_1 FILLER_47_2542 ();
 sg13g2_fill_2 FILLER_47_2551 ();
 sg13g2_decap_4 FILLER_47_2561 ();
 sg13g2_fill_1 FILLER_47_2565 ();
 sg13g2_decap_4 FILLER_47_2591 ();
 sg13g2_fill_2 FILLER_47_2595 ();
 sg13g2_decap_8 FILLER_47_2628 ();
 sg13g2_fill_2 FILLER_47_2635 ();
 sg13g2_fill_1 FILLER_47_2637 ();
 sg13g2_decap_4 FILLER_47_2643 ();
 sg13g2_fill_1 FILLER_47_2647 ();
 sg13g2_fill_2 FILLER_47_2652 ();
 sg13g2_fill_1 FILLER_47_2654 ();
 sg13g2_fill_2 FILLER_47_2663 ();
 sg13g2_decap_4 FILLER_47_2670 ();
 sg13g2_fill_2 FILLER_47_2685 ();
 sg13g2_fill_2 FILLER_47_2804 ();
 sg13g2_fill_1 FILLER_47_2827 ();
 sg13g2_decap_4 FILLER_47_2842 ();
 sg13g2_decap_4 FILLER_47_2865 ();
 sg13g2_decap_4 FILLER_47_2879 ();
 sg13g2_decap_4 FILLER_47_2901 ();
 sg13g2_fill_2 FILLER_47_2920 ();
 sg13g2_fill_1 FILLER_47_2922 ();
 sg13g2_fill_2 FILLER_47_2928 ();
 sg13g2_fill_1 FILLER_47_2930 ();
 sg13g2_fill_2 FILLER_47_2940 ();
 sg13g2_decap_8 FILLER_47_2946 ();
 sg13g2_decap_8 FILLER_47_2953 ();
 sg13g2_decap_8 FILLER_47_2960 ();
 sg13g2_decap_8 FILLER_47_2967 ();
 sg13g2_decap_8 FILLER_47_2974 ();
 sg13g2_decap_8 FILLER_47_2981 ();
 sg13g2_decap_8 FILLER_47_2988 ();
 sg13g2_decap_8 FILLER_47_2995 ();
 sg13g2_decap_8 FILLER_47_3002 ();
 sg13g2_decap_8 FILLER_47_3009 ();
 sg13g2_decap_8 FILLER_47_3016 ();
 sg13g2_decap_8 FILLER_47_3023 ();
 sg13g2_decap_8 FILLER_47_3030 ();
 sg13g2_decap_8 FILLER_47_3037 ();
 sg13g2_decap_8 FILLER_47_3044 ();
 sg13g2_decap_8 FILLER_47_3051 ();
 sg13g2_decap_8 FILLER_47_3058 ();
 sg13g2_decap_8 FILLER_47_3065 ();
 sg13g2_decap_8 FILLER_47_3072 ();
 sg13g2_decap_8 FILLER_47_3079 ();
 sg13g2_decap_8 FILLER_47_3086 ();
 sg13g2_decap_8 FILLER_47_3093 ();
 sg13g2_decap_8 FILLER_47_3100 ();
 sg13g2_decap_8 FILLER_47_3107 ();
 sg13g2_decap_8 FILLER_47_3114 ();
 sg13g2_decap_8 FILLER_47_3121 ();
 sg13g2_decap_8 FILLER_47_3128 ();
 sg13g2_decap_8 FILLER_47_3135 ();
 sg13g2_decap_8 FILLER_47_3142 ();
 sg13g2_decap_8 FILLER_47_3149 ();
 sg13g2_decap_8 FILLER_47_3156 ();
 sg13g2_decap_8 FILLER_47_3163 ();
 sg13g2_decap_8 FILLER_47_3170 ();
 sg13g2_decap_8 FILLER_47_3177 ();
 sg13g2_decap_8 FILLER_47_3184 ();
 sg13g2_decap_8 FILLER_47_3191 ();
 sg13g2_decap_8 FILLER_47_3198 ();
 sg13g2_decap_8 FILLER_47_3205 ();
 sg13g2_decap_8 FILLER_47_3212 ();
 sg13g2_decap_8 FILLER_47_3219 ();
 sg13g2_decap_8 FILLER_47_3226 ();
 sg13g2_decap_8 FILLER_47_3233 ();
 sg13g2_decap_8 FILLER_47_3240 ();
 sg13g2_decap_8 FILLER_47_3247 ();
 sg13g2_decap_8 FILLER_47_3254 ();
 sg13g2_decap_8 FILLER_47_3261 ();
 sg13g2_decap_8 FILLER_47_3268 ();
 sg13g2_decap_8 FILLER_47_3275 ();
 sg13g2_decap_8 FILLER_47_3282 ();
 sg13g2_decap_8 FILLER_47_3289 ();
 sg13g2_decap_8 FILLER_47_3296 ();
 sg13g2_decap_8 FILLER_47_3303 ();
 sg13g2_decap_8 FILLER_47_3310 ();
 sg13g2_decap_8 FILLER_47_3317 ();
 sg13g2_decap_8 FILLER_47_3324 ();
 sg13g2_decap_8 FILLER_47_3331 ();
 sg13g2_decap_8 FILLER_47_3338 ();
 sg13g2_decap_8 FILLER_47_3345 ();
 sg13g2_decap_8 FILLER_47_3352 ();
 sg13g2_decap_8 FILLER_47_3359 ();
 sg13g2_decap_8 FILLER_47_3366 ();
 sg13g2_decap_8 FILLER_47_3373 ();
 sg13g2_decap_8 FILLER_47_3380 ();
 sg13g2_decap_8 FILLER_47_3387 ();
 sg13g2_decap_8 FILLER_47_3394 ();
 sg13g2_decap_8 FILLER_47_3401 ();
 sg13g2_decap_8 FILLER_47_3408 ();
 sg13g2_decap_8 FILLER_47_3415 ();
 sg13g2_decap_8 FILLER_47_3422 ();
 sg13g2_decap_8 FILLER_47_3429 ();
 sg13g2_decap_8 FILLER_47_3436 ();
 sg13g2_decap_8 FILLER_47_3443 ();
 sg13g2_decap_8 FILLER_47_3450 ();
 sg13g2_decap_8 FILLER_47_3457 ();
 sg13g2_decap_8 FILLER_47_3464 ();
 sg13g2_decap_8 FILLER_47_3471 ();
 sg13g2_decap_8 FILLER_47_3478 ();
 sg13g2_decap_8 FILLER_47_3485 ();
 sg13g2_decap_8 FILLER_47_3492 ();
 sg13g2_decap_8 FILLER_47_3499 ();
 sg13g2_decap_8 FILLER_47_3506 ();
 sg13g2_decap_8 FILLER_47_3513 ();
 sg13g2_decap_8 FILLER_47_3520 ();
 sg13g2_decap_8 FILLER_47_3527 ();
 sg13g2_decap_8 FILLER_47_3534 ();
 sg13g2_decap_8 FILLER_47_3541 ();
 sg13g2_decap_8 FILLER_47_3548 ();
 sg13g2_decap_8 FILLER_47_3555 ();
 sg13g2_decap_8 FILLER_47_3562 ();
 sg13g2_decap_8 FILLER_47_3569 ();
 sg13g2_decap_4 FILLER_47_3576 ();
 sg13g2_fill_1 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_55 ();
 sg13g2_decap_4 FILLER_48_62 ();
 sg13g2_fill_2 FILLER_48_66 ();
 sg13g2_decap_8 FILLER_48_144 ();
 sg13g2_fill_1 FILLER_48_151 ();
 sg13g2_decap_8 FILLER_48_174 ();
 sg13g2_fill_1 FILLER_48_181 ();
 sg13g2_fill_1 FILLER_48_200 ();
 sg13g2_fill_2 FILLER_48_208 ();
 sg13g2_fill_1 FILLER_48_236 ();
 sg13g2_fill_2 FILLER_48_263 ();
 sg13g2_fill_1 FILLER_48_265 ();
 sg13g2_fill_2 FILLER_48_271 ();
 sg13g2_fill_1 FILLER_48_273 ();
 sg13g2_fill_2 FILLER_48_289 ();
 sg13g2_fill_1 FILLER_48_291 ();
 sg13g2_decap_4 FILLER_48_301 ();
 sg13g2_fill_2 FILLER_48_305 ();
 sg13g2_decap_4 FILLER_48_321 ();
 sg13g2_fill_2 FILLER_48_325 ();
 sg13g2_fill_2 FILLER_48_353 ();
 sg13g2_fill_2 FILLER_48_364 ();
 sg13g2_decap_8 FILLER_48_369 ();
 sg13g2_fill_1 FILLER_48_384 ();
 sg13g2_fill_2 FILLER_48_399 ();
 sg13g2_fill_1 FILLER_48_401 ();
 sg13g2_decap_4 FILLER_48_420 ();
 sg13g2_fill_2 FILLER_48_470 ();
 sg13g2_decap_8 FILLER_48_492 ();
 sg13g2_fill_2 FILLER_48_499 ();
 sg13g2_decap_8 FILLER_48_531 ();
 sg13g2_decap_8 FILLER_48_538 ();
 sg13g2_decap_8 FILLER_48_566 ();
 sg13g2_decap_8 FILLER_48_573 ();
 sg13g2_decap_4 FILLER_48_580 ();
 sg13g2_decap_8 FILLER_48_594 ();
 sg13g2_fill_1 FILLER_48_601 ();
 sg13g2_fill_1 FILLER_48_641 ();
 sg13g2_fill_1 FILLER_48_673 ();
 sg13g2_fill_1 FILLER_48_689 ();
 sg13g2_decap_8 FILLER_48_727 ();
 sg13g2_fill_2 FILLER_48_756 ();
 sg13g2_fill_1 FILLER_48_758 ();
 sg13g2_decap_8 FILLER_48_769 ();
 sg13g2_fill_2 FILLER_48_776 ();
 sg13g2_fill_1 FILLER_48_778 ();
 sg13g2_decap_8 FILLER_48_812 ();
 sg13g2_decap_8 FILLER_48_819 ();
 sg13g2_fill_1 FILLER_48_826 ();
 sg13g2_decap_8 FILLER_48_842 ();
 sg13g2_decap_8 FILLER_48_849 ();
 sg13g2_decap_4 FILLER_48_856 ();
 sg13g2_fill_1 FILLER_48_860 ();
 sg13g2_fill_2 FILLER_48_901 ();
 sg13g2_fill_1 FILLER_48_903 ();
 sg13g2_fill_1 FILLER_48_916 ();
 sg13g2_fill_2 FILLER_48_927 ();
 sg13g2_fill_1 FILLER_48_1013 ();
 sg13g2_fill_1 FILLER_48_1041 ();
 sg13g2_fill_2 FILLER_48_1093 ();
 sg13g2_decap_8 FILLER_48_1098 ();
 sg13g2_fill_2 FILLER_48_1105 ();
 sg13g2_fill_1 FILLER_48_1107 ();
 sg13g2_decap_8 FILLER_48_1115 ();
 sg13g2_decap_4 FILLER_48_1122 ();
 sg13g2_decap_4 FILLER_48_1152 ();
 sg13g2_fill_2 FILLER_48_1161 ();
 sg13g2_fill_1 FILLER_48_1163 ();
 sg13g2_decap_4 FILLER_48_1169 ();
 sg13g2_fill_2 FILLER_48_1177 ();
 sg13g2_decap_8 FILLER_48_1184 ();
 sg13g2_decap_8 FILLER_48_1191 ();
 sg13g2_decap_8 FILLER_48_1202 ();
 sg13g2_decap_8 FILLER_48_1209 ();
 sg13g2_decap_8 FILLER_48_1216 ();
 sg13g2_fill_2 FILLER_48_1223 ();
 sg13g2_fill_1 FILLER_48_1225 ();
 sg13g2_decap_8 FILLER_48_1231 ();
 sg13g2_fill_2 FILLER_48_1251 ();
 sg13g2_decap_4 FILLER_48_1261 ();
 sg13g2_fill_2 FILLER_48_1265 ();
 sg13g2_fill_1 FILLER_48_1306 ();
 sg13g2_fill_2 FILLER_48_1312 ();
 sg13g2_fill_1 FILLER_48_1314 ();
 sg13g2_fill_1 FILLER_48_1321 ();
 sg13g2_decap_4 FILLER_48_1348 ();
 sg13g2_fill_2 FILLER_48_1352 ();
 sg13g2_decap_8 FILLER_48_1357 ();
 sg13g2_decap_8 FILLER_48_1364 ();
 sg13g2_fill_2 FILLER_48_1371 ();
 sg13g2_fill_1 FILLER_48_1373 ();
 sg13g2_fill_2 FILLER_48_1413 ();
 sg13g2_fill_1 FILLER_48_1415 ();
 sg13g2_decap_8 FILLER_48_1435 ();
 sg13g2_decap_4 FILLER_48_1442 ();
 sg13g2_fill_1 FILLER_48_1476 ();
 sg13g2_fill_2 FILLER_48_1503 ();
 sg13g2_fill_1 FILLER_48_1505 ();
 sg13g2_decap_4 FILLER_48_1521 ();
 sg13g2_fill_2 FILLER_48_1537 ();
 sg13g2_fill_1 FILLER_48_1539 ();
 sg13g2_decap_4 FILLER_48_1548 ();
 sg13g2_fill_2 FILLER_48_1552 ();
 sg13g2_fill_1 FILLER_48_1562 ();
 sg13g2_fill_2 FILLER_48_1584 ();
 sg13g2_fill_1 FILLER_48_1586 ();
 sg13g2_decap_4 FILLER_48_1591 ();
 sg13g2_decap_4 FILLER_48_1600 ();
 sg13g2_fill_1 FILLER_48_1604 ();
 sg13g2_fill_1 FILLER_48_1609 ();
 sg13g2_decap_8 FILLER_48_1619 ();
 sg13g2_fill_2 FILLER_48_1645 ();
 sg13g2_fill_1 FILLER_48_1647 ();
 sg13g2_decap_4 FILLER_48_1654 ();
 sg13g2_fill_2 FILLER_48_1658 ();
 sg13g2_fill_2 FILLER_48_1677 ();
 sg13g2_fill_2 FILLER_48_1684 ();
 sg13g2_fill_1 FILLER_48_1686 ();
 sg13g2_decap_4 FILLER_48_1705 ();
 sg13g2_fill_2 FILLER_48_1736 ();
 sg13g2_fill_1 FILLER_48_1738 ();
 sg13g2_fill_2 FILLER_48_1744 ();
 sg13g2_fill_1 FILLER_48_1746 ();
 sg13g2_decap_4 FILLER_48_1772 ();
 sg13g2_fill_2 FILLER_48_1776 ();
 sg13g2_decap_8 FILLER_48_1789 ();
 sg13g2_decap_4 FILLER_48_1796 ();
 sg13g2_fill_1 FILLER_48_1800 ();
 sg13g2_decap_8 FILLER_48_1814 ();
 sg13g2_decap_4 FILLER_48_1821 ();
 sg13g2_fill_1 FILLER_48_1825 ();
 sg13g2_fill_2 FILLER_48_1852 ();
 sg13g2_fill_1 FILLER_48_1854 ();
 sg13g2_fill_1 FILLER_48_1873 ();
 sg13g2_fill_2 FILLER_48_1880 ();
 sg13g2_fill_1 FILLER_48_1882 ();
 sg13g2_fill_1 FILLER_48_1892 ();
 sg13g2_decap_8 FILLER_48_1902 ();
 sg13g2_decap_4 FILLER_48_1909 ();
 sg13g2_decap_8 FILLER_48_1946 ();
 sg13g2_decap_8 FILLER_48_1971 ();
 sg13g2_fill_1 FILLER_48_1992 ();
 sg13g2_decap_8 FILLER_48_2002 ();
 sg13g2_fill_2 FILLER_48_2009 ();
 sg13g2_decap_4 FILLER_48_2017 ();
 sg13g2_decap_8 FILLER_48_2045 ();
 sg13g2_fill_1 FILLER_48_2052 ();
 sg13g2_decap_8 FILLER_48_2071 ();
 sg13g2_decap_8 FILLER_48_2078 ();
 sg13g2_fill_1 FILLER_48_2085 ();
 sg13g2_fill_2 FILLER_48_2102 ();
 sg13g2_fill_1 FILLER_48_2104 ();
 sg13g2_fill_2 FILLER_48_2109 ();
 sg13g2_fill_1 FILLER_48_2111 ();
 sg13g2_decap_4 FILLER_48_2129 ();
 sg13g2_fill_2 FILLER_48_2141 ();
 sg13g2_decap_4 FILLER_48_2162 ();
 sg13g2_decap_8 FILLER_48_2180 ();
 sg13g2_decap_4 FILLER_48_2187 ();
 sg13g2_fill_2 FILLER_48_2191 ();
 sg13g2_decap_8 FILLER_48_2206 ();
 sg13g2_decap_8 FILLER_48_2221 ();
 sg13g2_fill_2 FILLER_48_2238 ();
 sg13g2_decap_4 FILLER_48_2255 ();
 sg13g2_decap_4 FILLER_48_2284 ();
 sg13g2_fill_1 FILLER_48_2288 ();
 sg13g2_fill_2 FILLER_48_2294 ();
 sg13g2_fill_1 FILLER_48_2296 ();
 sg13g2_decap_8 FILLER_48_2312 ();
 sg13g2_fill_2 FILLER_48_2319 ();
 sg13g2_fill_1 FILLER_48_2321 ();
 sg13g2_fill_2 FILLER_48_2335 ();
 sg13g2_fill_1 FILLER_48_2337 ();
 sg13g2_decap_8 FILLER_48_2342 ();
 sg13g2_fill_1 FILLER_48_2382 ();
 sg13g2_fill_1 FILLER_48_2395 ();
 sg13g2_fill_1 FILLER_48_2411 ();
 sg13g2_decap_4 FILLER_48_2447 ();
 sg13g2_decap_4 FILLER_48_2455 ();
 sg13g2_decap_8 FILLER_48_2474 ();
 sg13g2_decap_8 FILLER_48_2485 ();
 sg13g2_fill_1 FILLER_48_2492 ();
 sg13g2_fill_2 FILLER_48_2509 ();
 sg13g2_fill_1 FILLER_48_2511 ();
 sg13g2_fill_2 FILLER_48_2521 ();
 sg13g2_fill_1 FILLER_48_2523 ();
 sg13g2_decap_8 FILLER_48_2533 ();
 sg13g2_decap_8 FILLER_48_2544 ();
 sg13g2_fill_2 FILLER_48_2551 ();
 sg13g2_fill_1 FILLER_48_2553 ();
 sg13g2_decap_4 FILLER_48_2599 ();
 sg13g2_decap_4 FILLER_48_2606 ();
 sg13g2_fill_2 FILLER_48_2610 ();
 sg13g2_decap_8 FILLER_48_2625 ();
 sg13g2_decap_8 FILLER_48_2663 ();
 sg13g2_fill_2 FILLER_48_2670 ();
 sg13g2_fill_2 FILLER_48_2681 ();
 sg13g2_decap_8 FILLER_48_2693 ();
 sg13g2_decap_8 FILLER_48_2700 ();
 sg13g2_fill_2 FILLER_48_2707 ();
 sg13g2_fill_2 FILLER_48_2721 ();
 sg13g2_fill_1 FILLER_48_2723 ();
 sg13g2_fill_2 FILLER_48_2733 ();
 sg13g2_decap_8 FILLER_48_2758 ();
 sg13g2_decap_8 FILLER_48_2765 ();
 sg13g2_decap_4 FILLER_48_2776 ();
 sg13g2_fill_2 FILLER_48_2780 ();
 sg13g2_fill_2 FILLER_48_2804 ();
 sg13g2_fill_1 FILLER_48_2806 ();
 sg13g2_decap_8 FILLER_48_2821 ();
 sg13g2_decap_4 FILLER_48_2828 ();
 sg13g2_fill_1 FILLER_48_2844 ();
 sg13g2_decap_8 FILLER_48_2860 ();
 sg13g2_fill_1 FILLER_48_2883 ();
 sg13g2_fill_1 FILLER_48_2906 ();
 sg13g2_decap_8 FILLER_48_2965 ();
 sg13g2_decap_8 FILLER_48_2972 ();
 sg13g2_decap_8 FILLER_48_2979 ();
 sg13g2_decap_8 FILLER_48_2986 ();
 sg13g2_decap_8 FILLER_48_2993 ();
 sg13g2_decap_8 FILLER_48_3000 ();
 sg13g2_decap_8 FILLER_48_3007 ();
 sg13g2_decap_8 FILLER_48_3014 ();
 sg13g2_decap_8 FILLER_48_3021 ();
 sg13g2_decap_8 FILLER_48_3028 ();
 sg13g2_decap_8 FILLER_48_3035 ();
 sg13g2_decap_8 FILLER_48_3042 ();
 sg13g2_decap_8 FILLER_48_3049 ();
 sg13g2_decap_8 FILLER_48_3056 ();
 sg13g2_decap_8 FILLER_48_3063 ();
 sg13g2_decap_8 FILLER_48_3070 ();
 sg13g2_decap_8 FILLER_48_3077 ();
 sg13g2_decap_8 FILLER_48_3084 ();
 sg13g2_decap_8 FILLER_48_3091 ();
 sg13g2_decap_8 FILLER_48_3098 ();
 sg13g2_decap_8 FILLER_48_3105 ();
 sg13g2_decap_8 FILLER_48_3112 ();
 sg13g2_decap_8 FILLER_48_3119 ();
 sg13g2_decap_8 FILLER_48_3126 ();
 sg13g2_decap_8 FILLER_48_3133 ();
 sg13g2_decap_8 FILLER_48_3140 ();
 sg13g2_decap_8 FILLER_48_3147 ();
 sg13g2_decap_8 FILLER_48_3154 ();
 sg13g2_decap_8 FILLER_48_3161 ();
 sg13g2_decap_8 FILLER_48_3168 ();
 sg13g2_decap_8 FILLER_48_3175 ();
 sg13g2_decap_8 FILLER_48_3182 ();
 sg13g2_decap_8 FILLER_48_3189 ();
 sg13g2_decap_8 FILLER_48_3196 ();
 sg13g2_decap_8 FILLER_48_3203 ();
 sg13g2_decap_8 FILLER_48_3210 ();
 sg13g2_decap_8 FILLER_48_3217 ();
 sg13g2_decap_8 FILLER_48_3224 ();
 sg13g2_decap_8 FILLER_48_3231 ();
 sg13g2_decap_8 FILLER_48_3238 ();
 sg13g2_decap_8 FILLER_48_3245 ();
 sg13g2_decap_8 FILLER_48_3252 ();
 sg13g2_decap_8 FILLER_48_3259 ();
 sg13g2_decap_8 FILLER_48_3266 ();
 sg13g2_decap_8 FILLER_48_3273 ();
 sg13g2_decap_8 FILLER_48_3280 ();
 sg13g2_decap_8 FILLER_48_3287 ();
 sg13g2_decap_8 FILLER_48_3294 ();
 sg13g2_decap_8 FILLER_48_3301 ();
 sg13g2_decap_8 FILLER_48_3308 ();
 sg13g2_decap_8 FILLER_48_3315 ();
 sg13g2_decap_8 FILLER_48_3322 ();
 sg13g2_decap_8 FILLER_48_3329 ();
 sg13g2_decap_8 FILLER_48_3336 ();
 sg13g2_decap_8 FILLER_48_3343 ();
 sg13g2_decap_8 FILLER_48_3350 ();
 sg13g2_decap_8 FILLER_48_3357 ();
 sg13g2_decap_8 FILLER_48_3364 ();
 sg13g2_decap_8 FILLER_48_3371 ();
 sg13g2_decap_8 FILLER_48_3378 ();
 sg13g2_decap_8 FILLER_48_3385 ();
 sg13g2_decap_8 FILLER_48_3392 ();
 sg13g2_decap_8 FILLER_48_3399 ();
 sg13g2_decap_8 FILLER_48_3406 ();
 sg13g2_decap_8 FILLER_48_3413 ();
 sg13g2_decap_8 FILLER_48_3420 ();
 sg13g2_decap_8 FILLER_48_3427 ();
 sg13g2_decap_8 FILLER_48_3434 ();
 sg13g2_decap_8 FILLER_48_3441 ();
 sg13g2_decap_8 FILLER_48_3448 ();
 sg13g2_decap_8 FILLER_48_3455 ();
 sg13g2_decap_8 FILLER_48_3462 ();
 sg13g2_decap_8 FILLER_48_3469 ();
 sg13g2_decap_8 FILLER_48_3476 ();
 sg13g2_decap_8 FILLER_48_3483 ();
 sg13g2_decap_8 FILLER_48_3490 ();
 sg13g2_decap_8 FILLER_48_3497 ();
 sg13g2_decap_8 FILLER_48_3504 ();
 sg13g2_decap_8 FILLER_48_3511 ();
 sg13g2_decap_8 FILLER_48_3518 ();
 sg13g2_decap_8 FILLER_48_3525 ();
 sg13g2_decap_8 FILLER_48_3532 ();
 sg13g2_decap_8 FILLER_48_3539 ();
 sg13g2_decap_8 FILLER_48_3546 ();
 sg13g2_decap_8 FILLER_48_3553 ();
 sg13g2_decap_8 FILLER_48_3560 ();
 sg13g2_decap_8 FILLER_48_3567 ();
 sg13g2_decap_4 FILLER_48_3574 ();
 sg13g2_fill_2 FILLER_48_3578 ();
 sg13g2_fill_2 FILLER_49_0 ();
 sg13g2_fill_1 FILLER_49_28 ();
 sg13g2_fill_2 FILLER_49_44 ();
 sg13g2_fill_1 FILLER_49_46 ();
 sg13g2_fill_2 FILLER_49_59 ();
 sg13g2_fill_1 FILLER_49_61 ();
 sg13g2_decap_4 FILLER_49_92 ();
 sg13g2_fill_2 FILLER_49_96 ();
 sg13g2_fill_2 FILLER_49_152 ();
 sg13g2_fill_1 FILLER_49_154 ();
 sg13g2_fill_2 FILLER_49_160 ();
 sg13g2_fill_1 FILLER_49_162 ();
 sg13g2_fill_2 FILLER_49_189 ();
 sg13g2_fill_1 FILLER_49_191 ();
 sg13g2_fill_2 FILLER_49_220 ();
 sg13g2_fill_1 FILLER_49_222 ();
 sg13g2_fill_2 FILLER_49_232 ();
 sg13g2_fill_2 FILLER_49_266 ();
 sg13g2_fill_2 FILLER_49_273 ();
 sg13g2_decap_4 FILLER_49_280 ();
 sg13g2_fill_1 FILLER_49_284 ();
 sg13g2_fill_2 FILLER_49_329 ();
 sg13g2_fill_1 FILLER_49_331 ();
 sg13g2_fill_1 FILLER_49_337 ();
 sg13g2_fill_2 FILLER_49_342 ();
 sg13g2_fill_2 FILLER_49_379 ();
 sg13g2_fill_1 FILLER_49_415 ();
 sg13g2_fill_1 FILLER_49_425 ();
 sg13g2_fill_1 FILLER_49_430 ();
 sg13g2_fill_2 FILLER_49_471 ();
 sg13g2_fill_1 FILLER_49_473 ();
 sg13g2_fill_2 FILLER_49_479 ();
 sg13g2_fill_1 FILLER_49_481 ();
 sg13g2_decap_8 FILLER_49_487 ();
 sg13g2_fill_2 FILLER_49_509 ();
 sg13g2_fill_1 FILLER_49_511 ();
 sg13g2_decap_8 FILLER_49_520 ();
 sg13g2_decap_4 FILLER_49_527 ();
 sg13g2_fill_2 FILLER_49_531 ();
 sg13g2_decap_4 FILLER_49_545 ();
 sg13g2_fill_2 FILLER_49_623 ();
 sg13g2_decap_8 FILLER_49_629 ();
 sg13g2_decap_8 FILLER_49_636 ();
 sg13g2_fill_2 FILLER_49_643 ();
 sg13g2_fill_1 FILLER_49_645 ();
 sg13g2_fill_2 FILLER_49_669 ();
 sg13g2_fill_2 FILLER_49_711 ();
 sg13g2_fill_1 FILLER_49_713 ();
 sg13g2_fill_2 FILLER_49_720 ();
 sg13g2_decap_4 FILLER_49_727 ();
 sg13g2_fill_1 FILLER_49_736 ();
 sg13g2_fill_1 FILLER_49_742 ();
 sg13g2_decap_4 FILLER_49_769 ();
 sg13g2_fill_2 FILLER_49_773 ();
 sg13g2_fill_2 FILLER_49_780 ();
 sg13g2_fill_1 FILLER_49_787 ();
 sg13g2_decap_4 FILLER_49_806 ();
 sg13g2_decap_8 FILLER_49_814 ();
 sg13g2_fill_1 FILLER_49_821 ();
 sg13g2_fill_2 FILLER_49_835 ();
 sg13g2_decap_8 FILLER_49_842 ();
 sg13g2_fill_2 FILLER_49_855 ();
 sg13g2_fill_1 FILLER_49_857 ();
 sg13g2_decap_8 FILLER_49_874 ();
 sg13g2_decap_4 FILLER_49_881 ();
 sg13g2_fill_1 FILLER_49_885 ();
 sg13g2_fill_2 FILLER_49_891 ();
 sg13g2_decap_8 FILLER_49_898 ();
 sg13g2_fill_1 FILLER_49_938 ();
 sg13g2_fill_1 FILLER_49_958 ();
 sg13g2_fill_1 FILLER_49_968 ();
 sg13g2_fill_2 FILLER_49_999 ();
 sg13g2_decap_8 FILLER_49_1006 ();
 sg13g2_fill_1 FILLER_49_1013 ();
 sg13g2_fill_2 FILLER_49_1018 ();
 sg13g2_fill_1 FILLER_49_1020 ();
 sg13g2_fill_1 FILLER_49_1030 ();
 sg13g2_fill_2 FILLER_49_1062 ();
 sg13g2_decap_4 FILLER_49_1074 ();
 sg13g2_decap_4 FILLER_49_1091 ();
 sg13g2_fill_1 FILLER_49_1154 ();
 sg13g2_fill_1 FILLER_49_1241 ();
 sg13g2_fill_1 FILLER_49_1251 ();
 sg13g2_fill_2 FILLER_49_1257 ();
 sg13g2_fill_1 FILLER_49_1259 ();
 sg13g2_fill_2 FILLER_49_1274 ();
 sg13g2_fill_1 FILLER_49_1276 ();
 sg13g2_fill_1 FILLER_49_1324 ();
 sg13g2_fill_2 FILLER_49_1343 ();
 sg13g2_fill_1 FILLER_49_1345 ();
 sg13g2_decap_8 FILLER_49_1360 ();
 sg13g2_fill_2 FILLER_49_1367 ();
 sg13g2_decap_8 FILLER_49_1373 ();
 sg13g2_decap_8 FILLER_49_1380 ();
 sg13g2_decap_8 FILLER_49_1387 ();
 sg13g2_fill_2 FILLER_49_1394 ();
 sg13g2_decap_8 FILLER_49_1406 ();
 sg13g2_decap_8 FILLER_49_1413 ();
 sg13g2_fill_2 FILLER_49_1420 ();
 sg13g2_fill_1 FILLER_49_1422 ();
 sg13g2_decap_4 FILLER_49_1453 ();
 sg13g2_decap_8 FILLER_49_1462 ();
 sg13g2_fill_1 FILLER_49_1469 ();
 sg13g2_decap_4 FILLER_49_1483 ();
 sg13g2_fill_1 FILLER_49_1520 ();
 sg13g2_decap_8 FILLER_49_1541 ();
 sg13g2_decap_4 FILLER_49_1566 ();
 sg13g2_fill_2 FILLER_49_1570 ();
 sg13g2_fill_1 FILLER_49_1607 ();
 sg13g2_decap_4 FILLER_49_1613 ();
 sg13g2_fill_2 FILLER_49_1628 ();
 sg13g2_fill_2 FILLER_49_1649 ();
 sg13g2_fill_1 FILLER_49_1651 ();
 sg13g2_fill_2 FILLER_49_1656 ();
 sg13g2_fill_1 FILLER_49_1658 ();
 sg13g2_fill_1 FILLER_49_1664 ();
 sg13g2_decap_4 FILLER_49_1673 ();
 sg13g2_fill_2 FILLER_49_1677 ();
 sg13g2_fill_1 FILLER_49_1689 ();
 sg13g2_decap_8 FILLER_49_1708 ();
 sg13g2_decap_4 FILLER_49_1715 ();
 sg13g2_decap_8 FILLER_49_1747 ();
 sg13g2_fill_1 FILLER_49_1754 ();
 sg13g2_decap_4 FILLER_49_1794 ();
 sg13g2_decap_4 FILLER_49_1805 ();
 sg13g2_fill_1 FILLER_49_1809 ();
 sg13g2_decap_4 FILLER_49_1813 ();
 sg13g2_decap_8 FILLER_49_1835 ();
 sg13g2_decap_8 FILLER_49_1859 ();
 sg13g2_fill_1 FILLER_49_1901 ();
 sg13g2_decap_8 FILLER_49_1915 ();
 sg13g2_decap_8 FILLER_49_1922 ();
 sg13g2_fill_1 FILLER_49_1929 ();
 sg13g2_decap_8 FILLER_49_1934 ();
 sg13g2_decap_8 FILLER_49_1941 ();
 sg13g2_decap_4 FILLER_49_1948 ();
 sg13g2_fill_1 FILLER_49_1952 ();
 sg13g2_decap_8 FILLER_49_1970 ();
 sg13g2_fill_1 FILLER_49_1977 ();
 sg13g2_decap_4 FILLER_49_1995 ();
 sg13g2_fill_2 FILLER_49_2017 ();
 sg13g2_decap_4 FILLER_49_2032 ();
 sg13g2_fill_2 FILLER_49_2036 ();
 sg13g2_fill_2 FILLER_49_2043 ();
 sg13g2_fill_1 FILLER_49_2045 ();
 sg13g2_decap_4 FILLER_49_2050 ();
 sg13g2_fill_1 FILLER_49_2054 ();
 sg13g2_fill_1 FILLER_49_2059 ();
 sg13g2_decap_4 FILLER_49_2076 ();
 sg13g2_fill_2 FILLER_49_2080 ();
 sg13g2_decap_8 FILLER_49_2096 ();
 sg13g2_fill_2 FILLER_49_2121 ();
 sg13g2_fill_1 FILLER_49_2123 ();
 sg13g2_decap_8 FILLER_49_2132 ();
 sg13g2_fill_1 FILLER_49_2139 ();
 sg13g2_fill_2 FILLER_49_2155 ();
 sg13g2_fill_1 FILLER_49_2157 ();
 sg13g2_fill_2 FILLER_49_2187 ();
 sg13g2_fill_2 FILLER_49_2205 ();
 sg13g2_fill_1 FILLER_49_2207 ();
 sg13g2_decap_8 FILLER_49_2233 ();
 sg13g2_decap_4 FILLER_49_2240 ();
 sg13g2_fill_1 FILLER_49_2244 ();
 sg13g2_decap_4 FILLER_49_2249 ();
 sg13g2_fill_1 FILLER_49_2253 ();
 sg13g2_fill_2 FILLER_49_2269 ();
 sg13g2_fill_1 FILLER_49_2271 ();
 sg13g2_decap_8 FILLER_49_2280 ();
 sg13g2_decap_8 FILLER_49_2287 ();
 sg13g2_fill_2 FILLER_49_2294 ();
 sg13g2_decap_4 FILLER_49_2305 ();
 sg13g2_fill_2 FILLER_49_2309 ();
 sg13g2_fill_2 FILLER_49_2316 ();
 sg13g2_fill_1 FILLER_49_2318 ();
 sg13g2_fill_2 FILLER_49_2330 ();
 sg13g2_fill_1 FILLER_49_2332 ();
 sg13g2_decap_4 FILLER_49_2352 ();
 sg13g2_fill_2 FILLER_49_2356 ();
 sg13g2_decap_4 FILLER_49_2363 ();
 sg13g2_fill_1 FILLER_49_2367 ();
 sg13g2_decap_8 FILLER_49_2380 ();
 sg13g2_decap_8 FILLER_49_2387 ();
 sg13g2_fill_2 FILLER_49_2394 ();
 sg13g2_decap_4 FILLER_49_2406 ();
 sg13g2_fill_1 FILLER_49_2410 ();
 sg13g2_decap_4 FILLER_49_2416 ();
 sg13g2_fill_2 FILLER_49_2420 ();
 sg13g2_decap_8 FILLER_49_2432 ();
 sg13g2_decap_8 FILLER_49_2439 ();
 sg13g2_fill_2 FILLER_49_2454 ();
 sg13g2_fill_1 FILLER_49_2456 ();
 sg13g2_decap_8 FILLER_49_2471 ();
 sg13g2_decap_8 FILLER_49_2478 ();
 sg13g2_decap_4 FILLER_49_2565 ();
 sg13g2_fill_1 FILLER_49_2598 ();
 sg13g2_fill_2 FILLER_49_2617 ();
 sg13g2_decap_8 FILLER_49_2631 ();
 sg13g2_decap_4 FILLER_49_2638 ();
 sg13g2_fill_2 FILLER_49_2642 ();
 sg13g2_decap_8 FILLER_49_2659 ();
 sg13g2_decap_8 FILLER_49_2666 ();
 sg13g2_fill_2 FILLER_49_2673 ();
 sg13g2_decap_4 FILLER_49_2699 ();
 sg13g2_fill_1 FILLER_49_2703 ();
 sg13g2_decap_8 FILLER_49_2764 ();
 sg13g2_fill_2 FILLER_49_2771 ();
 sg13g2_decap_8 FILLER_49_2777 ();
 sg13g2_fill_1 FILLER_49_2784 ();
 sg13g2_fill_1 FILLER_49_2807 ();
 sg13g2_fill_2 FILLER_49_2838 ();
 sg13g2_fill_2 FILLER_49_2859 ();
 sg13g2_decap_8 FILLER_49_2877 ();
 sg13g2_fill_2 FILLER_49_2884 ();
 sg13g2_fill_1 FILLER_49_2886 ();
 sg13g2_fill_2 FILLER_49_2891 ();
 sg13g2_fill_1 FILLER_49_2893 ();
 sg13g2_fill_1 FILLER_49_2910 ();
 sg13g2_fill_1 FILLER_49_2916 ();
 sg13g2_decap_8 FILLER_49_2921 ();
 sg13g2_decap_8 FILLER_49_2928 ();
 sg13g2_decap_8 FILLER_49_2935 ();
 sg13g2_decap_8 FILLER_49_2955 ();
 sg13g2_decap_8 FILLER_49_2962 ();
 sg13g2_decap_8 FILLER_49_2969 ();
 sg13g2_decap_8 FILLER_49_2976 ();
 sg13g2_decap_8 FILLER_49_2983 ();
 sg13g2_decap_8 FILLER_49_2990 ();
 sg13g2_decap_8 FILLER_49_2997 ();
 sg13g2_decap_8 FILLER_49_3004 ();
 sg13g2_decap_8 FILLER_49_3011 ();
 sg13g2_decap_8 FILLER_49_3018 ();
 sg13g2_decap_8 FILLER_49_3025 ();
 sg13g2_decap_8 FILLER_49_3032 ();
 sg13g2_decap_8 FILLER_49_3039 ();
 sg13g2_decap_8 FILLER_49_3046 ();
 sg13g2_decap_8 FILLER_49_3053 ();
 sg13g2_decap_8 FILLER_49_3060 ();
 sg13g2_decap_8 FILLER_49_3067 ();
 sg13g2_decap_8 FILLER_49_3074 ();
 sg13g2_decap_8 FILLER_49_3081 ();
 sg13g2_decap_8 FILLER_49_3088 ();
 sg13g2_decap_8 FILLER_49_3095 ();
 sg13g2_decap_8 FILLER_49_3102 ();
 sg13g2_decap_8 FILLER_49_3109 ();
 sg13g2_decap_8 FILLER_49_3116 ();
 sg13g2_decap_8 FILLER_49_3123 ();
 sg13g2_decap_8 FILLER_49_3130 ();
 sg13g2_decap_8 FILLER_49_3137 ();
 sg13g2_decap_8 FILLER_49_3144 ();
 sg13g2_decap_8 FILLER_49_3151 ();
 sg13g2_decap_8 FILLER_49_3158 ();
 sg13g2_decap_8 FILLER_49_3165 ();
 sg13g2_decap_8 FILLER_49_3172 ();
 sg13g2_decap_8 FILLER_49_3179 ();
 sg13g2_decap_8 FILLER_49_3186 ();
 sg13g2_decap_8 FILLER_49_3193 ();
 sg13g2_decap_8 FILLER_49_3200 ();
 sg13g2_decap_8 FILLER_49_3207 ();
 sg13g2_decap_8 FILLER_49_3214 ();
 sg13g2_decap_8 FILLER_49_3221 ();
 sg13g2_decap_8 FILLER_49_3228 ();
 sg13g2_decap_8 FILLER_49_3235 ();
 sg13g2_decap_8 FILLER_49_3242 ();
 sg13g2_decap_8 FILLER_49_3249 ();
 sg13g2_decap_8 FILLER_49_3256 ();
 sg13g2_decap_8 FILLER_49_3263 ();
 sg13g2_decap_8 FILLER_49_3270 ();
 sg13g2_decap_8 FILLER_49_3277 ();
 sg13g2_decap_8 FILLER_49_3284 ();
 sg13g2_decap_8 FILLER_49_3291 ();
 sg13g2_decap_8 FILLER_49_3298 ();
 sg13g2_decap_8 FILLER_49_3305 ();
 sg13g2_decap_8 FILLER_49_3312 ();
 sg13g2_decap_8 FILLER_49_3319 ();
 sg13g2_decap_8 FILLER_49_3326 ();
 sg13g2_decap_8 FILLER_49_3333 ();
 sg13g2_decap_8 FILLER_49_3340 ();
 sg13g2_decap_8 FILLER_49_3347 ();
 sg13g2_decap_8 FILLER_49_3354 ();
 sg13g2_decap_8 FILLER_49_3361 ();
 sg13g2_decap_8 FILLER_49_3368 ();
 sg13g2_decap_8 FILLER_49_3375 ();
 sg13g2_decap_8 FILLER_49_3382 ();
 sg13g2_decap_8 FILLER_49_3389 ();
 sg13g2_decap_8 FILLER_49_3396 ();
 sg13g2_decap_8 FILLER_49_3403 ();
 sg13g2_decap_8 FILLER_49_3410 ();
 sg13g2_decap_8 FILLER_49_3417 ();
 sg13g2_decap_8 FILLER_49_3424 ();
 sg13g2_decap_8 FILLER_49_3431 ();
 sg13g2_decap_8 FILLER_49_3438 ();
 sg13g2_decap_8 FILLER_49_3445 ();
 sg13g2_decap_8 FILLER_49_3452 ();
 sg13g2_decap_8 FILLER_49_3459 ();
 sg13g2_decap_8 FILLER_49_3466 ();
 sg13g2_decap_8 FILLER_49_3473 ();
 sg13g2_decap_8 FILLER_49_3480 ();
 sg13g2_decap_8 FILLER_49_3487 ();
 sg13g2_decap_8 FILLER_49_3494 ();
 sg13g2_decap_8 FILLER_49_3501 ();
 sg13g2_decap_8 FILLER_49_3508 ();
 sg13g2_decap_8 FILLER_49_3515 ();
 sg13g2_decap_8 FILLER_49_3522 ();
 sg13g2_decap_8 FILLER_49_3529 ();
 sg13g2_decap_8 FILLER_49_3536 ();
 sg13g2_decap_8 FILLER_49_3543 ();
 sg13g2_decap_8 FILLER_49_3550 ();
 sg13g2_decap_8 FILLER_49_3557 ();
 sg13g2_decap_8 FILLER_49_3564 ();
 sg13g2_decap_8 FILLER_49_3571 ();
 sg13g2_fill_2 FILLER_49_3578 ();
 sg13g2_fill_2 FILLER_50_26 ();
 sg13g2_fill_1 FILLER_50_43 ();
 sg13g2_fill_2 FILLER_50_55 ();
 sg13g2_fill_2 FILLER_50_87 ();
 sg13g2_fill_1 FILLER_50_89 ();
 sg13g2_decap_4 FILLER_50_95 ();
 sg13g2_fill_1 FILLER_50_121 ();
 sg13g2_decap_8 FILLER_50_162 ();
 sg13g2_decap_4 FILLER_50_169 ();
 sg13g2_fill_1 FILLER_50_173 ();
 sg13g2_fill_1 FILLER_50_206 ();
 sg13g2_fill_2 FILLER_50_225 ();
 sg13g2_decap_8 FILLER_50_261 ();
 sg13g2_decap_8 FILLER_50_268 ();
 sg13g2_decap_8 FILLER_50_275 ();
 sg13g2_fill_1 FILLER_50_282 ();
 sg13g2_decap_8 FILLER_50_296 ();
 sg13g2_decap_4 FILLER_50_303 ();
 sg13g2_decap_4 FILLER_50_310 ();
 sg13g2_fill_1 FILLER_50_314 ();
 sg13g2_decap_4 FILLER_50_330 ();
 sg13g2_decap_8 FILLER_50_339 ();
 sg13g2_fill_2 FILLER_50_346 ();
 sg13g2_decap_8 FILLER_50_377 ();
 sg13g2_decap_8 FILLER_50_384 ();
 sg13g2_fill_2 FILLER_50_404 ();
 sg13g2_decap_8 FILLER_50_416 ();
 sg13g2_decap_8 FILLER_50_423 ();
 sg13g2_decap_4 FILLER_50_430 ();
 sg13g2_fill_2 FILLER_50_434 ();
 sg13g2_fill_2 FILLER_50_468 ();
 sg13g2_decap_4 FILLER_50_475 ();
 sg13g2_fill_1 FILLER_50_479 ();
 sg13g2_decap_4 FILLER_50_488 ();
 sg13g2_fill_1 FILLER_50_492 ();
 sg13g2_fill_1 FILLER_50_499 ();
 sg13g2_fill_2 FILLER_50_514 ();
 sg13g2_fill_1 FILLER_50_516 ();
 sg13g2_fill_2 FILLER_50_543 ();
 sg13g2_fill_1 FILLER_50_545 ();
 sg13g2_fill_1 FILLER_50_561 ();
 sg13g2_fill_1 FILLER_50_590 ();
 sg13g2_decap_4 FILLER_50_596 ();
 sg13g2_decap_8 FILLER_50_605 ();
 sg13g2_decap_8 FILLER_50_612 ();
 sg13g2_decap_8 FILLER_50_619 ();
 sg13g2_decap_4 FILLER_50_631 ();
 sg13g2_fill_1 FILLER_50_656 ();
 sg13g2_fill_2 FILLER_50_666 ();
 sg13g2_fill_2 FILLER_50_672 ();
 sg13g2_fill_1 FILLER_50_674 ();
 sg13g2_fill_2 FILLER_50_680 ();
 sg13g2_fill_1 FILLER_50_694 ();
 sg13g2_fill_2 FILLER_50_709 ();
 sg13g2_fill_1 FILLER_50_711 ();
 sg13g2_decap_8 FILLER_50_726 ();
 sg13g2_fill_2 FILLER_50_733 ();
 sg13g2_fill_1 FILLER_50_735 ();
 sg13g2_fill_2 FILLER_50_769 ();
 sg13g2_fill_1 FILLER_50_771 ();
 sg13g2_fill_2 FILLER_50_782 ();
 sg13g2_fill_1 FILLER_50_784 ();
 sg13g2_decap_4 FILLER_50_834 ();
 sg13g2_decap_8 FILLER_50_867 ();
 sg13g2_decap_4 FILLER_50_874 ();
 sg13g2_fill_2 FILLER_50_904 ();
 sg13g2_fill_1 FILLER_50_906 ();
 sg13g2_fill_2 FILLER_50_925 ();
 sg13g2_fill_1 FILLER_50_927 ();
 sg13g2_fill_2 FILLER_50_954 ();
 sg13g2_fill_1 FILLER_50_956 ();
 sg13g2_fill_2 FILLER_50_996 ();
 sg13g2_fill_1 FILLER_50_998 ();
 sg13g2_fill_1 FILLER_50_1007 ();
 sg13g2_decap_4 FILLER_50_1012 ();
 sg13g2_fill_1 FILLER_50_1059 ();
 sg13g2_decap_8 FILLER_50_1069 ();
 sg13g2_fill_1 FILLER_50_1076 ();
 sg13g2_decap_4 FILLER_50_1081 ();
 sg13g2_fill_1 FILLER_50_1085 ();
 sg13g2_decap_8 FILLER_50_1123 ();
 sg13g2_decap_8 FILLER_50_1130 ();
 sg13g2_fill_2 FILLER_50_1137 ();
 sg13g2_decap_8 FILLER_50_1154 ();
 sg13g2_decap_8 FILLER_50_1161 ();
 sg13g2_fill_2 FILLER_50_1168 ();
 sg13g2_decap_8 FILLER_50_1174 ();
 sg13g2_decap_4 FILLER_50_1181 ();
 sg13g2_fill_2 FILLER_50_1185 ();
 sg13g2_fill_2 FILLER_50_1193 ();
 sg13g2_decap_8 FILLER_50_1208 ();
 sg13g2_fill_2 FILLER_50_1215 ();
 sg13g2_fill_1 FILLER_50_1217 ();
 sg13g2_decap_4 FILLER_50_1222 ();
 sg13g2_fill_2 FILLER_50_1226 ();
 sg13g2_decap_4 FILLER_50_1283 ();
 sg13g2_fill_1 FILLER_50_1287 ();
 sg13g2_decap_8 FILLER_50_1292 ();
 sg13g2_decap_4 FILLER_50_1299 ();
 sg13g2_fill_1 FILLER_50_1303 ();
 sg13g2_decap_4 FILLER_50_1312 ();
 sg13g2_fill_1 FILLER_50_1346 ();
 sg13g2_decap_4 FILLER_50_1359 ();
 sg13g2_fill_2 FILLER_50_1363 ();
 sg13g2_fill_2 FILLER_50_1391 ();
 sg13g2_fill_1 FILLER_50_1393 ();
 sg13g2_decap_8 FILLER_50_1415 ();
 sg13g2_decap_4 FILLER_50_1422 ();
 sg13g2_fill_2 FILLER_50_1426 ();
 sg13g2_fill_1 FILLER_50_1436 ();
 sg13g2_fill_2 FILLER_50_1446 ();
 sg13g2_fill_2 FILLER_50_1458 ();
 sg13g2_fill_1 FILLER_50_1460 ();
 sg13g2_decap_8 FILLER_50_1492 ();
 sg13g2_fill_2 FILLER_50_1499 ();
 sg13g2_decap_8 FILLER_50_1506 ();
 sg13g2_decap_8 FILLER_50_1513 ();
 sg13g2_decap_8 FILLER_50_1520 ();
 sg13g2_fill_2 FILLER_50_1527 ();
 sg13g2_fill_1 FILLER_50_1529 ();
 sg13g2_decap_4 FILLER_50_1543 ();
 sg13g2_decap_8 FILLER_50_1573 ();
 sg13g2_decap_4 FILLER_50_1580 ();
 sg13g2_fill_2 FILLER_50_1584 ();
 sg13g2_fill_2 FILLER_50_1590 ();
 sg13g2_fill_2 FILLER_50_1597 ();
 sg13g2_decap_4 FILLER_50_1613 ();
 sg13g2_fill_2 FILLER_50_1622 ();
 sg13g2_fill_1 FILLER_50_1624 ();
 sg13g2_fill_1 FILLER_50_1636 ();
 sg13g2_fill_1 FILLER_50_1660 ();
 sg13g2_decap_8 FILLER_50_1678 ();
 sg13g2_decap_8 FILLER_50_1685 ();
 sg13g2_decap_8 FILLER_50_1692 ();
 sg13g2_fill_1 FILLER_50_1704 ();
 sg13g2_decap_8 FILLER_50_1711 ();
 sg13g2_fill_1 FILLER_50_1731 ();
 sg13g2_decap_4 FILLER_50_1743 ();
 sg13g2_fill_1 FILLER_50_1760 ();
 sg13g2_fill_2 FILLER_50_1770 ();
 sg13g2_decap_8 FILLER_50_1780 ();
 sg13g2_decap_4 FILLER_50_1792 ();
 sg13g2_fill_1 FILLER_50_1796 ();
 sg13g2_fill_2 FILLER_50_1810 ();
 sg13g2_decap_8 FILLER_50_1832 ();
 sg13g2_decap_8 FILLER_50_1839 ();
 sg13g2_decap_4 FILLER_50_1846 ();
 sg13g2_fill_1 FILLER_50_1850 ();
 sg13g2_decap_4 FILLER_50_1865 ();
 sg13g2_fill_1 FILLER_50_1869 ();
 sg13g2_decap_8 FILLER_50_1880 ();
 sg13g2_decap_8 FILLER_50_1906 ();
 sg13g2_fill_1 FILLER_50_1913 ();
 sg13g2_fill_2 FILLER_50_1918 ();
 sg13g2_fill_1 FILLER_50_1920 ();
 sg13g2_fill_1 FILLER_50_1941 ();
 sg13g2_decap_8 FILLER_50_1974 ();
 sg13g2_decap_8 FILLER_50_1981 ();
 sg13g2_fill_2 FILLER_50_1988 ();
 sg13g2_decap_8 FILLER_50_1996 ();
 sg13g2_decap_8 FILLER_50_2003 ();
 sg13g2_fill_1 FILLER_50_2010 ();
 sg13g2_fill_1 FILLER_50_2027 ();
 sg13g2_decap_8 FILLER_50_2048 ();
 sg13g2_decap_8 FILLER_50_2055 ();
 sg13g2_fill_2 FILLER_50_2062 ();
 sg13g2_fill_1 FILLER_50_2064 ();
 sg13g2_decap_8 FILLER_50_2076 ();
 sg13g2_decap_8 FILLER_50_2100 ();
 sg13g2_decap_8 FILLER_50_2107 ();
 sg13g2_decap_8 FILLER_50_2114 ();
 sg13g2_fill_2 FILLER_50_2121 ();
 sg13g2_decap_8 FILLER_50_2138 ();
 sg13g2_decap_4 FILLER_50_2145 ();
 sg13g2_fill_2 FILLER_50_2162 ();
 sg13g2_fill_1 FILLER_50_2164 ();
 sg13g2_decap_8 FILLER_50_2175 ();
 sg13g2_decap_8 FILLER_50_2187 ();
 sg13g2_decap_8 FILLER_50_2194 ();
 sg13g2_fill_2 FILLER_50_2206 ();
 sg13g2_decap_8 FILLER_50_2214 ();
 sg13g2_fill_2 FILLER_50_2221 ();
 sg13g2_fill_2 FILLER_50_2227 ();
 sg13g2_decap_8 FILLER_50_2237 ();
 sg13g2_fill_2 FILLER_50_2244 ();
 sg13g2_fill_1 FILLER_50_2246 ();
 sg13g2_decap_4 FILLER_50_2268 ();
 sg13g2_fill_2 FILLER_50_2276 ();
 sg13g2_fill_1 FILLER_50_2278 ();
 sg13g2_decap_8 FILLER_50_2284 ();
 sg13g2_fill_2 FILLER_50_2291 ();
 sg13g2_fill_1 FILLER_50_2293 ();
 sg13g2_decap_4 FILLER_50_2307 ();
 sg13g2_decap_4 FILLER_50_2315 ();
 sg13g2_fill_2 FILLER_50_2319 ();
 sg13g2_fill_1 FILLER_50_2362 ();
 sg13g2_fill_2 FILLER_50_2410 ();
 sg13g2_fill_1 FILLER_50_2412 ();
 sg13g2_fill_2 FILLER_50_2444 ();
 sg13g2_decap_4 FILLER_50_2465 ();
 sg13g2_fill_2 FILLER_50_2469 ();
 sg13g2_decap_8 FILLER_50_2499 ();
 sg13g2_fill_1 FILLER_50_2506 ();
 sg13g2_decap_8 FILLER_50_2530 ();
 sg13g2_decap_4 FILLER_50_2537 ();
 sg13g2_fill_1 FILLER_50_2541 ();
 sg13g2_decap_4 FILLER_50_2548 ();
 sg13g2_fill_2 FILLER_50_2552 ();
 sg13g2_fill_1 FILLER_50_2562 ();
 sg13g2_fill_1 FILLER_50_2568 ();
 sg13g2_decap_8 FILLER_50_2589 ();
 sg13g2_fill_2 FILLER_50_2614 ();
 sg13g2_fill_1 FILLER_50_2616 ();
 sg13g2_decap_4 FILLER_50_2630 ();
 sg13g2_fill_1 FILLER_50_2634 ();
 sg13g2_decap_8 FILLER_50_2640 ();
 sg13g2_fill_1 FILLER_50_2647 ();
 sg13g2_fill_1 FILLER_50_2670 ();
 sg13g2_decap_4 FILLER_50_2698 ();
 sg13g2_fill_1 FILLER_50_2702 ();
 sg13g2_fill_1 FILLER_50_2718 ();
 sg13g2_fill_2 FILLER_50_2728 ();
 sg13g2_fill_1 FILLER_50_2730 ();
 sg13g2_decap_8 FILLER_50_2742 ();
 sg13g2_decap_8 FILLER_50_2753 ();
 sg13g2_fill_2 FILLER_50_2760 ();
 sg13g2_fill_1 FILLER_50_2762 ();
 sg13g2_fill_2 FILLER_50_2841 ();
 sg13g2_decap_8 FILLER_50_2851 ();
 sg13g2_fill_2 FILLER_50_2858 ();
 sg13g2_decap_8 FILLER_50_2867 ();
 sg13g2_decap_4 FILLER_50_2874 ();
 sg13g2_fill_1 FILLER_50_2910 ();
 sg13g2_fill_2 FILLER_50_2915 ();
 sg13g2_fill_2 FILLER_50_2921 ();
 sg13g2_fill_1 FILLER_50_2923 ();
 sg13g2_decap_8 FILLER_50_2959 ();
 sg13g2_decap_4 FILLER_50_2966 ();
 sg13g2_fill_2 FILLER_50_2970 ();
 sg13g2_decap_8 FILLER_50_2981 ();
 sg13g2_decap_8 FILLER_50_2988 ();
 sg13g2_decap_8 FILLER_50_2995 ();
 sg13g2_decap_8 FILLER_50_3002 ();
 sg13g2_decap_8 FILLER_50_3009 ();
 sg13g2_decap_8 FILLER_50_3016 ();
 sg13g2_decap_8 FILLER_50_3023 ();
 sg13g2_decap_8 FILLER_50_3030 ();
 sg13g2_decap_8 FILLER_50_3037 ();
 sg13g2_decap_8 FILLER_50_3044 ();
 sg13g2_decap_8 FILLER_50_3051 ();
 sg13g2_decap_8 FILLER_50_3058 ();
 sg13g2_decap_8 FILLER_50_3065 ();
 sg13g2_decap_8 FILLER_50_3072 ();
 sg13g2_decap_8 FILLER_50_3079 ();
 sg13g2_decap_8 FILLER_50_3086 ();
 sg13g2_decap_8 FILLER_50_3093 ();
 sg13g2_decap_8 FILLER_50_3100 ();
 sg13g2_decap_8 FILLER_50_3107 ();
 sg13g2_decap_8 FILLER_50_3114 ();
 sg13g2_decap_8 FILLER_50_3121 ();
 sg13g2_decap_8 FILLER_50_3128 ();
 sg13g2_decap_8 FILLER_50_3135 ();
 sg13g2_decap_8 FILLER_50_3142 ();
 sg13g2_decap_8 FILLER_50_3149 ();
 sg13g2_decap_8 FILLER_50_3156 ();
 sg13g2_decap_8 FILLER_50_3163 ();
 sg13g2_decap_8 FILLER_50_3170 ();
 sg13g2_decap_8 FILLER_50_3177 ();
 sg13g2_decap_8 FILLER_50_3184 ();
 sg13g2_decap_8 FILLER_50_3191 ();
 sg13g2_decap_8 FILLER_50_3198 ();
 sg13g2_decap_8 FILLER_50_3205 ();
 sg13g2_decap_8 FILLER_50_3212 ();
 sg13g2_decap_8 FILLER_50_3219 ();
 sg13g2_decap_8 FILLER_50_3226 ();
 sg13g2_decap_8 FILLER_50_3233 ();
 sg13g2_decap_8 FILLER_50_3240 ();
 sg13g2_decap_8 FILLER_50_3247 ();
 sg13g2_decap_8 FILLER_50_3254 ();
 sg13g2_decap_8 FILLER_50_3261 ();
 sg13g2_decap_8 FILLER_50_3268 ();
 sg13g2_decap_8 FILLER_50_3275 ();
 sg13g2_decap_8 FILLER_50_3282 ();
 sg13g2_decap_8 FILLER_50_3289 ();
 sg13g2_decap_8 FILLER_50_3296 ();
 sg13g2_decap_8 FILLER_50_3303 ();
 sg13g2_decap_8 FILLER_50_3310 ();
 sg13g2_decap_8 FILLER_50_3317 ();
 sg13g2_decap_8 FILLER_50_3324 ();
 sg13g2_decap_8 FILLER_50_3331 ();
 sg13g2_decap_8 FILLER_50_3338 ();
 sg13g2_decap_8 FILLER_50_3345 ();
 sg13g2_decap_8 FILLER_50_3352 ();
 sg13g2_decap_8 FILLER_50_3359 ();
 sg13g2_decap_8 FILLER_50_3366 ();
 sg13g2_decap_8 FILLER_50_3373 ();
 sg13g2_decap_8 FILLER_50_3380 ();
 sg13g2_decap_8 FILLER_50_3387 ();
 sg13g2_decap_8 FILLER_50_3394 ();
 sg13g2_decap_8 FILLER_50_3401 ();
 sg13g2_decap_8 FILLER_50_3408 ();
 sg13g2_decap_8 FILLER_50_3415 ();
 sg13g2_decap_8 FILLER_50_3422 ();
 sg13g2_decap_8 FILLER_50_3429 ();
 sg13g2_decap_8 FILLER_50_3436 ();
 sg13g2_decap_8 FILLER_50_3443 ();
 sg13g2_decap_8 FILLER_50_3450 ();
 sg13g2_decap_8 FILLER_50_3457 ();
 sg13g2_decap_8 FILLER_50_3464 ();
 sg13g2_decap_8 FILLER_50_3471 ();
 sg13g2_decap_8 FILLER_50_3478 ();
 sg13g2_decap_8 FILLER_50_3485 ();
 sg13g2_decap_8 FILLER_50_3492 ();
 sg13g2_decap_8 FILLER_50_3499 ();
 sg13g2_decap_8 FILLER_50_3506 ();
 sg13g2_decap_8 FILLER_50_3513 ();
 sg13g2_decap_8 FILLER_50_3520 ();
 sg13g2_decap_8 FILLER_50_3527 ();
 sg13g2_decap_8 FILLER_50_3534 ();
 sg13g2_decap_8 FILLER_50_3541 ();
 sg13g2_decap_8 FILLER_50_3548 ();
 sg13g2_decap_8 FILLER_50_3555 ();
 sg13g2_decap_8 FILLER_50_3562 ();
 sg13g2_decap_8 FILLER_50_3569 ();
 sg13g2_decap_4 FILLER_50_3576 ();
 sg13g2_fill_2 FILLER_51_26 ();
 sg13g2_fill_1 FILLER_51_28 ();
 sg13g2_fill_2 FILLER_51_72 ();
 sg13g2_fill_1 FILLER_51_74 ();
 sg13g2_fill_1 FILLER_51_79 ();
 sg13g2_fill_1 FILLER_51_115 ();
 sg13g2_decap_8 FILLER_51_150 ();
 sg13g2_decap_8 FILLER_51_161 ();
 sg13g2_decap_4 FILLER_51_168 ();
 sg13g2_fill_2 FILLER_51_172 ();
 sg13g2_decap_4 FILLER_51_179 ();
 sg13g2_decap_4 FILLER_51_230 ();
 sg13g2_fill_2 FILLER_51_262 ();
 sg13g2_decap_8 FILLER_51_274 ();
 sg13g2_decap_8 FILLER_51_281 ();
 sg13g2_decap_4 FILLER_51_288 ();
 sg13g2_decap_8 FILLER_51_305 ();
 sg13g2_fill_1 FILLER_51_326 ();
 sg13g2_decap_8 FILLER_51_345 ();
 sg13g2_fill_2 FILLER_51_357 ();
 sg13g2_fill_1 FILLER_51_359 ();
 sg13g2_fill_2 FILLER_51_418 ();
 sg13g2_fill_1 FILLER_51_420 ();
 sg13g2_decap_4 FILLER_51_441 ();
 sg13g2_fill_2 FILLER_51_445 ();
 sg13g2_fill_1 FILLER_51_451 ();
 sg13g2_decap_8 FILLER_51_461 ();
 sg13g2_decap_8 FILLER_51_468 ();
 sg13g2_fill_2 FILLER_51_475 ();
 sg13g2_fill_2 FILLER_51_514 ();
 sg13g2_decap_4 FILLER_51_521 ();
 sg13g2_fill_1 FILLER_51_542 ();
 sg13g2_fill_1 FILLER_51_563 ();
 sg13g2_decap_8 FILLER_51_568 ();
 sg13g2_fill_1 FILLER_51_575 ();
 sg13g2_fill_1 FILLER_51_617 ();
 sg13g2_fill_2 FILLER_51_626 ();
 sg13g2_fill_2 FILLER_51_642 ();
 sg13g2_fill_2 FILLER_51_662 ();
 sg13g2_fill_1 FILLER_51_664 ();
 sg13g2_fill_2 FILLER_51_673 ();
 sg13g2_decap_4 FILLER_51_697 ();
 sg13g2_fill_2 FILLER_51_701 ();
 sg13g2_fill_1 FILLER_51_721 ();
 sg13g2_decap_4 FILLER_51_727 ();
 sg13g2_decap_4 FILLER_51_772 ();
 sg13g2_fill_1 FILLER_51_776 ();
 sg13g2_fill_2 FILLER_51_786 ();
 sg13g2_fill_1 FILLER_51_788 ();
 sg13g2_fill_1 FILLER_51_803 ();
 sg13g2_fill_2 FILLER_51_813 ();
 sg13g2_fill_1 FILLER_51_815 ();
 sg13g2_decap_4 FILLER_51_821 ();
 sg13g2_decap_4 FILLER_51_829 ();
 sg13g2_fill_1 FILLER_51_897 ();
 sg13g2_fill_2 FILLER_51_911 ();
 sg13g2_fill_2 FILLER_51_923 ();
 sg13g2_fill_1 FILLER_51_942 ();
 sg13g2_fill_1 FILLER_51_952 ();
 sg13g2_fill_2 FILLER_51_958 ();
 sg13g2_decap_8 FILLER_51_970 ();
 sg13g2_fill_1 FILLER_51_977 ();
 sg13g2_fill_2 FILLER_51_991 ();
 sg13g2_fill_1 FILLER_51_1019 ();
 sg13g2_fill_2 FILLER_51_1029 ();
 sg13g2_fill_2 FILLER_51_1060 ();
 sg13g2_fill_1 FILLER_51_1062 ();
 sg13g2_decap_4 FILLER_51_1115 ();
 sg13g2_decap_8 FILLER_51_1176 ();
 sg13g2_decap_8 FILLER_51_1183 ();
 sg13g2_fill_1 FILLER_51_1190 ();
 sg13g2_decap_4 FILLER_51_1195 ();
 sg13g2_fill_2 FILLER_51_1199 ();
 sg13g2_fill_2 FILLER_51_1210 ();
 sg13g2_fill_1 FILLER_51_1212 ();
 sg13g2_decap_8 FILLER_51_1226 ();
 sg13g2_decap_8 FILLER_51_1233 ();
 sg13g2_fill_1 FILLER_51_1240 ();
 sg13g2_decap_4 FILLER_51_1255 ();
 sg13g2_decap_8 FILLER_51_1284 ();
 sg13g2_fill_1 FILLER_51_1291 ();
 sg13g2_fill_2 FILLER_51_1323 ();
 sg13g2_fill_1 FILLER_51_1325 ();
 sg13g2_decap_4 FILLER_51_1352 ();
 sg13g2_fill_1 FILLER_51_1356 ();
 sg13g2_decap_8 FILLER_51_1388 ();
 sg13g2_fill_2 FILLER_51_1395 ();
 sg13g2_decap_8 FILLER_51_1407 ();
 sg13g2_decap_4 FILLER_51_1414 ();
 sg13g2_decap_8 FILLER_51_1422 ();
 sg13g2_fill_2 FILLER_51_1429 ();
 sg13g2_fill_1 FILLER_51_1441 ();
 sg13g2_decap_4 FILLER_51_1468 ();
 sg13g2_decap_8 FILLER_51_1481 ();
 sg13g2_decap_4 FILLER_51_1488 ();
 sg13g2_fill_1 FILLER_51_1492 ();
 sg13g2_decap_4 FILLER_51_1497 ();
 sg13g2_fill_1 FILLER_51_1511 ();
 sg13g2_decap_8 FILLER_51_1533 ();
 sg13g2_decap_8 FILLER_51_1540 ();
 sg13g2_fill_2 FILLER_51_1547 ();
 sg13g2_fill_1 FILLER_51_1560 ();
 sg13g2_decap_8 FILLER_51_1575 ();
 sg13g2_fill_1 FILLER_51_1582 ();
 sg13g2_fill_1 FILLER_51_1588 ();
 sg13g2_fill_2 FILLER_51_1593 ();
 sg13g2_fill_1 FILLER_51_1595 ();
 sg13g2_fill_2 FILLER_51_1604 ();
 sg13g2_fill_1 FILLER_51_1606 ();
 sg13g2_decap_8 FILLER_51_1612 ();
 sg13g2_decap_8 FILLER_51_1619 ();
 sg13g2_fill_2 FILLER_51_1626 ();
 sg13g2_fill_1 FILLER_51_1628 ();
 sg13g2_fill_1 FILLER_51_1650 ();
 sg13g2_decap_8 FILLER_51_1673 ();
 sg13g2_fill_2 FILLER_51_1680 ();
 sg13g2_decap_8 FILLER_51_1708 ();
 sg13g2_fill_2 FILLER_51_1715 ();
 sg13g2_decap_8 FILLER_51_1733 ();
 sg13g2_decap_8 FILLER_51_1740 ();
 sg13g2_decap_8 FILLER_51_1747 ();
 sg13g2_decap_4 FILLER_51_1754 ();
 sg13g2_fill_1 FILLER_51_1758 ();
 sg13g2_decap_8 FILLER_51_1773 ();
 sg13g2_fill_1 FILLER_51_1780 ();
 sg13g2_decap_8 FILLER_51_1802 ();
 sg13g2_decap_8 FILLER_51_1809 ();
 sg13g2_fill_1 FILLER_51_1816 ();
 sg13g2_fill_2 FILLER_51_1843 ();
 sg13g2_decap_8 FILLER_51_1867 ();
 sg13g2_decap_8 FILLER_51_1874 ();
 sg13g2_decap_4 FILLER_51_1881 ();
 sg13g2_fill_2 FILLER_51_1885 ();
 sg13g2_decap_8 FILLER_51_1927 ();
 sg13g2_decap_4 FILLER_51_1934 ();
 sg13g2_fill_1 FILLER_51_1938 ();
 sg13g2_fill_1 FILLER_51_1949 ();
 sg13g2_fill_1 FILLER_51_1955 ();
 sg13g2_decap_4 FILLER_51_1967 ();
 sg13g2_fill_2 FILLER_51_1987 ();
 sg13g2_decap_8 FILLER_51_2008 ();
 sg13g2_decap_8 FILLER_51_2015 ();
 sg13g2_fill_2 FILLER_51_2022 ();
 sg13g2_fill_1 FILLER_51_2024 ();
 sg13g2_decap_8 FILLER_51_2038 ();
 sg13g2_fill_2 FILLER_51_2045 ();
 sg13g2_fill_1 FILLER_51_2047 ();
 sg13g2_decap_4 FILLER_51_2057 ();
 sg13g2_fill_1 FILLER_51_2061 ();
 sg13g2_fill_1 FILLER_51_2075 ();
 sg13g2_decap_4 FILLER_51_2080 ();
 sg13g2_fill_1 FILLER_51_2084 ();
 sg13g2_fill_1 FILLER_51_2105 ();
 sg13g2_decap_4 FILLER_51_2124 ();
 sg13g2_fill_2 FILLER_51_2144 ();
 sg13g2_fill_1 FILLER_51_2163 ();
 sg13g2_decap_4 FILLER_51_2169 ();
 sg13g2_fill_1 FILLER_51_2173 ();
 sg13g2_fill_2 FILLER_51_2192 ();
 sg13g2_fill_1 FILLER_51_2194 ();
 sg13g2_fill_2 FILLER_51_2216 ();
 sg13g2_fill_1 FILLER_51_2218 ();
 sg13g2_fill_1 FILLER_51_2229 ();
 sg13g2_fill_2 FILLER_51_2245 ();
 sg13g2_fill_1 FILLER_51_2247 ();
 sg13g2_decap_8 FILLER_51_2256 ();
 sg13g2_decap_4 FILLER_51_2272 ();
 sg13g2_fill_2 FILLER_51_2294 ();
 sg13g2_fill_1 FILLER_51_2296 ();
 sg13g2_decap_4 FILLER_51_2316 ();
 sg13g2_fill_1 FILLER_51_2320 ();
 sg13g2_fill_2 FILLER_51_2328 ();
 sg13g2_fill_1 FILLER_51_2334 ();
 sg13g2_fill_2 FILLER_51_2344 ();
 sg13g2_decap_4 FILLER_51_2350 ();
 sg13g2_fill_2 FILLER_51_2354 ();
 sg13g2_fill_1 FILLER_51_2363 ();
 sg13g2_decap_8 FILLER_51_2386 ();
 sg13g2_decap_8 FILLER_51_2393 ();
 sg13g2_decap_8 FILLER_51_2400 ();
 sg13g2_decap_4 FILLER_51_2407 ();
 sg13g2_fill_2 FILLER_51_2429 ();
 sg13g2_decap_8 FILLER_51_2439 ();
 sg13g2_decap_8 FILLER_51_2446 ();
 sg13g2_fill_1 FILLER_51_2453 ();
 sg13g2_decap_8 FILLER_51_2466 ();
 sg13g2_fill_2 FILLER_51_2473 ();
 sg13g2_fill_1 FILLER_51_2475 ();
 sg13g2_fill_2 FILLER_51_2481 ();
 sg13g2_fill_1 FILLER_51_2483 ();
 sg13g2_decap_8 FILLER_51_2494 ();
 sg13g2_decap_8 FILLER_51_2501 ();
 sg13g2_fill_2 FILLER_51_2508 ();
 sg13g2_fill_2 FILLER_51_2519 ();
 sg13g2_fill_1 FILLER_51_2567 ();
 sg13g2_decap_4 FILLER_51_2594 ();
 sg13g2_decap_8 FILLER_51_2608 ();
 sg13g2_fill_1 FILLER_51_2624 ();
 sg13g2_decap_4 FILLER_51_2629 ();
 sg13g2_fill_2 FILLER_51_2642 ();
 sg13g2_fill_1 FILLER_51_2644 ();
 sg13g2_decap_4 FILLER_51_2649 ();
 sg13g2_fill_1 FILLER_51_2653 ();
 sg13g2_fill_2 FILLER_51_2674 ();
 sg13g2_fill_1 FILLER_51_2676 ();
 sg13g2_fill_1 FILLER_51_2703 ();
 sg13g2_fill_2 FILLER_51_2713 ();
 sg13g2_fill_2 FILLER_51_2724 ();
 sg13g2_fill_1 FILLER_51_2739 ();
 sg13g2_fill_2 FILLER_51_2766 ();
 sg13g2_decap_4 FILLER_51_2781 ();
 sg13g2_fill_2 FILLER_51_2785 ();
 sg13g2_fill_1 FILLER_51_2791 ();
 sg13g2_fill_2 FILLER_51_2810 ();
 sg13g2_fill_2 FILLER_51_2838 ();
 sg13g2_decap_4 FILLER_51_2844 ();
 sg13g2_fill_1 FILLER_51_2848 ();
 sg13g2_fill_2 FILLER_51_2887 ();
 sg13g2_fill_2 FILLER_51_2893 ();
 sg13g2_fill_2 FILLER_51_2919 ();
 sg13g2_fill_2 FILLER_51_2929 ();
 sg13g2_fill_1 FILLER_51_2931 ();
 sg13g2_fill_2 FILLER_51_2946 ();
 sg13g2_fill_1 FILLER_51_2953 ();
 sg13g2_fill_2 FILLER_51_2961 ();
 sg13g2_decap_8 FILLER_51_2989 ();
 sg13g2_decap_8 FILLER_51_2996 ();
 sg13g2_decap_8 FILLER_51_3003 ();
 sg13g2_decap_8 FILLER_51_3010 ();
 sg13g2_decap_8 FILLER_51_3017 ();
 sg13g2_decap_8 FILLER_51_3024 ();
 sg13g2_decap_8 FILLER_51_3031 ();
 sg13g2_decap_8 FILLER_51_3038 ();
 sg13g2_decap_8 FILLER_51_3045 ();
 sg13g2_decap_8 FILLER_51_3052 ();
 sg13g2_decap_8 FILLER_51_3059 ();
 sg13g2_decap_8 FILLER_51_3066 ();
 sg13g2_decap_8 FILLER_51_3073 ();
 sg13g2_decap_8 FILLER_51_3080 ();
 sg13g2_decap_8 FILLER_51_3087 ();
 sg13g2_decap_8 FILLER_51_3094 ();
 sg13g2_decap_8 FILLER_51_3101 ();
 sg13g2_decap_8 FILLER_51_3108 ();
 sg13g2_decap_8 FILLER_51_3115 ();
 sg13g2_decap_8 FILLER_51_3122 ();
 sg13g2_decap_8 FILLER_51_3129 ();
 sg13g2_decap_8 FILLER_51_3136 ();
 sg13g2_decap_8 FILLER_51_3143 ();
 sg13g2_decap_8 FILLER_51_3150 ();
 sg13g2_decap_8 FILLER_51_3157 ();
 sg13g2_decap_8 FILLER_51_3164 ();
 sg13g2_decap_8 FILLER_51_3171 ();
 sg13g2_decap_8 FILLER_51_3178 ();
 sg13g2_decap_8 FILLER_51_3185 ();
 sg13g2_decap_8 FILLER_51_3192 ();
 sg13g2_decap_8 FILLER_51_3199 ();
 sg13g2_decap_8 FILLER_51_3206 ();
 sg13g2_decap_8 FILLER_51_3213 ();
 sg13g2_decap_8 FILLER_51_3220 ();
 sg13g2_decap_8 FILLER_51_3227 ();
 sg13g2_decap_8 FILLER_51_3234 ();
 sg13g2_decap_8 FILLER_51_3241 ();
 sg13g2_decap_8 FILLER_51_3248 ();
 sg13g2_decap_8 FILLER_51_3255 ();
 sg13g2_decap_8 FILLER_51_3262 ();
 sg13g2_decap_8 FILLER_51_3269 ();
 sg13g2_decap_8 FILLER_51_3276 ();
 sg13g2_decap_8 FILLER_51_3283 ();
 sg13g2_decap_8 FILLER_51_3290 ();
 sg13g2_decap_8 FILLER_51_3297 ();
 sg13g2_decap_8 FILLER_51_3304 ();
 sg13g2_decap_8 FILLER_51_3311 ();
 sg13g2_decap_8 FILLER_51_3318 ();
 sg13g2_decap_8 FILLER_51_3325 ();
 sg13g2_decap_8 FILLER_51_3332 ();
 sg13g2_decap_8 FILLER_51_3339 ();
 sg13g2_decap_8 FILLER_51_3346 ();
 sg13g2_decap_8 FILLER_51_3353 ();
 sg13g2_decap_8 FILLER_51_3360 ();
 sg13g2_decap_8 FILLER_51_3367 ();
 sg13g2_decap_8 FILLER_51_3374 ();
 sg13g2_decap_8 FILLER_51_3381 ();
 sg13g2_decap_8 FILLER_51_3388 ();
 sg13g2_decap_8 FILLER_51_3395 ();
 sg13g2_decap_8 FILLER_51_3402 ();
 sg13g2_decap_8 FILLER_51_3409 ();
 sg13g2_decap_8 FILLER_51_3416 ();
 sg13g2_decap_8 FILLER_51_3423 ();
 sg13g2_decap_8 FILLER_51_3430 ();
 sg13g2_decap_8 FILLER_51_3437 ();
 sg13g2_decap_8 FILLER_51_3444 ();
 sg13g2_decap_8 FILLER_51_3451 ();
 sg13g2_decap_8 FILLER_51_3458 ();
 sg13g2_decap_8 FILLER_51_3465 ();
 sg13g2_decap_8 FILLER_51_3472 ();
 sg13g2_decap_8 FILLER_51_3479 ();
 sg13g2_decap_8 FILLER_51_3486 ();
 sg13g2_decap_8 FILLER_51_3493 ();
 sg13g2_decap_8 FILLER_51_3500 ();
 sg13g2_decap_8 FILLER_51_3507 ();
 sg13g2_decap_8 FILLER_51_3514 ();
 sg13g2_decap_8 FILLER_51_3521 ();
 sg13g2_decap_8 FILLER_51_3528 ();
 sg13g2_decap_8 FILLER_51_3535 ();
 sg13g2_decap_8 FILLER_51_3542 ();
 sg13g2_decap_8 FILLER_51_3549 ();
 sg13g2_decap_8 FILLER_51_3556 ();
 sg13g2_decap_8 FILLER_51_3563 ();
 sg13g2_decap_8 FILLER_51_3570 ();
 sg13g2_fill_2 FILLER_51_3577 ();
 sg13g2_fill_1 FILLER_51_3579 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_4 FILLER_52_14 ();
 sg13g2_fill_1 FILLER_52_18 ();
 sg13g2_fill_2 FILLER_52_45 ();
 sg13g2_fill_1 FILLER_52_47 ();
 sg13g2_fill_1 FILLER_52_65 ();
 sg13g2_decap_8 FILLER_52_71 ();
 sg13g2_decap_4 FILLER_52_78 ();
 sg13g2_decap_8 FILLER_52_105 ();
 sg13g2_fill_1 FILLER_52_112 ();
 sg13g2_decap_4 FILLER_52_193 ();
 sg13g2_fill_2 FILLER_52_224 ();
 sg13g2_fill_1 FILLER_52_226 ();
 sg13g2_fill_1 FILLER_52_266 ();
 sg13g2_fill_1 FILLER_52_273 ();
 sg13g2_fill_2 FILLER_52_310 ();
 sg13g2_fill_1 FILLER_52_312 ();
 sg13g2_decap_4 FILLER_52_339 ();
 sg13g2_fill_2 FILLER_52_360 ();
 sg13g2_fill_1 FILLER_52_362 ();
 sg13g2_decap_4 FILLER_52_377 ();
 sg13g2_fill_2 FILLER_52_381 ();
 sg13g2_decap_4 FILLER_52_409 ();
 sg13g2_fill_2 FILLER_52_413 ();
 sg13g2_decap_8 FILLER_52_418 ();
 sg13g2_fill_2 FILLER_52_467 ();
 sg13g2_fill_1 FILLER_52_469 ();
 sg13g2_decap_8 FILLER_52_474 ();
 sg13g2_decap_4 FILLER_52_481 ();
 sg13g2_fill_2 FILLER_52_485 ();
 sg13g2_fill_2 FILLER_52_494 ();
 sg13g2_fill_2 FILLER_52_510 ();
 sg13g2_fill_2 FILLER_52_538 ();
 sg13g2_fill_2 FILLER_52_549 ();
 sg13g2_fill_2 FILLER_52_581 ();
 sg13g2_fill_1 FILLER_52_583 ();
 sg13g2_fill_2 FILLER_52_598 ();
 sg13g2_fill_1 FILLER_52_600 ();
 sg13g2_decap_8 FILLER_52_605 ();
 sg13g2_decap_4 FILLER_52_612 ();
 sg13g2_fill_2 FILLER_52_616 ();
 sg13g2_decap_8 FILLER_52_631 ();
 sg13g2_decap_8 FILLER_52_638 ();
 sg13g2_fill_1 FILLER_52_645 ();
 sg13g2_fill_2 FILLER_52_667 ();
 sg13g2_fill_2 FILLER_52_733 ();
 sg13g2_fill_1 FILLER_52_735 ();
 sg13g2_decap_4 FILLER_52_746 ();
 sg13g2_fill_1 FILLER_52_750 ();
 sg13g2_fill_1 FILLER_52_759 ();
 sg13g2_fill_2 FILLER_52_788 ();
 sg13g2_fill_2 FILLER_52_816 ();
 sg13g2_fill_1 FILLER_52_818 ();
 sg13g2_fill_2 FILLER_52_852 ();
 sg13g2_decap_4 FILLER_52_892 ();
 sg13g2_decap_4 FILLER_52_912 ();
 sg13g2_fill_1 FILLER_52_916 ();
 sg13g2_fill_2 FILLER_52_943 ();
 sg13g2_decap_8 FILLER_52_958 ();
 sg13g2_decap_4 FILLER_52_965 ();
 sg13g2_decap_8 FILLER_52_979 ();
 sg13g2_fill_2 FILLER_52_986 ();
 sg13g2_fill_2 FILLER_52_1008 ();
 sg13g2_fill_2 FILLER_52_1019 ();
 sg13g2_fill_1 FILLER_52_1040 ();
 sg13g2_fill_2 FILLER_52_1076 ();
 sg13g2_fill_1 FILLER_52_1078 ();
 sg13g2_fill_2 FILLER_52_1088 ();
 sg13g2_fill_1 FILLER_52_1090 ();
 sg13g2_fill_2 FILLER_52_1110 ();
 sg13g2_fill_2 FILLER_52_1121 ();
 sg13g2_fill_1 FILLER_52_1123 ();
 sg13g2_fill_1 FILLER_52_1148 ();
 sg13g2_decap_4 FILLER_52_1170 ();
 sg13g2_fill_2 FILLER_52_1174 ();
 sg13g2_fill_1 FILLER_52_1184 ();
 sg13g2_fill_1 FILLER_52_1215 ();
 sg13g2_fill_1 FILLER_52_1225 ();
 sg13g2_fill_2 FILLER_52_1252 ();
 sg13g2_fill_2 FILLER_52_1259 ();
 sg13g2_fill_1 FILLER_52_1261 ();
 sg13g2_decap_8 FILLER_52_1270 ();
 sg13g2_decap_4 FILLER_52_1277 ();
 sg13g2_fill_1 FILLER_52_1281 ();
 sg13g2_fill_2 FILLER_52_1290 ();
 sg13g2_fill_1 FILLER_52_1292 ();
 sg13g2_decap_8 FILLER_52_1298 ();
 sg13g2_decap_4 FILLER_52_1332 ();
 sg13g2_fill_1 FILLER_52_1336 ();
 sg13g2_decap_8 FILLER_52_1341 ();
 sg13g2_fill_1 FILLER_52_1348 ();
 sg13g2_decap_8 FILLER_52_1353 ();
 sg13g2_decap_8 FILLER_52_1360 ();
 sg13g2_decap_8 FILLER_52_1367 ();
 sg13g2_fill_2 FILLER_52_1374 ();
 sg13g2_decap_8 FILLER_52_1384 ();
 sg13g2_fill_1 FILLER_52_1391 ();
 sg13g2_decap_4 FILLER_52_1402 ();
 sg13g2_decap_4 FILLER_52_1458 ();
 sg13g2_decap_4 FILLER_52_1472 ();
 sg13g2_decap_8 FILLER_52_1508 ();
 sg13g2_decap_8 FILLER_52_1515 ();
 sg13g2_decap_8 FILLER_52_1522 ();
 sg13g2_fill_2 FILLER_52_1529 ();
 sg13g2_fill_1 FILLER_52_1531 ();
 sg13g2_decap_8 FILLER_52_1540 ();
 sg13g2_fill_1 FILLER_52_1547 ();
 sg13g2_decap_4 FILLER_52_1556 ();
 sg13g2_decap_4 FILLER_52_1564 ();
 sg13g2_fill_2 FILLER_52_1568 ();
 sg13g2_fill_2 FILLER_52_1591 ();
 sg13g2_fill_1 FILLER_52_1593 ();
 sg13g2_decap_8 FILLER_52_1623 ();
 sg13g2_decap_4 FILLER_52_1630 ();
 sg13g2_fill_2 FILLER_52_1634 ();
 sg13g2_fill_1 FILLER_52_1654 ();
 sg13g2_decap_8 FILLER_52_1660 ();
 sg13g2_decap_8 FILLER_52_1667 ();
 sg13g2_decap_4 FILLER_52_1674 ();
 sg13g2_fill_1 FILLER_52_1678 ();
 sg13g2_decap_4 FILLER_52_1685 ();
 sg13g2_fill_2 FILLER_52_1695 ();
 sg13g2_fill_1 FILLER_52_1697 ();
 sg13g2_decap_4 FILLER_52_1708 ();
 sg13g2_fill_2 FILLER_52_1718 ();
 sg13g2_fill_2 FILLER_52_1734 ();
 sg13g2_fill_2 FILLER_52_1759 ();
 sg13g2_fill_2 FILLER_52_1779 ();
 sg13g2_decap_8 FILLER_52_1797 ();
 sg13g2_fill_1 FILLER_52_1804 ();
 sg13g2_decap_8 FILLER_52_1809 ();
 sg13g2_decap_8 FILLER_52_1816 ();
 sg13g2_decap_4 FILLER_52_1823 ();
 sg13g2_fill_1 FILLER_52_1827 ();
 sg13g2_fill_1 FILLER_52_1832 ();
 sg13g2_decap_8 FILLER_52_1837 ();
 sg13g2_fill_2 FILLER_52_1844 ();
 sg13g2_fill_1 FILLER_52_1846 ();
 sg13g2_fill_2 FILLER_52_1860 ();
 sg13g2_fill_1 FILLER_52_1862 ();
 sg13g2_decap_8 FILLER_52_1885 ();
 sg13g2_fill_2 FILLER_52_1892 ();
 sg13g2_fill_1 FILLER_52_1894 ();
 sg13g2_decap_8 FILLER_52_1910 ();
 sg13g2_fill_1 FILLER_52_1917 ();
 sg13g2_decap_8 FILLER_52_1943 ();
 sg13g2_fill_2 FILLER_52_1950 ();
 sg13g2_fill_1 FILLER_52_1965 ();
 sg13g2_fill_1 FILLER_52_1974 ();
 sg13g2_decap_4 FILLER_52_1980 ();
 sg13g2_fill_2 FILLER_52_1984 ();
 sg13g2_fill_1 FILLER_52_1996 ();
 sg13g2_decap_4 FILLER_52_2023 ();
 sg13g2_fill_2 FILLER_52_2038 ();
 sg13g2_decap_8 FILLER_52_2058 ();
 sg13g2_fill_2 FILLER_52_2065 ();
 sg13g2_fill_2 FILLER_52_2073 ();
 sg13g2_fill_1 FILLER_52_2075 ();
 sg13g2_decap_8 FILLER_52_2086 ();
 sg13g2_decap_8 FILLER_52_2093 ();
 sg13g2_decap_8 FILLER_52_2100 ();
 sg13g2_decap_4 FILLER_52_2112 ();
 sg13g2_decap_4 FILLER_52_2124 ();
 sg13g2_fill_2 FILLER_52_2142 ();
 sg13g2_fill_1 FILLER_52_2144 ();
 sg13g2_decap_8 FILLER_52_2151 ();
 sg13g2_decap_8 FILLER_52_2158 ();
 sg13g2_fill_2 FILLER_52_2165 ();
 sg13g2_fill_1 FILLER_52_2167 ();
 sg13g2_fill_1 FILLER_52_2175 ();
 sg13g2_decap_8 FILLER_52_2186 ();
 sg13g2_decap_4 FILLER_52_2193 ();
 sg13g2_fill_1 FILLER_52_2197 ();
 sg13g2_fill_1 FILLER_52_2213 ();
 sg13g2_fill_2 FILLER_52_2218 ();
 sg13g2_decap_8 FILLER_52_2242 ();
 sg13g2_decap_4 FILLER_52_2249 ();
 sg13g2_fill_1 FILLER_52_2253 ();
 sg13g2_fill_1 FILLER_52_2259 ();
 sg13g2_fill_2 FILLER_52_2268 ();
 sg13g2_decap_8 FILLER_52_2275 ();
 sg13g2_fill_2 FILLER_52_2290 ();
 sg13g2_fill_2 FILLER_52_2308 ();
 sg13g2_decap_4 FILLER_52_2315 ();
 sg13g2_fill_2 FILLER_52_2353 ();
 sg13g2_decap_8 FILLER_52_2381 ();
 sg13g2_fill_1 FILLER_52_2388 ();
 sg13g2_decap_8 FILLER_52_2394 ();
 sg13g2_fill_1 FILLER_52_2401 ();
 sg13g2_fill_1 FILLER_52_2415 ();
 sg13g2_fill_2 FILLER_52_2425 ();
 sg13g2_fill_1 FILLER_52_2427 ();
 sg13g2_decap_8 FILLER_52_2432 ();
 sg13g2_fill_1 FILLER_52_2439 ();
 sg13g2_decap_4 FILLER_52_2445 ();
 sg13g2_fill_1 FILLER_52_2457 ();
 sg13g2_decap_8 FILLER_52_2463 ();
 sg13g2_fill_1 FILLER_52_2470 ();
 sg13g2_decap_8 FILLER_52_2494 ();
 sg13g2_decap_8 FILLER_52_2524 ();
 sg13g2_fill_2 FILLER_52_2531 ();
 sg13g2_fill_2 FILLER_52_2537 ();
 sg13g2_fill_1 FILLER_52_2539 ();
 sg13g2_fill_2 FILLER_52_2588 ();
 sg13g2_fill_1 FILLER_52_2611 ();
 sg13g2_fill_1 FILLER_52_2632 ();
 sg13g2_fill_2 FILLER_52_2637 ();
 sg13g2_fill_1 FILLER_52_2639 ();
 sg13g2_decap_8 FILLER_52_2666 ();
 sg13g2_decap_8 FILLER_52_2673 ();
 sg13g2_decap_8 FILLER_52_2680 ();
 sg13g2_fill_1 FILLER_52_2687 ();
 sg13g2_decap_8 FILLER_52_2692 ();
 sg13g2_fill_2 FILLER_52_2713 ();
 sg13g2_decap_4 FILLER_52_2746 ();
 sg13g2_fill_1 FILLER_52_2750 ();
 sg13g2_decap_4 FILLER_52_2755 ();
 sg13g2_fill_1 FILLER_52_2759 ();
 sg13g2_decap_4 FILLER_52_2773 ();
 sg13g2_decap_4 FILLER_52_2795 ();
 sg13g2_fill_2 FILLER_52_2799 ();
 sg13g2_fill_1 FILLER_52_2806 ();
 sg13g2_decap_8 FILLER_52_2815 ();
 sg13g2_fill_2 FILLER_52_2830 ();
 sg13g2_fill_1 FILLER_52_2832 ();
 sg13g2_decap_8 FILLER_52_2838 ();
 sg13g2_decap_4 FILLER_52_2845 ();
 sg13g2_fill_2 FILLER_52_2849 ();
 sg13g2_fill_2 FILLER_52_2884 ();
 sg13g2_fill_1 FILLER_52_2886 ();
 sg13g2_decap_4 FILLER_52_2908 ();
 sg13g2_fill_1 FILLER_52_2912 ();
 sg13g2_fill_1 FILLER_52_2926 ();
 sg13g2_fill_1 FILLER_52_2948 ();
 sg13g2_fill_1 FILLER_52_2969 ();
 sg13g2_decap_8 FILLER_52_2984 ();
 sg13g2_decap_8 FILLER_52_2991 ();
 sg13g2_decap_8 FILLER_52_2998 ();
 sg13g2_decap_8 FILLER_52_3005 ();
 sg13g2_decap_8 FILLER_52_3012 ();
 sg13g2_decap_8 FILLER_52_3019 ();
 sg13g2_decap_8 FILLER_52_3026 ();
 sg13g2_decap_8 FILLER_52_3033 ();
 sg13g2_decap_8 FILLER_52_3040 ();
 sg13g2_decap_8 FILLER_52_3047 ();
 sg13g2_decap_8 FILLER_52_3054 ();
 sg13g2_decap_8 FILLER_52_3061 ();
 sg13g2_decap_8 FILLER_52_3068 ();
 sg13g2_decap_8 FILLER_52_3075 ();
 sg13g2_decap_8 FILLER_52_3082 ();
 sg13g2_decap_8 FILLER_52_3089 ();
 sg13g2_decap_8 FILLER_52_3096 ();
 sg13g2_decap_8 FILLER_52_3103 ();
 sg13g2_decap_8 FILLER_52_3110 ();
 sg13g2_decap_8 FILLER_52_3117 ();
 sg13g2_decap_8 FILLER_52_3124 ();
 sg13g2_decap_8 FILLER_52_3131 ();
 sg13g2_decap_8 FILLER_52_3138 ();
 sg13g2_decap_8 FILLER_52_3145 ();
 sg13g2_decap_8 FILLER_52_3152 ();
 sg13g2_decap_8 FILLER_52_3159 ();
 sg13g2_decap_8 FILLER_52_3166 ();
 sg13g2_decap_8 FILLER_52_3173 ();
 sg13g2_decap_8 FILLER_52_3180 ();
 sg13g2_decap_8 FILLER_52_3187 ();
 sg13g2_decap_8 FILLER_52_3194 ();
 sg13g2_decap_8 FILLER_52_3201 ();
 sg13g2_decap_8 FILLER_52_3208 ();
 sg13g2_decap_8 FILLER_52_3215 ();
 sg13g2_decap_8 FILLER_52_3222 ();
 sg13g2_decap_8 FILLER_52_3229 ();
 sg13g2_decap_8 FILLER_52_3236 ();
 sg13g2_decap_8 FILLER_52_3243 ();
 sg13g2_decap_8 FILLER_52_3250 ();
 sg13g2_decap_8 FILLER_52_3257 ();
 sg13g2_decap_8 FILLER_52_3264 ();
 sg13g2_decap_8 FILLER_52_3271 ();
 sg13g2_decap_8 FILLER_52_3278 ();
 sg13g2_decap_8 FILLER_52_3285 ();
 sg13g2_decap_8 FILLER_52_3292 ();
 sg13g2_decap_8 FILLER_52_3299 ();
 sg13g2_decap_8 FILLER_52_3306 ();
 sg13g2_decap_8 FILLER_52_3313 ();
 sg13g2_decap_8 FILLER_52_3320 ();
 sg13g2_decap_8 FILLER_52_3327 ();
 sg13g2_decap_8 FILLER_52_3334 ();
 sg13g2_decap_8 FILLER_52_3341 ();
 sg13g2_decap_8 FILLER_52_3348 ();
 sg13g2_decap_8 FILLER_52_3355 ();
 sg13g2_decap_8 FILLER_52_3362 ();
 sg13g2_decap_8 FILLER_52_3369 ();
 sg13g2_decap_8 FILLER_52_3376 ();
 sg13g2_decap_8 FILLER_52_3383 ();
 sg13g2_decap_8 FILLER_52_3390 ();
 sg13g2_decap_8 FILLER_52_3397 ();
 sg13g2_decap_8 FILLER_52_3404 ();
 sg13g2_decap_8 FILLER_52_3411 ();
 sg13g2_decap_8 FILLER_52_3418 ();
 sg13g2_decap_8 FILLER_52_3425 ();
 sg13g2_decap_8 FILLER_52_3432 ();
 sg13g2_decap_8 FILLER_52_3439 ();
 sg13g2_decap_8 FILLER_52_3446 ();
 sg13g2_decap_8 FILLER_52_3453 ();
 sg13g2_decap_8 FILLER_52_3460 ();
 sg13g2_decap_8 FILLER_52_3467 ();
 sg13g2_decap_8 FILLER_52_3474 ();
 sg13g2_decap_8 FILLER_52_3481 ();
 sg13g2_decap_8 FILLER_52_3488 ();
 sg13g2_decap_8 FILLER_52_3495 ();
 sg13g2_decap_8 FILLER_52_3502 ();
 sg13g2_decap_8 FILLER_52_3509 ();
 sg13g2_decap_8 FILLER_52_3516 ();
 sg13g2_decap_8 FILLER_52_3523 ();
 sg13g2_decap_8 FILLER_52_3530 ();
 sg13g2_decap_8 FILLER_52_3537 ();
 sg13g2_decap_8 FILLER_52_3544 ();
 sg13g2_decap_8 FILLER_52_3551 ();
 sg13g2_decap_8 FILLER_52_3558 ();
 sg13g2_decap_8 FILLER_52_3565 ();
 sg13g2_decap_8 FILLER_52_3572 ();
 sg13g2_fill_1 FILLER_52_3579 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_fill_1 FILLER_53_7 ();
 sg13g2_fill_1 FILLER_53_25 ();
 sg13g2_fill_2 FILLER_53_31 ();
 sg13g2_fill_1 FILLER_53_33 ();
 sg13g2_fill_2 FILLER_53_57 ();
 sg13g2_fill_2 FILLER_53_80 ();
 sg13g2_fill_2 FILLER_53_127 ();
 sg13g2_fill_1 FILLER_53_129 ();
 sg13g2_fill_1 FILLER_53_139 ();
 sg13g2_fill_1 FILLER_53_145 ();
 sg13g2_decap_8 FILLER_53_150 ();
 sg13g2_decap_8 FILLER_53_157 ();
 sg13g2_decap_8 FILLER_53_164 ();
 sg13g2_decap_8 FILLER_53_171 ();
 sg13g2_fill_2 FILLER_53_182 ();
 sg13g2_fill_1 FILLER_53_184 ();
 sg13g2_decap_4 FILLER_53_224 ();
 sg13g2_fill_1 FILLER_53_261 ();
 sg13g2_fill_1 FILLER_53_272 ();
 sg13g2_fill_2 FILLER_53_283 ();
 sg13g2_fill_2 FILLER_53_299 ();
 sg13g2_fill_1 FILLER_53_301 ();
 sg13g2_fill_2 FILLER_53_315 ();
 sg13g2_fill_1 FILLER_53_317 ();
 sg13g2_fill_1 FILLER_53_323 ();
 sg13g2_fill_1 FILLER_53_328 ();
 sg13g2_fill_2 FILLER_53_350 ();
 sg13g2_fill_2 FILLER_53_369 ();
 sg13g2_fill_1 FILLER_53_393 ();
 sg13g2_fill_2 FILLER_53_398 ();
 sg13g2_fill_1 FILLER_53_400 ();
 sg13g2_decap_8 FILLER_53_424 ();
 sg13g2_fill_1 FILLER_53_431 ();
 sg13g2_fill_2 FILLER_53_435 ();
 sg13g2_fill_2 FILLER_53_442 ();
 sg13g2_fill_1 FILLER_53_444 ();
 sg13g2_decap_4 FILLER_53_485 ();
 sg13g2_fill_2 FILLER_53_489 ();
 sg13g2_fill_1 FILLER_53_537 ();
 sg13g2_fill_1 FILLER_53_548 ();
 sg13g2_fill_2 FILLER_53_559 ();
 sg13g2_decap_8 FILLER_53_565 ();
 sg13g2_fill_1 FILLER_53_572 ();
 sg13g2_fill_2 FILLER_53_599 ();
 sg13g2_fill_1 FILLER_53_601 ();
 sg13g2_fill_2 FILLER_53_605 ();
 sg13g2_fill_1 FILLER_53_607 ();
 sg13g2_fill_2 FILLER_53_620 ();
 sg13g2_decap_8 FILLER_53_626 ();
 sg13g2_decap_8 FILLER_53_633 ();
 sg13g2_decap_8 FILLER_53_640 ();
 sg13g2_fill_1 FILLER_53_673 ();
 sg13g2_fill_1 FILLER_53_677 ();
 sg13g2_fill_1 FILLER_53_692 ();
 sg13g2_decap_8 FILLER_53_698 ();
 sg13g2_fill_1 FILLER_53_705 ();
 sg13g2_decap_8 FILLER_53_719 ();
 sg13g2_fill_1 FILLER_53_726 ();
 sg13g2_fill_1 FILLER_53_732 ();
 sg13g2_decap_8 FILLER_53_749 ();
 sg13g2_decap_4 FILLER_53_756 ();
 sg13g2_fill_1 FILLER_53_825 ();
 sg13g2_fill_1 FILLER_53_854 ();
 sg13g2_fill_2 FILLER_53_892 ();
 sg13g2_decap_8 FILLER_53_932 ();
 sg13g2_fill_2 FILLER_53_939 ();
 sg13g2_fill_1 FILLER_53_941 ();
 sg13g2_decap_8 FILLER_53_948 ();
 sg13g2_fill_2 FILLER_53_955 ();
 sg13g2_fill_2 FILLER_53_988 ();
 sg13g2_fill_1 FILLER_53_990 ();
 sg13g2_fill_1 FILLER_53_1026 ();
 sg13g2_fill_1 FILLER_53_1032 ();
 sg13g2_fill_2 FILLER_53_1051 ();
 sg13g2_fill_1 FILLER_53_1053 ();
 sg13g2_fill_1 FILLER_53_1077 ();
 sg13g2_fill_2 FILLER_53_1082 ();
 sg13g2_fill_1 FILLER_53_1089 ();
 sg13g2_fill_2 FILLER_53_1100 ();
 sg13g2_fill_2 FILLER_53_1115 ();
 sg13g2_fill_2 FILLER_53_1123 ();
 sg13g2_fill_1 FILLER_53_1125 ();
 sg13g2_fill_2 FILLER_53_1139 ();
 sg13g2_fill_1 FILLER_53_1141 ();
 sg13g2_decap_8 FILLER_53_1152 ();
 sg13g2_fill_1 FILLER_53_1159 ();
 sg13g2_decap_4 FILLER_53_1164 ();
 sg13g2_fill_2 FILLER_53_1176 ();
 sg13g2_decap_8 FILLER_53_1183 ();
 sg13g2_decap_8 FILLER_53_1222 ();
 sg13g2_fill_2 FILLER_53_1229 ();
 sg13g2_fill_1 FILLER_53_1231 ();
 sg13g2_fill_2 FILLER_53_1249 ();
 sg13g2_decap_8 FILLER_53_1296 ();
 sg13g2_decap_4 FILLER_53_1303 ();
 sg13g2_decap_4 FILLER_53_1312 ();
 sg13g2_decap_4 FILLER_53_1321 ();
 sg13g2_fill_2 FILLER_53_1325 ();
 sg13g2_decap_4 FILLER_53_1364 ();
 sg13g2_decap_4 FILLER_53_1381 ();
 sg13g2_fill_1 FILLER_53_1385 ();
 sg13g2_fill_1 FILLER_53_1399 ();
 sg13g2_decap_8 FILLER_53_1424 ();
 sg13g2_decap_4 FILLER_53_1431 ();
 sg13g2_decap_4 FILLER_53_1439 ();
 sg13g2_decap_8 FILLER_53_1447 ();
 sg13g2_decap_4 FILLER_53_1454 ();
 sg13g2_decap_8 FILLER_53_1473 ();
 sg13g2_decap_4 FILLER_53_1480 ();
 sg13g2_fill_1 FILLER_53_1484 ();
 sg13g2_decap_8 FILLER_53_1490 ();
 sg13g2_fill_2 FILLER_53_1497 ();
 sg13g2_fill_2 FILLER_53_1531 ();
 sg13g2_fill_1 FILLER_53_1533 ();
 sg13g2_decap_4 FILLER_53_1564 ();
 sg13g2_fill_2 FILLER_53_1568 ();
 sg13g2_decap_4 FILLER_53_1587 ();
 sg13g2_fill_1 FILLER_53_1591 ();
 sg13g2_fill_2 FILLER_53_1600 ();
 sg13g2_decap_8 FILLER_53_1654 ();
 sg13g2_decap_4 FILLER_53_1661 ();
 sg13g2_decap_4 FILLER_53_1675 ();
 sg13g2_fill_2 FILLER_53_1679 ();
 sg13g2_decap_4 FILLER_53_1695 ();
 sg13g2_fill_2 FILLER_53_1699 ();
 sg13g2_fill_2 FILLER_53_1706 ();
 sg13g2_fill_1 FILLER_53_1708 ();
 sg13g2_decap_8 FILLER_53_1729 ();
 sg13g2_decap_8 FILLER_53_1736 ();
 sg13g2_fill_2 FILLER_53_1755 ();
 sg13g2_decap_8 FILLER_53_1778 ();
 sg13g2_decap_8 FILLER_53_1785 ();
 sg13g2_fill_2 FILLER_53_1792 ();
 sg13g2_decap_4 FILLER_53_1820 ();
 sg13g2_fill_2 FILLER_53_1837 ();
 sg13g2_fill_1 FILLER_53_1839 ();
 sg13g2_decap_8 FILLER_53_1845 ();
 sg13g2_decap_8 FILLER_53_1852 ();
 sg13g2_fill_2 FILLER_53_1859 ();
 sg13g2_decap_8 FILLER_53_1886 ();
 sg13g2_decap_4 FILLER_53_1893 ();
 sg13g2_fill_1 FILLER_53_1897 ();
 sg13g2_decap_8 FILLER_53_1906 ();
 sg13g2_fill_2 FILLER_53_1913 ();
 sg13g2_fill_1 FILLER_53_1915 ();
 sg13g2_fill_2 FILLER_53_1940 ();
 sg13g2_fill_2 FILLER_53_1946 ();
 sg13g2_fill_1 FILLER_53_1948 ();
 sg13g2_decap_8 FILLER_53_1953 ();
 sg13g2_fill_2 FILLER_53_1960 ();
 sg13g2_decap_8 FILLER_53_1996 ();
 sg13g2_fill_2 FILLER_53_2003 ();
 sg13g2_fill_1 FILLER_53_2005 ();
 sg13g2_decap_8 FILLER_53_2011 ();
 sg13g2_decap_4 FILLER_53_2018 ();
 sg13g2_fill_2 FILLER_53_2022 ();
 sg13g2_decap_8 FILLER_53_2036 ();
 sg13g2_decap_4 FILLER_53_2043 ();
 sg13g2_fill_1 FILLER_53_2047 ();
 sg13g2_fill_2 FILLER_53_2063 ();
 sg13g2_fill_1 FILLER_53_2065 ();
 sg13g2_fill_2 FILLER_53_2070 ();
 sg13g2_decap_8 FILLER_53_2076 ();
 sg13g2_decap_8 FILLER_53_2091 ();
 sg13g2_fill_1 FILLER_53_2098 ();
 sg13g2_decap_8 FILLER_53_2118 ();
 sg13g2_fill_2 FILLER_53_2125 ();
 sg13g2_fill_2 FILLER_53_2136 ();
 sg13g2_fill_1 FILLER_53_2138 ();
 sg13g2_decap_4 FILLER_53_2152 ();
 sg13g2_fill_1 FILLER_53_2156 ();
 sg13g2_fill_2 FILLER_53_2191 ();
 sg13g2_fill_1 FILLER_53_2193 ();
 sg13g2_decap_8 FILLER_53_2208 ();
 sg13g2_decap_8 FILLER_53_2215 ();
 sg13g2_decap_4 FILLER_53_2222 ();
 sg13g2_fill_2 FILLER_53_2230 ();
 sg13g2_decap_8 FILLER_53_2240 ();
 sg13g2_fill_2 FILLER_53_2255 ();
 sg13g2_fill_2 FILLER_53_2278 ();
 sg13g2_fill_1 FILLER_53_2280 ();
 sg13g2_decap_8 FILLER_53_2286 ();
 sg13g2_fill_2 FILLER_53_2293 ();
 sg13g2_fill_1 FILLER_53_2300 ();
 sg13g2_fill_1 FILLER_53_2306 ();
 sg13g2_decap_8 FILLER_53_2317 ();
 sg13g2_decap_8 FILLER_53_2324 ();
 sg13g2_fill_2 FILLER_53_2331 ();
 sg13g2_decap_8 FILLER_53_2345 ();
 sg13g2_fill_2 FILLER_53_2352 ();
 sg13g2_fill_2 FILLER_53_2359 ();
 sg13g2_decap_4 FILLER_53_2378 ();
 sg13g2_fill_1 FILLER_53_2382 ();
 sg13g2_decap_8 FILLER_53_2399 ();
 sg13g2_fill_2 FILLER_53_2406 ();
 sg13g2_fill_1 FILLER_53_2408 ();
 sg13g2_fill_2 FILLER_53_2414 ();
 sg13g2_decap_4 FILLER_53_2428 ();
 sg13g2_fill_1 FILLER_53_2432 ();
 sg13g2_decap_4 FILLER_53_2442 ();
 sg13g2_decap_8 FILLER_53_2468 ();
 sg13g2_fill_1 FILLER_53_2475 ();
 sg13g2_fill_1 FILLER_53_2516 ();
 sg13g2_fill_1 FILLER_53_2567 ();
 sg13g2_decap_8 FILLER_53_2602 ();
 sg13g2_decap_4 FILLER_53_2624 ();
 sg13g2_fill_2 FILLER_53_2643 ();
 sg13g2_fill_1 FILLER_53_2645 ();
 sg13g2_fill_2 FILLER_53_2684 ();
 sg13g2_fill_2 FILLER_53_2696 ();
 sg13g2_decap_4 FILLER_53_2703 ();
 sg13g2_fill_2 FILLER_53_2707 ();
 sg13g2_decap_8 FILLER_53_2717 ();
 sg13g2_fill_2 FILLER_53_2724 ();
 sg13g2_decap_8 FILLER_53_2740 ();
 sg13g2_decap_4 FILLER_53_2747 ();
 sg13g2_fill_1 FILLER_53_2751 ();
 sg13g2_decap_4 FILLER_53_2764 ();
 sg13g2_fill_2 FILLER_53_2768 ();
 sg13g2_fill_2 FILLER_53_2823 ();
 sg13g2_fill_2 FILLER_53_2830 ();
 sg13g2_fill_2 FILLER_53_2837 ();
 sg13g2_fill_1 FILLER_53_2839 ();
 sg13g2_fill_2 FILLER_53_2849 ();
 sg13g2_fill_1 FILLER_53_2851 ();
 sg13g2_fill_2 FILLER_53_2865 ();
 sg13g2_fill_1 FILLER_53_2867 ();
 sg13g2_fill_1 FILLER_53_2889 ();
 sg13g2_decap_4 FILLER_53_2912 ();
 sg13g2_fill_1 FILLER_53_2916 ();
 sg13g2_fill_2 FILLER_53_2925 ();
 sg13g2_decap_8 FILLER_53_2940 ();
 sg13g2_decap_4 FILLER_53_2947 ();
 sg13g2_fill_1 FILLER_53_2951 ();
 sg13g2_fill_2 FILLER_53_2996 ();
 sg13g2_decap_8 FILLER_53_3024 ();
 sg13g2_decap_8 FILLER_53_3031 ();
 sg13g2_decap_4 FILLER_53_3038 ();
 sg13g2_decap_8 FILLER_53_3046 ();
 sg13g2_decap_8 FILLER_53_3053 ();
 sg13g2_decap_8 FILLER_53_3060 ();
 sg13g2_decap_8 FILLER_53_3067 ();
 sg13g2_decap_8 FILLER_53_3074 ();
 sg13g2_decap_8 FILLER_53_3081 ();
 sg13g2_decap_8 FILLER_53_3088 ();
 sg13g2_decap_8 FILLER_53_3095 ();
 sg13g2_decap_8 FILLER_53_3102 ();
 sg13g2_decap_8 FILLER_53_3109 ();
 sg13g2_decap_8 FILLER_53_3116 ();
 sg13g2_decap_8 FILLER_53_3123 ();
 sg13g2_decap_8 FILLER_53_3130 ();
 sg13g2_decap_8 FILLER_53_3137 ();
 sg13g2_decap_8 FILLER_53_3144 ();
 sg13g2_decap_8 FILLER_53_3151 ();
 sg13g2_decap_8 FILLER_53_3158 ();
 sg13g2_decap_8 FILLER_53_3165 ();
 sg13g2_decap_8 FILLER_53_3172 ();
 sg13g2_decap_8 FILLER_53_3179 ();
 sg13g2_decap_8 FILLER_53_3186 ();
 sg13g2_decap_8 FILLER_53_3193 ();
 sg13g2_decap_8 FILLER_53_3200 ();
 sg13g2_decap_8 FILLER_53_3207 ();
 sg13g2_decap_8 FILLER_53_3214 ();
 sg13g2_decap_8 FILLER_53_3221 ();
 sg13g2_decap_8 FILLER_53_3228 ();
 sg13g2_decap_8 FILLER_53_3235 ();
 sg13g2_decap_8 FILLER_53_3242 ();
 sg13g2_decap_8 FILLER_53_3249 ();
 sg13g2_decap_8 FILLER_53_3256 ();
 sg13g2_decap_8 FILLER_53_3263 ();
 sg13g2_decap_8 FILLER_53_3270 ();
 sg13g2_decap_8 FILLER_53_3277 ();
 sg13g2_decap_8 FILLER_53_3284 ();
 sg13g2_decap_8 FILLER_53_3291 ();
 sg13g2_decap_8 FILLER_53_3298 ();
 sg13g2_decap_8 FILLER_53_3305 ();
 sg13g2_decap_8 FILLER_53_3312 ();
 sg13g2_decap_8 FILLER_53_3319 ();
 sg13g2_decap_8 FILLER_53_3326 ();
 sg13g2_decap_8 FILLER_53_3333 ();
 sg13g2_decap_8 FILLER_53_3340 ();
 sg13g2_decap_8 FILLER_53_3347 ();
 sg13g2_decap_8 FILLER_53_3354 ();
 sg13g2_decap_8 FILLER_53_3361 ();
 sg13g2_decap_8 FILLER_53_3368 ();
 sg13g2_decap_8 FILLER_53_3375 ();
 sg13g2_decap_8 FILLER_53_3382 ();
 sg13g2_decap_8 FILLER_53_3389 ();
 sg13g2_decap_8 FILLER_53_3396 ();
 sg13g2_decap_8 FILLER_53_3403 ();
 sg13g2_decap_8 FILLER_53_3410 ();
 sg13g2_decap_8 FILLER_53_3417 ();
 sg13g2_decap_8 FILLER_53_3424 ();
 sg13g2_decap_8 FILLER_53_3431 ();
 sg13g2_decap_8 FILLER_53_3438 ();
 sg13g2_decap_8 FILLER_53_3445 ();
 sg13g2_decap_8 FILLER_53_3452 ();
 sg13g2_decap_8 FILLER_53_3459 ();
 sg13g2_decap_8 FILLER_53_3466 ();
 sg13g2_decap_8 FILLER_53_3473 ();
 sg13g2_decap_8 FILLER_53_3480 ();
 sg13g2_decap_8 FILLER_53_3487 ();
 sg13g2_decap_8 FILLER_53_3494 ();
 sg13g2_decap_8 FILLER_53_3501 ();
 sg13g2_decap_8 FILLER_53_3508 ();
 sg13g2_decap_8 FILLER_53_3515 ();
 sg13g2_decap_8 FILLER_53_3522 ();
 sg13g2_decap_8 FILLER_53_3529 ();
 sg13g2_decap_8 FILLER_53_3536 ();
 sg13g2_decap_8 FILLER_53_3543 ();
 sg13g2_decap_8 FILLER_53_3550 ();
 sg13g2_decap_8 FILLER_53_3557 ();
 sg13g2_decap_8 FILLER_53_3564 ();
 sg13g2_decap_8 FILLER_53_3571 ();
 sg13g2_fill_2 FILLER_53_3578 ();
 sg13g2_fill_1 FILLER_54_0 ();
 sg13g2_fill_2 FILLER_54_27 ();
 sg13g2_fill_2 FILLER_54_43 ();
 sg13g2_decap_4 FILLER_54_62 ();
 sg13g2_decap_4 FILLER_54_74 ();
 sg13g2_fill_2 FILLER_54_78 ();
 sg13g2_fill_1 FILLER_54_97 ();
 sg13g2_fill_1 FILLER_54_107 ();
 sg13g2_decap_4 FILLER_54_169 ();
 sg13g2_decap_8 FILLER_54_177 ();
 sg13g2_decap_8 FILLER_54_184 ();
 sg13g2_decap_4 FILLER_54_191 ();
 sg13g2_decap_4 FILLER_54_200 ();
 sg13g2_fill_1 FILLER_54_204 ();
 sg13g2_decap_8 FILLER_54_223 ();
 sg13g2_fill_2 FILLER_54_230 ();
 sg13g2_decap_8 FILLER_54_322 ();
 sg13g2_decap_4 FILLER_54_329 ();
 sg13g2_fill_1 FILLER_54_360 ();
 sg13g2_decap_8 FILLER_54_436 ();
 sg13g2_fill_2 FILLER_54_447 ();
 sg13g2_fill_1 FILLER_54_459 ();
 sg13g2_fill_1 FILLER_54_469 ();
 sg13g2_fill_1 FILLER_54_475 ();
 sg13g2_fill_2 FILLER_54_481 ();
 sg13g2_fill_1 FILLER_54_483 ();
 sg13g2_fill_2 FILLER_54_499 ();
 sg13g2_fill_2 FILLER_54_546 ();
 sg13g2_fill_2 FILLER_54_574 ();
 sg13g2_fill_1 FILLER_54_576 ();
 sg13g2_fill_1 FILLER_54_582 ();
 sg13g2_fill_1 FILLER_54_601 ();
 sg13g2_fill_2 FILLER_54_605 ();
 sg13g2_decap_8 FILLER_54_641 ();
 sg13g2_fill_1 FILLER_54_648 ();
 sg13g2_decap_8 FILLER_54_664 ();
 sg13g2_fill_1 FILLER_54_677 ();
 sg13g2_fill_2 FILLER_54_744 ();
 sg13g2_decap_4 FILLER_54_754 ();
 sg13g2_decap_8 FILLER_54_781 ();
 sg13g2_fill_1 FILLER_54_818 ();
 sg13g2_fill_1 FILLER_54_846 ();
 sg13g2_fill_2 FILLER_54_896 ();
 sg13g2_fill_1 FILLER_54_898 ();
 sg13g2_fill_2 FILLER_54_970 ();
 sg13g2_fill_1 FILLER_54_977 ();
 sg13g2_fill_2 FILLER_54_987 ();
 sg13g2_fill_1 FILLER_54_989 ();
 sg13g2_fill_2 FILLER_54_996 ();
 sg13g2_fill_1 FILLER_54_998 ();
 sg13g2_fill_2 FILLER_54_1005 ();
 sg13g2_fill_1 FILLER_54_1016 ();
 sg13g2_fill_1 FILLER_54_1040 ();
 sg13g2_fill_2 FILLER_54_1050 ();
 sg13g2_fill_1 FILLER_54_1078 ();
 sg13g2_fill_2 FILLER_54_1127 ();
 sg13g2_decap_4 FILLER_54_1188 ();
 sg13g2_fill_2 FILLER_54_1197 ();
 sg13g2_fill_1 FILLER_54_1199 ();
 sg13g2_fill_2 FILLER_54_1224 ();
 sg13g2_fill_1 FILLER_54_1226 ();
 sg13g2_decap_4 FILLER_54_1247 ();
 sg13g2_fill_1 FILLER_54_1251 ();
 sg13g2_fill_2 FILLER_54_1260 ();
 sg13g2_decap_8 FILLER_54_1267 ();
 sg13g2_decap_4 FILLER_54_1274 ();
 sg13g2_fill_2 FILLER_54_1278 ();
 sg13g2_decap_8 FILLER_54_1288 ();
 sg13g2_fill_2 FILLER_54_1295 ();
 sg13g2_fill_1 FILLER_54_1332 ();
 sg13g2_decap_8 FILLER_54_1357 ();
 sg13g2_decap_8 FILLER_54_1364 ();
 sg13g2_fill_2 FILLER_54_1371 ();
 sg13g2_fill_1 FILLER_54_1373 ();
 sg13g2_decap_8 FILLER_54_1378 ();
 sg13g2_decap_4 FILLER_54_1385 ();
 sg13g2_fill_1 FILLER_54_1389 ();
 sg13g2_fill_2 FILLER_54_1412 ();
 sg13g2_decap_4 FILLER_54_1419 ();
 sg13g2_decap_4 FILLER_54_1428 ();
 sg13g2_fill_1 FILLER_54_1453 ();
 sg13g2_fill_1 FILLER_54_1501 ();
 sg13g2_fill_1 FILLER_54_1514 ();
 sg13g2_decap_4 FILLER_54_1519 ();
 sg13g2_fill_1 FILLER_54_1523 ();
 sg13g2_fill_1 FILLER_54_1542 ();
 sg13g2_fill_2 FILLER_54_1546 ();
 sg13g2_fill_1 FILLER_54_1548 ();
 sg13g2_decap_4 FILLER_54_1553 ();
 sg13g2_fill_2 FILLER_54_1557 ();
 sg13g2_fill_1 FILLER_54_1564 ();
 sg13g2_decap_8 FILLER_54_1570 ();
 sg13g2_decap_8 FILLER_54_1577 ();
 sg13g2_fill_2 FILLER_54_1584 ();
 sg13g2_fill_1 FILLER_54_1586 ();
 sg13g2_decap_8 FILLER_54_1602 ();
 sg13g2_decap_8 FILLER_54_1609 ();
 sg13g2_decap_8 FILLER_54_1616 ();
 sg13g2_fill_2 FILLER_54_1623 ();
 sg13g2_fill_1 FILLER_54_1625 ();
 sg13g2_fill_2 FILLER_54_1631 ();
 sg13g2_decap_8 FILLER_54_1648 ();
 sg13g2_fill_1 FILLER_54_1655 ();
 sg13g2_fill_2 FILLER_54_1683 ();
 sg13g2_fill_1 FILLER_54_1685 ();
 sg13g2_fill_2 FILLER_54_1692 ();
 sg13g2_fill_1 FILLER_54_1694 ();
 sg13g2_decap_8 FILLER_54_1706 ();
 sg13g2_decap_4 FILLER_54_1713 ();
 sg13g2_fill_2 FILLER_54_1717 ();
 sg13g2_fill_2 FILLER_54_1735 ();
 sg13g2_decap_4 FILLER_54_1743 ();
 sg13g2_fill_1 FILLER_54_1747 ();
 sg13g2_fill_2 FILLER_54_1770 ();
 sg13g2_decap_8 FILLER_54_1781 ();
 sg13g2_decap_8 FILLER_54_1807 ();
 sg13g2_decap_8 FILLER_54_1814 ();
 sg13g2_fill_1 FILLER_54_1821 ();
 sg13g2_decap_8 FILLER_54_1827 ();
 sg13g2_fill_2 FILLER_54_1834 ();
 sg13g2_fill_1 FILLER_54_1836 ();
 sg13g2_fill_2 FILLER_54_1842 ();
 sg13g2_fill_1 FILLER_54_1844 ();
 sg13g2_fill_2 FILLER_54_1879 ();
 sg13g2_fill_1 FILLER_54_1881 ();
 sg13g2_decap_8 FILLER_54_1888 ();
 sg13g2_decap_8 FILLER_54_1911 ();
 sg13g2_decap_8 FILLER_54_1918 ();
 sg13g2_fill_1 FILLER_54_1925 ();
 sg13g2_decap_8 FILLER_54_1935 ();
 sg13g2_fill_1 FILLER_54_1942 ();
 sg13g2_decap_8 FILLER_54_1952 ();
 sg13g2_fill_2 FILLER_54_1959 ();
 sg13g2_decap_8 FILLER_54_1966 ();
 sg13g2_decap_4 FILLER_54_1973 ();
 sg13g2_fill_1 FILLER_54_1977 ();
 sg13g2_decap_8 FILLER_54_1991 ();
 sg13g2_fill_2 FILLER_54_1998 ();
 sg13g2_fill_1 FILLER_54_2000 ();
 sg13g2_fill_1 FILLER_54_2019 ();
 sg13g2_fill_2 FILLER_54_2033 ();
 sg13g2_fill_2 FILLER_54_2040 ();
 sg13g2_fill_1 FILLER_54_2042 ();
 sg13g2_decap_8 FILLER_54_2051 ();
 sg13g2_decap_4 FILLER_54_2058 ();
 sg13g2_fill_1 FILLER_54_2062 ();
 sg13g2_fill_2 FILLER_54_2105 ();
 sg13g2_fill_2 FILLER_54_2117 ();
 sg13g2_fill_1 FILLER_54_2119 ();
 sg13g2_fill_2 FILLER_54_2125 ();
 sg13g2_fill_1 FILLER_54_2127 ();
 sg13g2_fill_2 FILLER_54_2140 ();
 sg13g2_decap_4 FILLER_54_2156 ();
 sg13g2_fill_1 FILLER_54_2160 ();
 sg13g2_fill_2 FILLER_54_2169 ();
 sg13g2_fill_1 FILLER_54_2171 ();
 sg13g2_decap_8 FILLER_54_2180 ();
 sg13g2_fill_2 FILLER_54_2187 ();
 sg13g2_decap_4 FILLER_54_2213 ();
 sg13g2_fill_1 FILLER_54_2217 ();
 sg13g2_fill_2 FILLER_54_2244 ();
 sg13g2_fill_1 FILLER_54_2246 ();
 sg13g2_decap_8 FILLER_54_2267 ();
 sg13g2_decap_4 FILLER_54_2274 ();
 sg13g2_decap_4 FILLER_54_2297 ();
 sg13g2_decap_4 FILLER_54_2314 ();
 sg13g2_decap_4 FILLER_54_2322 ();
 sg13g2_fill_2 FILLER_54_2326 ();
 sg13g2_decap_4 FILLER_54_2377 ();
 sg13g2_fill_2 FILLER_54_2381 ();
 sg13g2_fill_2 FILLER_54_2393 ();
 sg13g2_decap_8 FILLER_54_2403 ();
 sg13g2_decap_4 FILLER_54_2410 ();
 sg13g2_fill_1 FILLER_54_2414 ();
 sg13g2_fill_2 FILLER_54_2436 ();
 sg13g2_fill_1 FILLER_54_2438 ();
 sg13g2_decap_4 FILLER_54_2471 ();
 sg13g2_decap_4 FILLER_54_2479 ();
 sg13g2_fill_2 FILLER_54_2489 ();
 sg13g2_fill_1 FILLER_54_2505 ();
 sg13g2_fill_2 FILLER_54_2543 ();
 sg13g2_fill_1 FILLER_54_2545 ();
 sg13g2_fill_2 FILLER_54_2557 ();
 sg13g2_fill_1 FILLER_54_2559 ();
 sg13g2_decap_4 FILLER_54_2582 ();
 sg13g2_fill_1 FILLER_54_2586 ();
 sg13g2_decap_8 FILLER_54_2591 ();
 sg13g2_decap_8 FILLER_54_2598 ();
 sg13g2_decap_8 FILLER_54_2605 ();
 sg13g2_fill_1 FILLER_54_2612 ();
 sg13g2_decap_8 FILLER_54_2642 ();
 sg13g2_decap_8 FILLER_54_2649 ();
 sg13g2_fill_2 FILLER_54_2656 ();
 sg13g2_fill_1 FILLER_54_2676 ();
 sg13g2_fill_2 FILLER_54_2681 ();
 sg13g2_fill_1 FILLER_54_2683 ();
 sg13g2_fill_2 FILLER_54_2714 ();
 sg13g2_fill_1 FILLER_54_2716 ();
 sg13g2_fill_1 FILLER_54_2732 ();
 sg13g2_decap_8 FILLER_54_2741 ();
 sg13g2_fill_1 FILLER_54_2753 ();
 sg13g2_decap_8 FILLER_54_2763 ();
 sg13g2_decap_8 FILLER_54_2770 ();
 sg13g2_fill_2 FILLER_54_2782 ();
 sg13g2_fill_1 FILLER_54_2784 ();
 sg13g2_fill_2 FILLER_54_2790 ();
 sg13g2_fill_1 FILLER_54_2800 ();
 sg13g2_decap_8 FILLER_54_2805 ();
 sg13g2_fill_2 FILLER_54_2812 ();
 sg13g2_fill_1 FILLER_54_2822 ();
 sg13g2_fill_2 FILLER_54_2866 ();
 sg13g2_fill_1 FILLER_54_2868 ();
 sg13g2_fill_2 FILLER_54_2891 ();
 sg13g2_fill_1 FILLER_54_2893 ();
 sg13g2_fill_2 FILLER_54_2898 ();
 sg13g2_fill_1 FILLER_54_2900 ();
 sg13g2_decap_8 FILLER_54_2905 ();
 sg13g2_fill_2 FILLER_54_2912 ();
 sg13g2_fill_2 FILLER_54_2918 ();
 sg13g2_fill_2 FILLER_54_2928 ();
 sg13g2_fill_1 FILLER_54_2930 ();
 sg13g2_decap_8 FILLER_54_2935 ();
 sg13g2_decap_8 FILLER_54_2942 ();
 sg13g2_decap_4 FILLER_54_2949 ();
 sg13g2_decap_4 FILLER_54_2969 ();
 sg13g2_fill_2 FILLER_54_2973 ();
 sg13g2_decap_8 FILLER_54_2988 ();
 sg13g2_decap_8 FILLER_54_2995 ();
 sg13g2_decap_8 FILLER_54_3002 ();
 sg13g2_decap_8 FILLER_54_3013 ();
 sg13g2_decap_8 FILLER_54_3020 ();
 sg13g2_decap_4 FILLER_54_3027 ();
 sg13g2_decap_8 FILLER_54_3057 ();
 sg13g2_decap_8 FILLER_54_3064 ();
 sg13g2_decap_8 FILLER_54_3071 ();
 sg13g2_decap_8 FILLER_54_3078 ();
 sg13g2_decap_8 FILLER_54_3085 ();
 sg13g2_decap_8 FILLER_54_3092 ();
 sg13g2_decap_8 FILLER_54_3099 ();
 sg13g2_decap_8 FILLER_54_3106 ();
 sg13g2_decap_8 FILLER_54_3113 ();
 sg13g2_decap_8 FILLER_54_3120 ();
 sg13g2_decap_8 FILLER_54_3127 ();
 sg13g2_decap_8 FILLER_54_3134 ();
 sg13g2_decap_8 FILLER_54_3141 ();
 sg13g2_decap_8 FILLER_54_3148 ();
 sg13g2_decap_8 FILLER_54_3155 ();
 sg13g2_decap_8 FILLER_54_3162 ();
 sg13g2_decap_8 FILLER_54_3169 ();
 sg13g2_decap_8 FILLER_54_3176 ();
 sg13g2_decap_8 FILLER_54_3183 ();
 sg13g2_decap_8 FILLER_54_3190 ();
 sg13g2_decap_8 FILLER_54_3197 ();
 sg13g2_decap_8 FILLER_54_3204 ();
 sg13g2_decap_8 FILLER_54_3211 ();
 sg13g2_decap_8 FILLER_54_3218 ();
 sg13g2_decap_8 FILLER_54_3225 ();
 sg13g2_decap_8 FILLER_54_3232 ();
 sg13g2_decap_8 FILLER_54_3239 ();
 sg13g2_decap_8 FILLER_54_3246 ();
 sg13g2_decap_8 FILLER_54_3253 ();
 sg13g2_decap_8 FILLER_54_3260 ();
 sg13g2_decap_8 FILLER_54_3267 ();
 sg13g2_decap_8 FILLER_54_3274 ();
 sg13g2_decap_8 FILLER_54_3281 ();
 sg13g2_decap_8 FILLER_54_3288 ();
 sg13g2_decap_8 FILLER_54_3295 ();
 sg13g2_decap_8 FILLER_54_3302 ();
 sg13g2_decap_8 FILLER_54_3309 ();
 sg13g2_decap_8 FILLER_54_3316 ();
 sg13g2_decap_8 FILLER_54_3323 ();
 sg13g2_decap_8 FILLER_54_3330 ();
 sg13g2_decap_8 FILLER_54_3337 ();
 sg13g2_decap_8 FILLER_54_3344 ();
 sg13g2_decap_8 FILLER_54_3351 ();
 sg13g2_decap_8 FILLER_54_3358 ();
 sg13g2_decap_8 FILLER_54_3365 ();
 sg13g2_decap_8 FILLER_54_3372 ();
 sg13g2_decap_8 FILLER_54_3379 ();
 sg13g2_decap_8 FILLER_54_3386 ();
 sg13g2_decap_8 FILLER_54_3393 ();
 sg13g2_decap_8 FILLER_54_3400 ();
 sg13g2_decap_8 FILLER_54_3407 ();
 sg13g2_decap_8 FILLER_54_3414 ();
 sg13g2_decap_8 FILLER_54_3421 ();
 sg13g2_decap_8 FILLER_54_3428 ();
 sg13g2_decap_8 FILLER_54_3435 ();
 sg13g2_decap_8 FILLER_54_3442 ();
 sg13g2_decap_8 FILLER_54_3449 ();
 sg13g2_decap_8 FILLER_54_3456 ();
 sg13g2_decap_8 FILLER_54_3463 ();
 sg13g2_decap_8 FILLER_54_3470 ();
 sg13g2_decap_8 FILLER_54_3477 ();
 sg13g2_decap_8 FILLER_54_3484 ();
 sg13g2_decap_8 FILLER_54_3491 ();
 sg13g2_decap_8 FILLER_54_3498 ();
 sg13g2_decap_8 FILLER_54_3505 ();
 sg13g2_decap_8 FILLER_54_3512 ();
 sg13g2_decap_8 FILLER_54_3519 ();
 sg13g2_decap_8 FILLER_54_3526 ();
 sg13g2_decap_8 FILLER_54_3533 ();
 sg13g2_decap_8 FILLER_54_3540 ();
 sg13g2_decap_8 FILLER_54_3547 ();
 sg13g2_decap_8 FILLER_54_3554 ();
 sg13g2_decap_8 FILLER_54_3561 ();
 sg13g2_decap_8 FILLER_54_3568 ();
 sg13g2_decap_4 FILLER_54_3575 ();
 sg13g2_fill_1 FILLER_54_3579 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_fill_2 FILLER_55_7 ();
 sg13g2_fill_1 FILLER_55_9 ();
 sg13g2_decap_4 FILLER_55_56 ();
 sg13g2_fill_2 FILLER_55_80 ();
 sg13g2_fill_1 FILLER_55_82 ();
 sg13g2_fill_1 FILLER_55_117 ();
 sg13g2_decap_8 FILLER_55_138 ();
 sg13g2_fill_2 FILLER_55_145 ();
 sg13g2_decap_4 FILLER_55_156 ();
 sg13g2_decap_4 FILLER_55_212 ();
 sg13g2_fill_2 FILLER_55_225 ();
 sg13g2_fill_1 FILLER_55_227 ();
 sg13g2_fill_2 FILLER_55_255 ();
 sg13g2_fill_2 FILLER_55_286 ();
 sg13g2_fill_1 FILLER_55_288 ();
 sg13g2_fill_2 FILLER_55_300 ();
 sg13g2_fill_1 FILLER_55_328 ();
 sg13g2_fill_2 FILLER_55_355 ();
 sg13g2_fill_2 FILLER_55_361 ();
 sg13g2_fill_1 FILLER_55_363 ();
 sg13g2_decap_8 FILLER_55_368 ();
 sg13g2_fill_2 FILLER_55_375 ();
 sg13g2_fill_1 FILLER_55_377 ();
 sg13g2_fill_2 FILLER_55_404 ();
 sg13g2_fill_1 FILLER_55_406 ();
 sg13g2_fill_2 FILLER_55_421 ();
 sg13g2_fill_1 FILLER_55_423 ();
 sg13g2_fill_2 FILLER_55_463 ();
 sg13g2_fill_2 FILLER_55_494 ();
 sg13g2_decap_4 FILLER_55_511 ();
 sg13g2_decap_8 FILLER_55_520 ();
 sg13g2_fill_2 FILLER_55_527 ();
 sg13g2_fill_1 FILLER_55_537 ();
 sg13g2_decap_8 FILLER_55_543 ();
 sg13g2_fill_1 FILLER_55_550 ();
 sg13g2_decap_4 FILLER_55_619 ();
 sg13g2_fill_2 FILLER_55_635 ();
 sg13g2_fill_1 FILLER_55_637 ();
 sg13g2_fill_2 FILLER_55_649 ();
 sg13g2_decap_8 FILLER_55_664 ();
 sg13g2_decap_4 FILLER_55_671 ();
 sg13g2_fill_2 FILLER_55_675 ();
 sg13g2_fill_2 FILLER_55_682 ();
 sg13g2_decap_4 FILLER_55_688 ();
 sg13g2_fill_1 FILLER_55_692 ();
 sg13g2_fill_1 FILLER_55_697 ();
 sg13g2_fill_2 FILLER_55_703 ();
 sg13g2_fill_1 FILLER_55_710 ();
 sg13g2_decap_8 FILLER_55_715 ();
 sg13g2_decap_8 FILLER_55_722 ();
 sg13g2_decap_4 FILLER_55_729 ();
 sg13g2_fill_2 FILLER_55_733 ();
 sg13g2_fill_2 FILLER_55_747 ();
 sg13g2_fill_1 FILLER_55_749 ();
 sg13g2_fill_2 FILLER_55_807 ();
 sg13g2_fill_1 FILLER_55_809 ();
 sg13g2_fill_1 FILLER_55_819 ();
 sg13g2_fill_1 FILLER_55_867 ();
 sg13g2_decap_4 FILLER_55_877 ();
 sg13g2_decap_4 FILLER_55_885 ();
 sg13g2_fill_2 FILLER_55_905 ();
 sg13g2_decap_4 FILLER_55_925 ();
 sg13g2_fill_1 FILLER_55_929 ();
 sg13g2_decap_4 FILLER_55_943 ();
 sg13g2_fill_2 FILLER_55_998 ();
 sg13g2_fill_2 FILLER_55_1010 ();
 sg13g2_fill_1 FILLER_55_1012 ();
 sg13g2_fill_2 FILLER_55_1022 ();
 sg13g2_fill_1 FILLER_55_1024 ();
 sg13g2_decap_4 FILLER_55_1051 ();
 sg13g2_fill_1 FILLER_55_1055 ();
 sg13g2_fill_1 FILLER_55_1064 ();
 sg13g2_fill_1 FILLER_55_1082 ();
 sg13g2_decap_8 FILLER_55_1096 ();
 sg13g2_fill_1 FILLER_55_1103 ();
 sg13g2_decap_8 FILLER_55_1108 ();
 sg13g2_fill_2 FILLER_55_1115 ();
 sg13g2_fill_2 FILLER_55_1123 ();
 sg13g2_fill_1 FILLER_55_1125 ();
 sg13g2_decap_8 FILLER_55_1130 ();
 sg13g2_decap_8 FILLER_55_1137 ();
 sg13g2_fill_1 FILLER_55_1144 ();
 sg13g2_decap_8 FILLER_55_1164 ();
 sg13g2_decap_8 FILLER_55_1174 ();
 sg13g2_decap_8 FILLER_55_1181 ();
 sg13g2_decap_8 FILLER_55_1188 ();
 sg13g2_fill_2 FILLER_55_1195 ();
 sg13g2_fill_2 FILLER_55_1223 ();
 sg13g2_decap_4 FILLER_55_1234 ();
 sg13g2_decap_4 FILLER_55_1243 ();
 sg13g2_fill_2 FILLER_55_1261 ();
 sg13g2_fill_1 FILLER_55_1263 ();
 sg13g2_fill_1 FILLER_55_1275 ();
 sg13g2_decap_8 FILLER_55_1289 ();
 sg13g2_fill_2 FILLER_55_1296 ();
 sg13g2_fill_1 FILLER_55_1298 ();
 sg13g2_decap_4 FILLER_55_1303 ();
 sg13g2_fill_1 FILLER_55_1307 ();
 sg13g2_decap_8 FILLER_55_1348 ();
 sg13g2_fill_1 FILLER_55_1456 ();
 sg13g2_fill_2 FILLER_55_1465 ();
 sg13g2_fill_1 FILLER_55_1467 ();
 sg13g2_decap_8 FILLER_55_1473 ();
 sg13g2_fill_2 FILLER_55_1480 ();
 sg13g2_fill_1 FILLER_55_1482 ();
 sg13g2_fill_1 FILLER_55_1492 ();
 sg13g2_decap_8 FILLER_55_1514 ();
 sg13g2_fill_1 FILLER_55_1521 ();
 sg13g2_fill_1 FILLER_55_1532 ();
 sg13g2_fill_2 FILLER_55_1543 ();
 sg13g2_fill_2 FILLER_55_1550 ();
 sg13g2_fill_2 FILLER_55_1560 ();
 sg13g2_fill_1 FILLER_55_1562 ();
 sg13g2_fill_2 FILLER_55_1581 ();
 sg13g2_decap_4 FILLER_55_1587 ();
 sg13g2_fill_1 FILLER_55_1591 ();
 sg13g2_fill_2 FILLER_55_1597 ();
 sg13g2_fill_1 FILLER_55_1599 ();
 sg13g2_fill_1 FILLER_55_1613 ();
 sg13g2_fill_1 FILLER_55_1632 ();
 sg13g2_decap_4 FILLER_55_1642 ();
 sg13g2_fill_1 FILLER_55_1646 ();
 sg13g2_decap_8 FILLER_55_1656 ();
 sg13g2_fill_1 FILLER_55_1668 ();
 sg13g2_decap_4 FILLER_55_1674 ();
 sg13g2_decap_4 FILLER_55_1683 ();
 sg13g2_fill_1 FILLER_55_1707 ();
 sg13g2_decap_8 FILLER_55_1718 ();
 sg13g2_fill_2 FILLER_55_1725 ();
 sg13g2_decap_4 FILLER_55_1751 ();
 sg13g2_fill_1 FILLER_55_1755 ();
 sg13g2_fill_2 FILLER_55_1761 ();
 sg13g2_fill_1 FILLER_55_1763 ();
 sg13g2_fill_1 FILLER_55_1770 ();
 sg13g2_fill_2 FILLER_55_1779 ();
 sg13g2_fill_1 FILLER_55_1781 ();
 sg13g2_fill_1 FILLER_55_1802 ();
 sg13g2_decap_8 FILLER_55_1811 ();
 sg13g2_decap_4 FILLER_55_1818 ();
 sg13g2_fill_1 FILLER_55_1822 ();
 sg13g2_fill_2 FILLER_55_1834 ();
 sg13g2_fill_1 FILLER_55_1877 ();
 sg13g2_decap_8 FILLER_55_1886 ();
 sg13g2_fill_2 FILLER_55_1893 ();
 sg13g2_fill_1 FILLER_55_1914 ();
 sg13g2_decap_4 FILLER_55_1928 ();
 sg13g2_fill_2 FILLER_55_1973 ();
 sg13g2_fill_1 FILLER_55_1975 ();
 sg13g2_fill_1 FILLER_55_1989 ();
 sg13g2_decap_8 FILLER_55_1998 ();
 sg13g2_fill_2 FILLER_55_2005 ();
 sg13g2_decap_8 FILLER_55_2015 ();
 sg13g2_fill_2 FILLER_55_2032 ();
 sg13g2_decap_4 FILLER_55_2039 ();
 sg13g2_fill_2 FILLER_55_2043 ();
 sg13g2_decap_4 FILLER_55_2050 ();
 sg13g2_fill_2 FILLER_55_2054 ();
 sg13g2_decap_8 FILLER_55_2074 ();
 sg13g2_decap_8 FILLER_55_2086 ();
 sg13g2_decap_8 FILLER_55_2093 ();
 sg13g2_decap_4 FILLER_55_2100 ();
 sg13g2_fill_2 FILLER_55_2104 ();
 sg13g2_fill_2 FILLER_55_2111 ();
 sg13g2_fill_1 FILLER_55_2113 ();
 sg13g2_fill_1 FILLER_55_2130 ();
 sg13g2_fill_2 FILLER_55_2135 ();
 sg13g2_fill_2 FILLER_55_2142 ();
 sg13g2_decap_4 FILLER_55_2157 ();
 sg13g2_fill_2 FILLER_55_2161 ();
 sg13g2_decap_8 FILLER_55_2182 ();
 sg13g2_fill_2 FILLER_55_2189 ();
 sg13g2_fill_2 FILLER_55_2195 ();
 sg13g2_fill_1 FILLER_55_2197 ();
 sg13g2_fill_1 FILLER_55_2202 ();
 sg13g2_decap_8 FILLER_55_2208 ();
 sg13g2_decap_4 FILLER_55_2215 ();
 sg13g2_fill_1 FILLER_55_2219 ();
 sg13g2_decap_4 FILLER_55_2235 ();
 sg13g2_decap_8 FILLER_55_2244 ();
 sg13g2_decap_4 FILLER_55_2251 ();
 sg13g2_fill_1 FILLER_55_2255 ();
 sg13g2_fill_1 FILLER_55_2271 ();
 sg13g2_decap_8 FILLER_55_2276 ();
 sg13g2_decap_8 FILLER_55_2283 ();
 sg13g2_decap_8 FILLER_55_2290 ();
 sg13g2_decap_4 FILLER_55_2305 ();
 sg13g2_fill_2 FILLER_55_2331 ();
 sg13g2_decap_8 FILLER_55_2342 ();
 sg13g2_decap_4 FILLER_55_2349 ();
 sg13g2_fill_1 FILLER_55_2353 ();
 sg13g2_decap_8 FILLER_55_2368 ();
 sg13g2_decap_4 FILLER_55_2375 ();
 sg13g2_fill_2 FILLER_55_2391 ();
 sg13g2_fill_1 FILLER_55_2393 ();
 sg13g2_fill_1 FILLER_55_2402 ();
 sg13g2_decap_8 FILLER_55_2437 ();
 sg13g2_fill_1 FILLER_55_2444 ();
 sg13g2_decap_4 FILLER_55_2491 ();
 sg13g2_fill_2 FILLER_55_2515 ();
 sg13g2_fill_2 FILLER_55_2521 ();
 sg13g2_fill_1 FILLER_55_2523 ();
 sg13g2_fill_1 FILLER_55_2544 ();
 sg13g2_decap_8 FILLER_55_2618 ();
 sg13g2_decap_8 FILLER_55_2625 ();
 sg13g2_fill_1 FILLER_55_2637 ();
 sg13g2_decap_8 FILLER_55_2643 ();
 sg13g2_decap_8 FILLER_55_2664 ();
 sg13g2_decap_4 FILLER_55_2687 ();
 sg13g2_fill_2 FILLER_55_2691 ();
 sg13g2_decap_4 FILLER_55_2697 ();
 sg13g2_decap_8 FILLER_55_2705 ();
 sg13g2_decap_4 FILLER_55_2712 ();
 sg13g2_fill_1 FILLER_55_2716 ();
 sg13g2_decap_8 FILLER_55_2729 ();
 sg13g2_fill_2 FILLER_55_2736 ();
 sg13g2_fill_2 FILLER_55_2751 ();
 sg13g2_fill_1 FILLER_55_2753 ();
 sg13g2_fill_2 FILLER_55_2762 ();
 sg13g2_fill_1 FILLER_55_2764 ();
 sg13g2_fill_1 FILLER_55_2770 ();
 sg13g2_decap_8 FILLER_55_2775 ();
 sg13g2_fill_2 FILLER_55_2782 ();
 sg13g2_fill_1 FILLER_55_2784 ();
 sg13g2_fill_2 FILLER_55_2801 ();
 sg13g2_fill_2 FILLER_55_2807 ();
 sg13g2_fill_1 FILLER_55_2809 ();
 sg13g2_fill_2 FILLER_55_2827 ();
 sg13g2_fill_1 FILLER_55_2833 ();
 sg13g2_decap_8 FILLER_55_2838 ();
 sg13g2_decap_8 FILLER_55_2845 ();
 sg13g2_fill_2 FILLER_55_2852 ();
 sg13g2_fill_1 FILLER_55_2854 ();
 sg13g2_decap_8 FILLER_55_2879 ();
 sg13g2_decap_4 FILLER_55_2886 ();
 sg13g2_decap_4 FILLER_55_2902 ();
 sg13g2_fill_2 FILLER_55_2915 ();
 sg13g2_fill_1 FILLER_55_2947 ();
 sg13g2_fill_1 FILLER_55_2970 ();
 sg13g2_decap_8 FILLER_55_2997 ();
 sg13g2_decap_8 FILLER_55_3004 ();
 sg13g2_decap_8 FILLER_55_3011 ();
 sg13g2_decap_8 FILLER_55_3018 ();
 sg13g2_decap_8 FILLER_55_3025 ();
 sg13g2_decap_8 FILLER_55_3032 ();
 sg13g2_decap_8 FILLER_55_3039 ();
 sg13g2_decap_8 FILLER_55_3046 ();
 sg13g2_decap_8 FILLER_55_3053 ();
 sg13g2_decap_8 FILLER_55_3060 ();
 sg13g2_decap_8 FILLER_55_3067 ();
 sg13g2_decap_8 FILLER_55_3074 ();
 sg13g2_decap_8 FILLER_55_3081 ();
 sg13g2_decap_8 FILLER_55_3088 ();
 sg13g2_decap_8 FILLER_55_3095 ();
 sg13g2_decap_8 FILLER_55_3102 ();
 sg13g2_decap_8 FILLER_55_3109 ();
 sg13g2_decap_8 FILLER_55_3116 ();
 sg13g2_decap_8 FILLER_55_3123 ();
 sg13g2_decap_8 FILLER_55_3130 ();
 sg13g2_decap_8 FILLER_55_3137 ();
 sg13g2_decap_8 FILLER_55_3144 ();
 sg13g2_decap_8 FILLER_55_3151 ();
 sg13g2_decap_8 FILLER_55_3158 ();
 sg13g2_decap_8 FILLER_55_3165 ();
 sg13g2_decap_8 FILLER_55_3172 ();
 sg13g2_decap_8 FILLER_55_3179 ();
 sg13g2_decap_8 FILLER_55_3186 ();
 sg13g2_decap_8 FILLER_55_3193 ();
 sg13g2_decap_8 FILLER_55_3200 ();
 sg13g2_decap_8 FILLER_55_3207 ();
 sg13g2_decap_8 FILLER_55_3214 ();
 sg13g2_decap_8 FILLER_55_3221 ();
 sg13g2_decap_8 FILLER_55_3228 ();
 sg13g2_decap_8 FILLER_55_3235 ();
 sg13g2_decap_8 FILLER_55_3242 ();
 sg13g2_decap_8 FILLER_55_3249 ();
 sg13g2_decap_8 FILLER_55_3256 ();
 sg13g2_decap_8 FILLER_55_3263 ();
 sg13g2_decap_8 FILLER_55_3270 ();
 sg13g2_decap_8 FILLER_55_3277 ();
 sg13g2_decap_8 FILLER_55_3284 ();
 sg13g2_decap_8 FILLER_55_3291 ();
 sg13g2_decap_8 FILLER_55_3298 ();
 sg13g2_decap_8 FILLER_55_3305 ();
 sg13g2_decap_8 FILLER_55_3312 ();
 sg13g2_decap_8 FILLER_55_3319 ();
 sg13g2_decap_8 FILLER_55_3326 ();
 sg13g2_decap_8 FILLER_55_3333 ();
 sg13g2_decap_8 FILLER_55_3340 ();
 sg13g2_decap_8 FILLER_55_3347 ();
 sg13g2_decap_8 FILLER_55_3354 ();
 sg13g2_decap_8 FILLER_55_3361 ();
 sg13g2_decap_8 FILLER_55_3368 ();
 sg13g2_decap_8 FILLER_55_3375 ();
 sg13g2_decap_8 FILLER_55_3382 ();
 sg13g2_decap_8 FILLER_55_3389 ();
 sg13g2_decap_8 FILLER_55_3396 ();
 sg13g2_decap_8 FILLER_55_3403 ();
 sg13g2_decap_8 FILLER_55_3410 ();
 sg13g2_decap_8 FILLER_55_3417 ();
 sg13g2_decap_8 FILLER_55_3424 ();
 sg13g2_decap_8 FILLER_55_3431 ();
 sg13g2_decap_8 FILLER_55_3438 ();
 sg13g2_decap_8 FILLER_55_3445 ();
 sg13g2_decap_8 FILLER_55_3452 ();
 sg13g2_decap_8 FILLER_55_3459 ();
 sg13g2_decap_8 FILLER_55_3466 ();
 sg13g2_decap_8 FILLER_55_3473 ();
 sg13g2_decap_8 FILLER_55_3480 ();
 sg13g2_decap_8 FILLER_55_3487 ();
 sg13g2_decap_8 FILLER_55_3494 ();
 sg13g2_decap_8 FILLER_55_3501 ();
 sg13g2_decap_8 FILLER_55_3508 ();
 sg13g2_decap_8 FILLER_55_3515 ();
 sg13g2_decap_8 FILLER_55_3522 ();
 sg13g2_decap_8 FILLER_55_3529 ();
 sg13g2_decap_8 FILLER_55_3536 ();
 sg13g2_decap_8 FILLER_55_3543 ();
 sg13g2_decap_8 FILLER_55_3550 ();
 sg13g2_decap_8 FILLER_55_3557 ();
 sg13g2_decap_8 FILLER_55_3564 ();
 sg13g2_decap_8 FILLER_55_3571 ();
 sg13g2_fill_2 FILLER_55_3578 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_33 ();
 sg13g2_fill_2 FILLER_56_48 ();
 sg13g2_fill_1 FILLER_56_58 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_fill_1 FILLER_56_91 ();
 sg13g2_decap_8 FILLER_56_111 ();
 sg13g2_decap_4 FILLER_56_118 ();
 sg13g2_decap_8 FILLER_56_130 ();
 sg13g2_decap_4 FILLER_56_137 ();
 sg13g2_fill_1 FILLER_56_141 ();
 sg13g2_decap_4 FILLER_56_168 ();
 sg13g2_fill_1 FILLER_56_187 ();
 sg13g2_fill_2 FILLER_56_202 ();
 sg13g2_decap_8 FILLER_56_217 ();
 sg13g2_fill_1 FILLER_56_224 ();
 sg13g2_fill_2 FILLER_56_251 ();
 sg13g2_fill_1 FILLER_56_262 ();
 sg13g2_fill_2 FILLER_56_279 ();
 sg13g2_fill_2 FILLER_56_296 ();
 sg13g2_decap_8 FILLER_56_325 ();
 sg13g2_decap_4 FILLER_56_332 ();
 sg13g2_fill_1 FILLER_56_351 ();
 sg13g2_decap_4 FILLER_56_381 ();
 sg13g2_decap_4 FILLER_56_395 ();
 sg13g2_decap_8 FILLER_56_434 ();
 sg13g2_decap_4 FILLER_56_441 ();
 sg13g2_fill_1 FILLER_56_445 ();
 sg13g2_fill_2 FILLER_56_469 ();
 sg13g2_fill_1 FILLER_56_476 ();
 sg13g2_fill_2 FILLER_56_506 ();
 sg13g2_fill_1 FILLER_56_508 ();
 sg13g2_decap_8 FILLER_56_517 ();
 sg13g2_decap_4 FILLER_56_550 ();
 sg13g2_decap_8 FILLER_56_559 ();
 sg13g2_decap_4 FILLER_56_566 ();
 sg13g2_fill_2 FILLER_56_570 ();
 sg13g2_decap_8 FILLER_56_576 ();
 sg13g2_decap_4 FILLER_56_583 ();
 sg13g2_fill_2 FILLER_56_587 ();
 sg13g2_decap_4 FILLER_56_598 ();
 sg13g2_decap_4 FILLER_56_605 ();
 sg13g2_decap_8 FILLER_56_631 ();
 sg13g2_fill_2 FILLER_56_638 ();
 sg13g2_fill_1 FILLER_56_640 ();
 sg13g2_fill_1 FILLER_56_644 ();
 sg13g2_fill_2 FILLER_56_659 ();
 sg13g2_decap_4 FILLER_56_667 ();
 sg13g2_fill_1 FILLER_56_671 ();
 sg13g2_fill_2 FILLER_56_694 ();
 sg13g2_fill_1 FILLER_56_711 ();
 sg13g2_fill_2 FILLER_56_764 ();
 sg13g2_fill_1 FILLER_56_766 ();
 sg13g2_decap_8 FILLER_56_776 ();
 sg13g2_decap_8 FILLER_56_783 ();
 sg13g2_decap_8 FILLER_56_790 ();
 sg13g2_decap_4 FILLER_56_797 ();
 sg13g2_fill_2 FILLER_56_829 ();
 sg13g2_fill_1 FILLER_56_836 ();
 sg13g2_fill_2 FILLER_56_852 ();
 sg13g2_fill_2 FILLER_56_870 ();
 sg13g2_decap_8 FILLER_56_877 ();
 sg13g2_decap_8 FILLER_56_924 ();
 sg13g2_decap_8 FILLER_56_950 ();
 sg13g2_fill_1 FILLER_56_957 ();
 sg13g2_decap_4 FILLER_56_961 ();
 sg13g2_fill_2 FILLER_56_965 ();
 sg13g2_decap_8 FILLER_56_976 ();
 sg13g2_decap_8 FILLER_56_983 ();
 sg13g2_fill_2 FILLER_56_1057 ();
 sg13g2_fill_1 FILLER_56_1059 ();
 sg13g2_fill_2 FILLER_56_1101 ();
 sg13g2_fill_1 FILLER_56_1142 ();
 sg13g2_fill_2 FILLER_56_1199 ();
 sg13g2_fill_1 FILLER_56_1201 ();
 sg13g2_fill_2 FILLER_56_1214 ();
 sg13g2_fill_2 FILLER_56_1231 ();
 sg13g2_fill_1 FILLER_56_1242 ();
 sg13g2_decap_8 FILLER_56_1314 ();
 sg13g2_fill_1 FILLER_56_1321 ();
 sg13g2_decap_8 FILLER_56_1353 ();
 sg13g2_decap_8 FILLER_56_1360 ();
 sg13g2_decap_8 FILLER_56_1367 ();
 sg13g2_decap_8 FILLER_56_1378 ();
 sg13g2_decap_8 FILLER_56_1385 ();
 sg13g2_fill_1 FILLER_56_1392 ();
 sg13g2_decap_8 FILLER_56_1404 ();
 sg13g2_fill_2 FILLER_56_1411 ();
 sg13g2_fill_1 FILLER_56_1413 ();
 sg13g2_fill_2 FILLER_56_1418 ();
 sg13g2_decap_8 FILLER_56_1428 ();
 sg13g2_decap_4 FILLER_56_1435 ();
 sg13g2_fill_1 FILLER_56_1439 ();
 sg13g2_decap_8 FILLER_56_1446 ();
 sg13g2_decap_8 FILLER_56_1453 ();
 sg13g2_decap_4 FILLER_56_1460 ();
 sg13g2_fill_2 FILLER_56_1464 ();
 sg13g2_decap_8 FILLER_56_1481 ();
 sg13g2_decap_8 FILLER_56_1488 ();
 sg13g2_fill_2 FILLER_56_1495 ();
 sg13g2_decap_4 FILLER_56_1523 ();
 sg13g2_fill_1 FILLER_56_1527 ();
 sg13g2_decap_8 FILLER_56_1533 ();
 sg13g2_decap_8 FILLER_56_1540 ();
 sg13g2_decap_8 FILLER_56_1547 ();
 sg13g2_decap_8 FILLER_56_1554 ();
 sg13g2_fill_2 FILLER_56_1561 ();
 sg13g2_fill_1 FILLER_56_1563 ();
 sg13g2_fill_2 FILLER_56_1573 ();
 sg13g2_fill_2 FILLER_56_1580 ();
 sg13g2_decap_4 FILLER_56_1587 ();
 sg13g2_fill_2 FILLER_56_1591 ();
 sg13g2_decap_8 FILLER_56_1598 ();
 sg13g2_fill_2 FILLER_56_1605 ();
 sg13g2_fill_2 FILLER_56_1624 ();
 sg13g2_fill_1 FILLER_56_1626 ();
 sg13g2_fill_2 FILLER_56_1637 ();
 sg13g2_fill_1 FILLER_56_1639 ();
 sg13g2_fill_2 FILLER_56_1663 ();
 sg13g2_fill_1 FILLER_56_1665 ();
 sg13g2_fill_1 FILLER_56_1674 ();
 sg13g2_decap_4 FILLER_56_1683 ();
 sg13g2_fill_1 FILLER_56_1687 ();
 sg13g2_fill_2 FILLER_56_1712 ();
 sg13g2_fill_1 FILLER_56_1714 ();
 sg13g2_decap_4 FILLER_56_1726 ();
 sg13g2_decap_8 FILLER_56_1740 ();
 sg13g2_decap_8 FILLER_56_1747 ();
 sg13g2_decap_4 FILLER_56_1754 ();
 sg13g2_fill_2 FILLER_56_1758 ();
 sg13g2_decap_8 FILLER_56_1773 ();
 sg13g2_decap_4 FILLER_56_1780 ();
 sg13g2_fill_1 FILLER_56_1784 ();
 sg13g2_decap_8 FILLER_56_1802 ();
 sg13g2_decap_8 FILLER_56_1809 ();
 sg13g2_decap_8 FILLER_56_1816 ();
 sg13g2_decap_4 FILLER_56_1842 ();
 sg13g2_decap_8 FILLER_56_1880 ();
 sg13g2_fill_1 FILLER_56_1887 ();
 sg13g2_fill_2 FILLER_56_1902 ();
 sg13g2_fill_1 FILLER_56_1904 ();
 sg13g2_fill_1 FILLER_56_1918 ();
 sg13g2_fill_2 FILLER_56_1925 ();
 sg13g2_fill_1 FILLER_56_1927 ();
 sg13g2_decap_8 FILLER_56_1933 ();
 sg13g2_fill_1 FILLER_56_1940 ();
 sg13g2_fill_1 FILLER_56_1955 ();
 sg13g2_decap_8 FILLER_56_1966 ();
 sg13g2_decap_4 FILLER_56_1973 ();
 sg13g2_fill_2 FILLER_56_1993 ();
 sg13g2_fill_1 FILLER_56_1995 ();
 sg13g2_fill_1 FILLER_56_2001 ();
 sg13g2_fill_1 FILLER_56_2012 ();
 sg13g2_decap_8 FILLER_56_2021 ();
 sg13g2_decap_8 FILLER_56_2028 ();
 sg13g2_decap_4 FILLER_56_2035 ();
 sg13g2_fill_2 FILLER_56_2047 ();
 sg13g2_fill_2 FILLER_56_2070 ();
 sg13g2_decap_8 FILLER_56_2078 ();
 sg13g2_fill_1 FILLER_56_2085 ();
 sg13g2_decap_4 FILLER_56_2092 ();
 sg13g2_fill_1 FILLER_56_2096 ();
 sg13g2_fill_1 FILLER_56_2127 ();
 sg13g2_fill_1 FILLER_56_2142 ();
 sg13g2_decap_4 FILLER_56_2168 ();
 sg13g2_decap_8 FILLER_56_2176 ();
 sg13g2_decap_8 FILLER_56_2214 ();
 sg13g2_fill_2 FILLER_56_2221 ();
 sg13g2_fill_2 FILLER_56_2238 ();
 sg13g2_decap_8 FILLER_56_2251 ();
 sg13g2_fill_2 FILLER_56_2266 ();
 sg13g2_fill_1 FILLER_56_2268 ();
 sg13g2_decap_8 FILLER_56_2283 ();
 sg13g2_fill_2 FILLER_56_2290 ();
 sg13g2_decap_4 FILLER_56_2317 ();
 sg13g2_fill_2 FILLER_56_2329 ();
 sg13g2_decap_8 FILLER_56_2339 ();
 sg13g2_decap_4 FILLER_56_2346 ();
 sg13g2_decap_8 FILLER_56_2376 ();
 sg13g2_decap_8 FILLER_56_2383 ();
 sg13g2_decap_4 FILLER_56_2390 ();
 sg13g2_fill_1 FILLER_56_2394 ();
 sg13g2_fill_2 FILLER_56_2404 ();
 sg13g2_decap_8 FILLER_56_2411 ();
 sg13g2_decap_4 FILLER_56_2418 ();
 sg13g2_fill_1 FILLER_56_2422 ();
 sg13g2_decap_4 FILLER_56_2435 ();
 sg13g2_fill_2 FILLER_56_2439 ();
 sg13g2_fill_1 FILLER_56_2454 ();
 sg13g2_decap_8 FILLER_56_2470 ();
 sg13g2_decap_8 FILLER_56_2477 ();
 sg13g2_fill_2 FILLER_56_2484 ();
 sg13g2_fill_1 FILLER_56_2486 ();
 sg13g2_decap_4 FILLER_56_2491 ();
 sg13g2_fill_1 FILLER_56_2495 ();
 sg13g2_decap_4 FILLER_56_2505 ();
 sg13g2_fill_1 FILLER_56_2509 ();
 sg13g2_fill_2 FILLER_56_2524 ();
 sg13g2_decap_8 FILLER_56_2548 ();
 sg13g2_fill_1 FILLER_56_2555 ();
 sg13g2_decap_8 FILLER_56_2560 ();
 sg13g2_fill_2 FILLER_56_2567 ();
 sg13g2_fill_1 FILLER_56_2569 ();
 sg13g2_decap_8 FILLER_56_2574 ();
 sg13g2_decap_4 FILLER_56_2585 ();
 sg13g2_fill_1 FILLER_56_2589 ();
 sg13g2_fill_1 FILLER_56_2593 ();
 sg13g2_fill_2 FILLER_56_2603 ();
 sg13g2_fill_1 FILLER_56_2605 ();
 sg13g2_decap_8 FILLER_56_2614 ();
 sg13g2_fill_1 FILLER_56_2621 ();
 sg13g2_decap_8 FILLER_56_2660 ();
 sg13g2_fill_1 FILLER_56_2667 ();
 sg13g2_decap_8 FILLER_56_2672 ();
 sg13g2_decap_8 FILLER_56_2679 ();
 sg13g2_fill_2 FILLER_56_2686 ();
 sg13g2_fill_1 FILLER_56_2688 ();
 sg13g2_decap_8 FILLER_56_2709 ();
 sg13g2_decap_8 FILLER_56_2732 ();
 sg13g2_fill_2 FILLER_56_2739 ();
 sg13g2_decap_4 FILLER_56_2758 ();
 sg13g2_fill_1 FILLER_56_2762 ();
 sg13g2_decap_4 FILLER_56_2792 ();
 sg13g2_fill_1 FILLER_56_2796 ();
 sg13g2_decap_8 FILLER_56_2808 ();
 sg13g2_decap_4 FILLER_56_2815 ();
 sg13g2_fill_2 FILLER_56_2819 ();
 sg13g2_fill_2 FILLER_56_2848 ();
 sg13g2_fill_1 FILLER_56_2850 ();
 sg13g2_decap_8 FILLER_56_2877 ();
 sg13g2_decap_8 FILLER_56_2892 ();
 sg13g2_fill_2 FILLER_56_2899 ();
 sg13g2_fill_2 FILLER_56_2923 ();
 sg13g2_fill_1 FILLER_56_2925 ();
 sg13g2_decap_4 FILLER_56_2930 ();
 sg13g2_fill_1 FILLER_56_2934 ();
 sg13g2_decap_8 FILLER_56_2940 ();
 sg13g2_decap_4 FILLER_56_2947 ();
 sg13g2_fill_1 FILLER_56_2951 ();
 sg13g2_fill_1 FILLER_56_2970 ();
 sg13g2_fill_2 FILLER_56_2980 ();
 sg13g2_decap_8 FILLER_56_2986 ();
 sg13g2_decap_8 FILLER_56_2993 ();
 sg13g2_decap_8 FILLER_56_3000 ();
 sg13g2_decap_4 FILLER_56_3007 ();
 sg13g2_fill_2 FILLER_56_3011 ();
 sg13g2_decap_8 FILLER_56_3024 ();
 sg13g2_decap_8 FILLER_56_3031 ();
 sg13g2_decap_8 FILLER_56_3038 ();
 sg13g2_decap_8 FILLER_56_3045 ();
 sg13g2_decap_8 FILLER_56_3052 ();
 sg13g2_decap_8 FILLER_56_3059 ();
 sg13g2_decap_8 FILLER_56_3066 ();
 sg13g2_decap_8 FILLER_56_3073 ();
 sg13g2_decap_8 FILLER_56_3080 ();
 sg13g2_decap_8 FILLER_56_3087 ();
 sg13g2_decap_8 FILLER_56_3094 ();
 sg13g2_decap_8 FILLER_56_3101 ();
 sg13g2_decap_8 FILLER_56_3108 ();
 sg13g2_decap_8 FILLER_56_3115 ();
 sg13g2_decap_8 FILLER_56_3122 ();
 sg13g2_decap_8 FILLER_56_3129 ();
 sg13g2_decap_8 FILLER_56_3136 ();
 sg13g2_decap_8 FILLER_56_3143 ();
 sg13g2_decap_8 FILLER_56_3150 ();
 sg13g2_decap_8 FILLER_56_3157 ();
 sg13g2_decap_8 FILLER_56_3164 ();
 sg13g2_decap_8 FILLER_56_3171 ();
 sg13g2_decap_8 FILLER_56_3178 ();
 sg13g2_decap_8 FILLER_56_3185 ();
 sg13g2_decap_8 FILLER_56_3192 ();
 sg13g2_decap_8 FILLER_56_3199 ();
 sg13g2_decap_8 FILLER_56_3206 ();
 sg13g2_decap_8 FILLER_56_3213 ();
 sg13g2_decap_8 FILLER_56_3220 ();
 sg13g2_decap_8 FILLER_56_3227 ();
 sg13g2_decap_8 FILLER_56_3234 ();
 sg13g2_decap_8 FILLER_56_3241 ();
 sg13g2_decap_8 FILLER_56_3248 ();
 sg13g2_decap_8 FILLER_56_3255 ();
 sg13g2_decap_8 FILLER_56_3262 ();
 sg13g2_decap_8 FILLER_56_3269 ();
 sg13g2_decap_8 FILLER_56_3276 ();
 sg13g2_decap_8 FILLER_56_3283 ();
 sg13g2_decap_8 FILLER_56_3290 ();
 sg13g2_decap_8 FILLER_56_3297 ();
 sg13g2_decap_8 FILLER_56_3304 ();
 sg13g2_decap_8 FILLER_56_3311 ();
 sg13g2_decap_8 FILLER_56_3318 ();
 sg13g2_decap_8 FILLER_56_3325 ();
 sg13g2_decap_8 FILLER_56_3332 ();
 sg13g2_decap_8 FILLER_56_3339 ();
 sg13g2_decap_8 FILLER_56_3346 ();
 sg13g2_decap_8 FILLER_56_3353 ();
 sg13g2_decap_8 FILLER_56_3360 ();
 sg13g2_decap_8 FILLER_56_3367 ();
 sg13g2_decap_8 FILLER_56_3374 ();
 sg13g2_decap_8 FILLER_56_3381 ();
 sg13g2_decap_8 FILLER_56_3388 ();
 sg13g2_decap_8 FILLER_56_3395 ();
 sg13g2_decap_8 FILLER_56_3402 ();
 sg13g2_decap_8 FILLER_56_3409 ();
 sg13g2_decap_8 FILLER_56_3416 ();
 sg13g2_decap_8 FILLER_56_3423 ();
 sg13g2_decap_8 FILLER_56_3430 ();
 sg13g2_decap_8 FILLER_56_3437 ();
 sg13g2_decap_8 FILLER_56_3444 ();
 sg13g2_decap_8 FILLER_56_3451 ();
 sg13g2_decap_8 FILLER_56_3458 ();
 sg13g2_decap_8 FILLER_56_3465 ();
 sg13g2_decap_8 FILLER_56_3472 ();
 sg13g2_decap_8 FILLER_56_3479 ();
 sg13g2_decap_8 FILLER_56_3486 ();
 sg13g2_decap_8 FILLER_56_3493 ();
 sg13g2_decap_8 FILLER_56_3500 ();
 sg13g2_decap_8 FILLER_56_3507 ();
 sg13g2_decap_8 FILLER_56_3514 ();
 sg13g2_decap_8 FILLER_56_3521 ();
 sg13g2_decap_8 FILLER_56_3528 ();
 sg13g2_decap_8 FILLER_56_3535 ();
 sg13g2_decap_8 FILLER_56_3542 ();
 sg13g2_decap_8 FILLER_56_3549 ();
 sg13g2_decap_8 FILLER_56_3556 ();
 sg13g2_decap_8 FILLER_56_3563 ();
 sg13g2_decap_8 FILLER_56_3570 ();
 sg13g2_fill_2 FILLER_56_3577 ();
 sg13g2_fill_1 FILLER_56_3579 ();
 sg13g2_fill_2 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_2 ();
 sg13g2_fill_1 FILLER_57_29 ();
 sg13g2_decap_4 FILLER_57_58 ();
 sg13g2_fill_1 FILLER_57_72 ();
 sg13g2_decap_8 FILLER_57_78 ();
 sg13g2_decap_8 FILLER_57_85 ();
 sg13g2_decap_4 FILLER_57_92 ();
 sg13g2_fill_1 FILLER_57_114 ();
 sg13g2_decap_4 FILLER_57_125 ();
 sg13g2_fill_1 FILLER_57_129 ();
 sg13g2_fill_2 FILLER_57_136 ();
 sg13g2_fill_1 FILLER_57_151 ();
 sg13g2_fill_2 FILLER_57_156 ();
 sg13g2_fill_1 FILLER_57_158 ();
 sg13g2_decap_8 FILLER_57_223 ();
 sg13g2_fill_2 FILLER_57_230 ();
 sg13g2_decap_4 FILLER_57_237 ();
 sg13g2_fill_2 FILLER_57_256 ();
 sg13g2_fill_1 FILLER_57_263 ();
 sg13g2_decap_8 FILLER_57_269 ();
 sg13g2_decap_8 FILLER_57_276 ();
 sg13g2_fill_1 FILLER_57_283 ();
 sg13g2_fill_2 FILLER_57_320 ();
 sg13g2_fill_1 FILLER_57_322 ();
 sg13g2_decap_4 FILLER_57_328 ();
 sg13g2_fill_2 FILLER_57_332 ();
 sg13g2_fill_1 FILLER_57_348 ();
 sg13g2_fill_2 FILLER_57_359 ();
 sg13g2_fill_2 FILLER_57_365 ();
 sg13g2_decap_8 FILLER_57_397 ();
 sg13g2_decap_4 FILLER_57_404 ();
 sg13g2_fill_2 FILLER_57_408 ();
 sg13g2_decap_8 FILLER_57_414 ();
 sg13g2_decap_8 FILLER_57_421 ();
 sg13g2_decap_4 FILLER_57_428 ();
 sg13g2_fill_2 FILLER_57_458 ();
 sg13g2_fill_1 FILLER_57_460 ();
 sg13g2_decap_4 FILLER_57_527 ();
 sg13g2_fill_2 FILLER_57_531 ();
 sg13g2_decap_4 FILLER_57_551 ();
 sg13g2_fill_1 FILLER_57_555 ();
 sg13g2_fill_2 FILLER_57_561 ();
 sg13g2_decap_8 FILLER_57_568 ();
 sg13g2_fill_2 FILLER_57_575 ();
 sg13g2_fill_2 FILLER_57_582 ();
 sg13g2_fill_1 FILLER_57_584 ();
 sg13g2_decap_8 FILLER_57_590 ();
 sg13g2_fill_2 FILLER_57_597 ();
 sg13g2_decap_4 FILLER_57_614 ();
 sg13g2_fill_2 FILLER_57_635 ();
 sg13g2_fill_1 FILLER_57_637 ();
 sg13g2_decap_8 FILLER_57_667 ();
 sg13g2_decap_8 FILLER_57_674 ();
 sg13g2_fill_1 FILLER_57_681 ();
 sg13g2_decap_8 FILLER_57_688 ();
 sg13g2_fill_2 FILLER_57_695 ();
 sg13g2_fill_1 FILLER_57_726 ();
 sg13g2_decap_4 FILLER_57_753 ();
 sg13g2_fill_1 FILLER_57_757 ();
 sg13g2_fill_2 FILLER_57_771 ();
 sg13g2_decap_8 FILLER_57_811 ();
 sg13g2_fill_1 FILLER_57_818 ();
 sg13g2_fill_2 FILLER_57_867 ();
 sg13g2_fill_1 FILLER_57_881 ();
 sg13g2_fill_2 FILLER_57_887 ();
 sg13g2_fill_2 FILLER_57_898 ();
 sg13g2_decap_4 FILLER_57_904 ();
 sg13g2_fill_1 FILLER_57_908 ();
 sg13g2_decap_8 FILLER_57_978 ();
 sg13g2_decap_4 FILLER_57_985 ();
 sg13g2_fill_1 FILLER_57_989 ();
 sg13g2_fill_1 FILLER_57_999 ();
 sg13g2_fill_1 FILLER_57_1010 ();
 sg13g2_fill_2 FILLER_57_1020 ();
 sg13g2_fill_1 FILLER_57_1022 ();
 sg13g2_decap_4 FILLER_57_1031 ();
 sg13g2_fill_2 FILLER_57_1035 ();
 sg13g2_fill_1 FILLER_57_1055 ();
 sg13g2_fill_2 FILLER_57_1075 ();
 sg13g2_fill_1 FILLER_57_1077 ();
 sg13g2_fill_1 FILLER_57_1110 ();
 sg13g2_fill_2 FILLER_57_1114 ();
 sg13g2_fill_1 FILLER_57_1116 ();
 sg13g2_fill_1 FILLER_57_1131 ();
 sg13g2_fill_1 FILLER_57_1141 ();
 sg13g2_fill_2 FILLER_57_1169 ();
 sg13g2_decap_4 FILLER_57_1250 ();
 sg13g2_fill_1 FILLER_57_1254 ();
 sg13g2_fill_2 FILLER_57_1264 ();
 sg13g2_fill_2 FILLER_57_1275 ();
 sg13g2_fill_1 FILLER_57_1277 ();
 sg13g2_fill_1 FILLER_57_1283 ();
 sg13g2_decap_8 FILLER_57_1298 ();
 sg13g2_decap_8 FILLER_57_1305 ();
 sg13g2_fill_2 FILLER_57_1312 ();
 sg13g2_fill_2 FILLER_57_1335 ();
 sg13g2_decap_8 FILLER_57_1346 ();
 sg13g2_fill_2 FILLER_57_1353 ();
 sg13g2_fill_1 FILLER_57_1407 ();
 sg13g2_fill_2 FILLER_57_1430 ();
 sg13g2_fill_1 FILLER_57_1432 ();
 sg13g2_fill_1 FILLER_57_1438 ();
 sg13g2_fill_2 FILLER_57_1462 ();
 sg13g2_fill_1 FILLER_57_1500 ();
 sg13g2_fill_1 FILLER_57_1515 ();
 sg13g2_fill_1 FILLER_57_1530 ();
 sg13g2_fill_2 FILLER_57_1543 ();
 sg13g2_decap_8 FILLER_57_1559 ();
 sg13g2_fill_2 FILLER_57_1566 ();
 sg13g2_fill_2 FILLER_57_1589 ();
 sg13g2_fill_1 FILLER_57_1591 ();
 sg13g2_fill_2 FILLER_57_1618 ();
 sg13g2_decap_4 FILLER_57_1642 ();
 sg13g2_fill_2 FILLER_57_1646 ();
 sg13g2_decap_4 FILLER_57_1661 ();
 sg13g2_fill_2 FILLER_57_1665 ();
 sg13g2_decap_4 FILLER_57_1674 ();
 sg13g2_fill_1 FILLER_57_1678 ();
 sg13g2_fill_2 FILLER_57_1696 ();
 sg13g2_decap_8 FILLER_57_1711 ();
 sg13g2_fill_2 FILLER_57_1718 ();
 sg13g2_fill_1 FILLER_57_1720 ();
 sg13g2_fill_2 FILLER_57_1743 ();
 sg13g2_fill_2 FILLER_57_1758 ();
 sg13g2_fill_2 FILLER_57_1765 ();
 sg13g2_decap_8 FILLER_57_1773 ();
 sg13g2_fill_1 FILLER_57_1780 ();
 sg13g2_decap_8 FILLER_57_1794 ();
 sg13g2_decap_4 FILLER_57_1817 ();
 sg13g2_decap_4 FILLER_57_1836 ();
 sg13g2_fill_2 FILLER_57_1840 ();
 sg13g2_fill_2 FILLER_57_1859 ();
 sg13g2_fill_1 FILLER_57_1861 ();
 sg13g2_fill_1 FILLER_57_1884 ();
 sg13g2_decap_8 FILLER_57_1907 ();
 sg13g2_decap_8 FILLER_57_1939 ();
 sg13g2_fill_2 FILLER_57_1946 ();
 sg13g2_fill_1 FILLER_57_1960 ();
 sg13g2_fill_1 FILLER_57_1977 ();
 sg13g2_fill_1 FILLER_57_2000 ();
 sg13g2_fill_2 FILLER_57_2055 ();
 sg13g2_decap_4 FILLER_57_2071 ();
 sg13g2_fill_2 FILLER_57_2080 ();
 sg13g2_fill_1 FILLER_57_2082 ();
 sg13g2_decap_8 FILLER_57_2100 ();
 sg13g2_decap_8 FILLER_57_2107 ();
 sg13g2_fill_2 FILLER_57_2114 ();
 sg13g2_fill_1 FILLER_57_2125 ();
 sg13g2_decap_4 FILLER_57_2130 ();
 sg13g2_decap_8 FILLER_57_2138 ();
 sg13g2_fill_2 FILLER_57_2145 ();
 sg13g2_decap_8 FILLER_57_2157 ();
 sg13g2_decap_4 FILLER_57_2164 ();
 sg13g2_fill_1 FILLER_57_2177 ();
 sg13g2_decap_8 FILLER_57_2188 ();
 sg13g2_decap_4 FILLER_57_2195 ();
 sg13g2_fill_2 FILLER_57_2199 ();
 sg13g2_decap_8 FILLER_57_2216 ();
 sg13g2_fill_2 FILLER_57_2223 ();
 sg13g2_fill_1 FILLER_57_2225 ();
 sg13g2_decap_4 FILLER_57_2234 ();
 sg13g2_fill_1 FILLER_57_2238 ();
 sg13g2_decap_8 FILLER_57_2248 ();
 sg13g2_decap_8 FILLER_57_2255 ();
 sg13g2_fill_2 FILLER_57_2262 ();
 sg13g2_decap_8 FILLER_57_2291 ();
 sg13g2_fill_1 FILLER_57_2298 ();
 sg13g2_decap_4 FILLER_57_2303 ();
 sg13g2_fill_1 FILLER_57_2312 ();
 sg13g2_decap_8 FILLER_57_2323 ();
 sg13g2_fill_2 FILLER_57_2330 ();
 sg13g2_fill_1 FILLER_57_2332 ();
 sg13g2_decap_4 FILLER_57_2350 ();
 sg13g2_fill_2 FILLER_57_2354 ();
 sg13g2_decap_8 FILLER_57_2371 ();
 sg13g2_fill_1 FILLER_57_2386 ();
 sg13g2_fill_1 FILLER_57_2391 ();
 sg13g2_decap_8 FILLER_57_2442 ();
 sg13g2_decap_4 FILLER_57_2449 ();
 sg13g2_fill_1 FILLER_57_2472 ();
 sg13g2_fill_2 FILLER_57_2528 ();
 sg13g2_fill_1 FILLER_57_2530 ();
 sg13g2_fill_2 FILLER_57_2565 ();
 sg13g2_decap_8 FILLER_57_2605 ();
 sg13g2_fill_2 FILLER_57_2612 ();
 sg13g2_fill_1 FILLER_57_2614 ();
 sg13g2_decap_8 FILLER_57_2633 ();
 sg13g2_decap_8 FILLER_57_2640 ();
 sg13g2_fill_2 FILLER_57_2647 ();
 sg13g2_fill_2 FILLER_57_2653 ();
 sg13g2_fill_1 FILLER_57_2655 ();
 sg13g2_decap_4 FILLER_57_2660 ();
 sg13g2_fill_1 FILLER_57_2664 ();
 sg13g2_decap_4 FILLER_57_2681 ();
 sg13g2_fill_2 FILLER_57_2685 ();
 sg13g2_decap_8 FILLER_57_2697 ();
 sg13g2_fill_2 FILLER_57_2704 ();
 sg13g2_fill_1 FILLER_57_2706 ();
 sg13g2_decap_8 FILLER_57_2722 ();
 sg13g2_fill_2 FILLER_57_2745 ();
 sg13g2_decap_8 FILLER_57_2763 ();
 sg13g2_fill_2 FILLER_57_2775 ();
 sg13g2_fill_1 FILLER_57_2777 ();
 sg13g2_decap_4 FILLER_57_2799 ();
 sg13g2_decap_4 FILLER_57_2807 ();
 sg13g2_decap_4 FILLER_57_2838 ();
 sg13g2_fill_1 FILLER_57_2842 ();
 sg13g2_fill_1 FILLER_57_2848 ();
 sg13g2_fill_2 FILLER_57_2854 ();
 sg13g2_decap_8 FILLER_57_2869 ();
 sg13g2_fill_2 FILLER_57_2876 ();
 sg13g2_fill_1 FILLER_57_2878 ();
 sg13g2_decap_8 FILLER_57_2890 ();
 sg13g2_decap_8 FILLER_57_2897 ();
 sg13g2_fill_2 FILLER_57_2904 ();
 sg13g2_fill_1 FILLER_57_2906 ();
 sg13g2_decap_4 FILLER_57_2912 ();
 sg13g2_fill_2 FILLER_57_2916 ();
 sg13g2_decap_8 FILLER_57_2930 ();
 sg13g2_decap_4 FILLER_57_2937 ();
 sg13g2_fill_1 FILLER_57_2941 ();
 sg13g2_fill_2 FILLER_57_2965 ();
 sg13g2_fill_1 FILLER_57_2967 ();
 sg13g2_decap_8 FILLER_57_2994 ();
 sg13g2_decap_8 FILLER_57_3001 ();
 sg13g2_decap_8 FILLER_57_3008 ();
 sg13g2_decap_8 FILLER_57_3015 ();
 sg13g2_decap_8 FILLER_57_3022 ();
 sg13g2_decap_8 FILLER_57_3029 ();
 sg13g2_decap_8 FILLER_57_3036 ();
 sg13g2_decap_8 FILLER_57_3043 ();
 sg13g2_decap_8 FILLER_57_3050 ();
 sg13g2_decap_8 FILLER_57_3057 ();
 sg13g2_decap_8 FILLER_57_3064 ();
 sg13g2_decap_8 FILLER_57_3071 ();
 sg13g2_decap_8 FILLER_57_3078 ();
 sg13g2_decap_8 FILLER_57_3085 ();
 sg13g2_decap_8 FILLER_57_3092 ();
 sg13g2_decap_8 FILLER_57_3099 ();
 sg13g2_decap_8 FILLER_57_3106 ();
 sg13g2_decap_8 FILLER_57_3113 ();
 sg13g2_decap_8 FILLER_57_3120 ();
 sg13g2_decap_8 FILLER_57_3127 ();
 sg13g2_decap_8 FILLER_57_3134 ();
 sg13g2_decap_8 FILLER_57_3141 ();
 sg13g2_decap_8 FILLER_57_3148 ();
 sg13g2_decap_8 FILLER_57_3155 ();
 sg13g2_decap_8 FILLER_57_3162 ();
 sg13g2_decap_8 FILLER_57_3169 ();
 sg13g2_decap_8 FILLER_57_3176 ();
 sg13g2_decap_8 FILLER_57_3183 ();
 sg13g2_decap_8 FILLER_57_3190 ();
 sg13g2_decap_8 FILLER_57_3197 ();
 sg13g2_decap_8 FILLER_57_3204 ();
 sg13g2_decap_8 FILLER_57_3211 ();
 sg13g2_decap_8 FILLER_57_3218 ();
 sg13g2_decap_8 FILLER_57_3225 ();
 sg13g2_decap_8 FILLER_57_3232 ();
 sg13g2_decap_8 FILLER_57_3239 ();
 sg13g2_decap_8 FILLER_57_3246 ();
 sg13g2_decap_8 FILLER_57_3253 ();
 sg13g2_decap_8 FILLER_57_3260 ();
 sg13g2_decap_8 FILLER_57_3267 ();
 sg13g2_decap_8 FILLER_57_3274 ();
 sg13g2_decap_8 FILLER_57_3281 ();
 sg13g2_decap_8 FILLER_57_3288 ();
 sg13g2_decap_8 FILLER_57_3295 ();
 sg13g2_decap_8 FILLER_57_3302 ();
 sg13g2_decap_8 FILLER_57_3309 ();
 sg13g2_decap_8 FILLER_57_3316 ();
 sg13g2_decap_8 FILLER_57_3323 ();
 sg13g2_decap_8 FILLER_57_3330 ();
 sg13g2_decap_8 FILLER_57_3337 ();
 sg13g2_decap_8 FILLER_57_3344 ();
 sg13g2_decap_8 FILLER_57_3351 ();
 sg13g2_decap_8 FILLER_57_3358 ();
 sg13g2_decap_8 FILLER_57_3365 ();
 sg13g2_decap_8 FILLER_57_3372 ();
 sg13g2_decap_8 FILLER_57_3379 ();
 sg13g2_decap_8 FILLER_57_3386 ();
 sg13g2_decap_8 FILLER_57_3393 ();
 sg13g2_decap_8 FILLER_57_3400 ();
 sg13g2_decap_8 FILLER_57_3407 ();
 sg13g2_decap_8 FILLER_57_3414 ();
 sg13g2_decap_8 FILLER_57_3421 ();
 sg13g2_decap_8 FILLER_57_3428 ();
 sg13g2_decap_8 FILLER_57_3435 ();
 sg13g2_decap_8 FILLER_57_3442 ();
 sg13g2_decap_8 FILLER_57_3449 ();
 sg13g2_decap_8 FILLER_57_3456 ();
 sg13g2_decap_8 FILLER_57_3463 ();
 sg13g2_decap_8 FILLER_57_3470 ();
 sg13g2_decap_8 FILLER_57_3477 ();
 sg13g2_decap_8 FILLER_57_3484 ();
 sg13g2_decap_8 FILLER_57_3491 ();
 sg13g2_decap_8 FILLER_57_3498 ();
 sg13g2_decap_8 FILLER_57_3505 ();
 sg13g2_decap_8 FILLER_57_3512 ();
 sg13g2_decap_8 FILLER_57_3519 ();
 sg13g2_decap_8 FILLER_57_3526 ();
 sg13g2_decap_8 FILLER_57_3533 ();
 sg13g2_decap_8 FILLER_57_3540 ();
 sg13g2_decap_8 FILLER_57_3547 ();
 sg13g2_decap_8 FILLER_57_3554 ();
 sg13g2_decap_8 FILLER_57_3561 ();
 sg13g2_decap_8 FILLER_57_3568 ();
 sg13g2_decap_4 FILLER_57_3575 ();
 sg13g2_fill_1 FILLER_57_3579 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_18 ();
 sg13g2_fill_2 FILLER_58_25 ();
 sg13g2_fill_2 FILLER_58_36 ();
 sg13g2_decap_4 FILLER_58_58 ();
 sg13g2_fill_1 FILLER_58_62 ();
 sg13g2_decap_8 FILLER_58_90 ();
 sg13g2_decap_4 FILLER_58_97 ();
 sg13g2_fill_2 FILLER_58_235 ();
 sg13g2_fill_1 FILLER_58_237 ();
 sg13g2_fill_1 FILLER_58_286 ();
 sg13g2_fill_2 FILLER_58_296 ();
 sg13g2_fill_2 FILLER_58_311 ();
 sg13g2_fill_1 FILLER_58_313 ();
 sg13g2_fill_2 FILLER_58_379 ();
 sg13g2_fill_1 FILLER_58_381 ();
 sg13g2_fill_2 FILLER_58_391 ();
 sg13g2_fill_2 FILLER_58_396 ();
 sg13g2_decap_4 FILLER_58_402 ();
 sg13g2_fill_2 FILLER_58_411 ();
 sg13g2_fill_1 FILLER_58_413 ();
 sg13g2_fill_2 FILLER_58_422 ();
 sg13g2_decap_4 FILLER_58_437 ();
 sg13g2_fill_1 FILLER_58_483 ();
 sg13g2_decap_8 FILLER_58_489 ();
 sg13g2_fill_2 FILLER_58_496 ();
 sg13g2_fill_1 FILLER_58_498 ();
 sg13g2_fill_1 FILLER_58_513 ();
 sg13g2_fill_2 FILLER_58_519 ();
 sg13g2_decap_4 FILLER_58_526 ();
 sg13g2_fill_2 FILLER_58_530 ();
 sg13g2_fill_2 FILLER_58_546 ();
 sg13g2_fill_1 FILLER_58_548 ();
 sg13g2_decap_4 FILLER_58_598 ();
 sg13g2_decap_4 FILLER_58_618 ();
 sg13g2_fill_2 FILLER_58_622 ();
 sg13g2_fill_2 FILLER_58_630 ();
 sg13g2_decap_8 FILLER_58_658 ();
 sg13g2_fill_1 FILLER_58_665 ();
 sg13g2_fill_1 FILLER_58_691 ();
 sg13g2_fill_2 FILLER_58_747 ();
 sg13g2_decap_8 FILLER_58_766 ();
 sg13g2_fill_2 FILLER_58_773 ();
 sg13g2_fill_1 FILLER_58_775 ();
 sg13g2_decap_8 FILLER_58_788 ();
 sg13g2_fill_2 FILLER_58_800 ();
 sg13g2_decap_4 FILLER_58_818 ();
 sg13g2_fill_1 FILLER_58_822 ();
 sg13g2_fill_2 FILLER_58_828 ();
 sg13g2_fill_2 FILLER_58_849 ();
 sg13g2_fill_1 FILLER_58_851 ();
 sg13g2_fill_2 FILLER_58_861 ();
 sg13g2_decap_8 FILLER_58_895 ();
 sg13g2_fill_1 FILLER_58_902 ();
 sg13g2_fill_1 FILLER_58_929 ();
 sg13g2_fill_2 FILLER_58_943 ();
 sg13g2_fill_1 FILLER_58_945 ();
 sg13g2_fill_1 FILLER_58_1015 ();
 sg13g2_decap_8 FILLER_58_1020 ();
 sg13g2_fill_2 FILLER_58_1027 ();
 sg13g2_fill_2 FILLER_58_1060 ();
 sg13g2_decap_4 FILLER_58_1071 ();
 sg13g2_fill_1 FILLER_58_1075 ();
 sg13g2_decap_8 FILLER_58_1081 ();
 sg13g2_fill_2 FILLER_58_1119 ();
 sg13g2_fill_1 FILLER_58_1121 ();
 sg13g2_fill_2 FILLER_58_1146 ();
 sg13g2_fill_1 FILLER_58_1148 ();
 sg13g2_fill_2 FILLER_58_1167 ();
 sg13g2_fill_2 FILLER_58_1181 ();
 sg13g2_fill_1 FILLER_58_1183 ();
 sg13g2_fill_2 FILLER_58_1224 ();
 sg13g2_fill_1 FILLER_58_1226 ();
 sg13g2_fill_2 FILLER_58_1232 ();
 sg13g2_fill_1 FILLER_58_1234 ();
 sg13g2_decap_8 FILLER_58_1264 ();
 sg13g2_fill_2 FILLER_58_1306 ();
 sg13g2_decap_8 FILLER_58_1330 ();
 sg13g2_fill_2 FILLER_58_1337 ();
 sg13g2_decap_8 FILLER_58_1342 ();
 sg13g2_decap_4 FILLER_58_1375 ();
 sg13g2_fill_1 FILLER_58_1388 ();
 sg13g2_fill_1 FILLER_58_1400 ();
 sg13g2_decap_8 FILLER_58_1411 ();
 sg13g2_fill_2 FILLER_58_1418 ();
 sg13g2_fill_2 FILLER_58_1436 ();
 sg13g2_decap_8 FILLER_58_1464 ();
 sg13g2_fill_1 FILLER_58_1471 ();
 sg13g2_decap_4 FILLER_58_1498 ();
 sg13g2_fill_2 FILLER_58_1502 ();
 sg13g2_fill_2 FILLER_58_1516 ();
 sg13g2_fill_1 FILLER_58_1518 ();
 sg13g2_decap_4 FILLER_58_1589 ();
 sg13g2_decap_8 FILLER_58_1607 ();
 sg13g2_fill_2 FILLER_58_1614 ();
 sg13g2_fill_1 FILLER_58_1624 ();
 sg13g2_fill_2 FILLER_58_1638 ();
 sg13g2_fill_2 FILLER_58_1670 ();
 sg13g2_fill_1 FILLER_58_1672 ();
 sg13g2_fill_2 FILLER_58_1693 ();
 sg13g2_fill_2 FILLER_58_1717 ();
 sg13g2_fill_1 FILLER_58_1719 ();
 sg13g2_fill_2 FILLER_58_1728 ();
 sg13g2_decap_4 FILLER_58_1749 ();
 sg13g2_fill_1 FILLER_58_1753 ();
 sg13g2_decap_4 FILLER_58_1776 ();
 sg13g2_fill_2 FILLER_58_1780 ();
 sg13g2_decap_8 FILLER_58_1790 ();
 sg13g2_fill_2 FILLER_58_1805 ();
 sg13g2_fill_1 FILLER_58_1837 ();
 sg13g2_fill_2 FILLER_58_1844 ();
 sg13g2_fill_1 FILLER_58_1846 ();
 sg13g2_fill_2 FILLER_58_1877 ();
 sg13g2_fill_1 FILLER_58_1879 ();
 sg13g2_decap_8 FILLER_58_1889 ();
 sg13g2_fill_1 FILLER_58_1896 ();
 sg13g2_decap_8 FILLER_58_1918 ();
 sg13g2_decap_8 FILLER_58_1925 ();
 sg13g2_decap_4 FILLER_58_1932 ();
 sg13g2_decap_8 FILLER_58_1952 ();
 sg13g2_decap_8 FILLER_58_1959 ();
 sg13g2_decap_8 FILLER_58_1966 ();
 sg13g2_fill_2 FILLER_58_1973 ();
 sg13g2_decap_4 FILLER_58_1996 ();
 sg13g2_fill_2 FILLER_58_2000 ();
 sg13g2_decap_8 FILLER_58_2005 ();
 sg13g2_decap_4 FILLER_58_2012 ();
 sg13g2_fill_2 FILLER_58_2016 ();
 sg13g2_fill_2 FILLER_58_2027 ();
 sg13g2_decap_4 FILLER_58_2034 ();
 sg13g2_fill_1 FILLER_58_2038 ();
 sg13g2_fill_1 FILLER_58_2052 ();
 sg13g2_fill_1 FILLER_58_2058 ();
 sg13g2_decap_4 FILLER_58_2069 ();
 sg13g2_decap_4 FILLER_58_2091 ();
 sg13g2_fill_1 FILLER_58_2107 ();
 sg13g2_decap_8 FILLER_58_2119 ();
 sg13g2_decap_8 FILLER_58_2126 ();
 sg13g2_decap_4 FILLER_58_2133 ();
 sg13g2_fill_1 FILLER_58_2137 ();
 sg13g2_decap_4 FILLER_58_2153 ();
 sg13g2_decap_4 FILLER_58_2180 ();
 sg13g2_fill_1 FILLER_58_2184 ();
 sg13g2_decap_4 FILLER_58_2190 ();
 sg13g2_fill_2 FILLER_58_2194 ();
 sg13g2_decap_8 FILLER_58_2213 ();
 sg13g2_decap_8 FILLER_58_2220 ();
 sg13g2_fill_1 FILLER_58_2227 ();
 sg13g2_fill_1 FILLER_58_2246 ();
 sg13g2_decap_8 FILLER_58_2250 ();
 sg13g2_fill_2 FILLER_58_2257 ();
 sg13g2_fill_1 FILLER_58_2259 ();
 sg13g2_fill_1 FILLER_58_2272 ();
 sg13g2_decap_8 FILLER_58_2283 ();
 sg13g2_decap_4 FILLER_58_2290 ();
 sg13g2_fill_1 FILLER_58_2294 ();
 sg13g2_fill_1 FILLER_58_2321 ();
 sg13g2_decap_8 FILLER_58_2348 ();
 sg13g2_fill_1 FILLER_58_2355 ();
 sg13g2_fill_2 FILLER_58_2379 ();
 sg13g2_decap_4 FILLER_58_2394 ();
 sg13g2_fill_1 FILLER_58_2398 ();
 sg13g2_fill_1 FILLER_58_2404 ();
 sg13g2_fill_2 FILLER_58_2410 ();
 sg13g2_fill_1 FILLER_58_2412 ();
 sg13g2_fill_2 FILLER_58_2431 ();
 sg13g2_fill_1 FILLER_58_2441 ();
 sg13g2_fill_2 FILLER_58_2447 ();
 sg13g2_decap_8 FILLER_58_2474 ();
 sg13g2_decap_8 FILLER_58_2481 ();
 sg13g2_decap_4 FILLER_58_2488 ();
 sg13g2_decap_8 FILLER_58_2496 ();
 sg13g2_decap_4 FILLER_58_2503 ();
 sg13g2_fill_1 FILLER_58_2507 ();
 sg13g2_decap_8 FILLER_58_2532 ();
 sg13g2_fill_2 FILLER_58_2539 ();
 sg13g2_decap_8 FILLER_58_2567 ();
 sg13g2_decap_8 FILLER_58_2574 ();
 sg13g2_decap_4 FILLER_58_2581 ();
 sg13g2_fill_1 FILLER_58_2585 ();
 sg13g2_fill_2 FILLER_58_2599 ();
 sg13g2_decap_8 FILLER_58_2611 ();
 sg13g2_decap_4 FILLER_58_2618 ();
 sg13g2_fill_2 FILLER_58_2622 ();
 sg13g2_decap_8 FILLER_58_2634 ();
 sg13g2_decap_8 FILLER_58_2641 ();
 sg13g2_fill_2 FILLER_58_2648 ();
 sg13g2_fill_1 FILLER_58_2658 ();
 sg13g2_fill_2 FILLER_58_2669 ();
 sg13g2_decap_8 FILLER_58_2685 ();
 sg13g2_fill_2 FILLER_58_2696 ();
 sg13g2_fill_2 FILLER_58_2702 ();
 sg13g2_fill_1 FILLER_58_2704 ();
 sg13g2_decap_4 FILLER_58_2710 ();
 sg13g2_fill_1 FILLER_58_2714 ();
 sg13g2_decap_8 FILLER_58_2723 ();
 sg13g2_decap_8 FILLER_58_2735 ();
 sg13g2_decap_4 FILLER_58_2742 ();
 sg13g2_decap_8 FILLER_58_2759 ();
 sg13g2_decap_8 FILLER_58_2778 ();
 sg13g2_decap_8 FILLER_58_2790 ();
 sg13g2_decap_8 FILLER_58_2797 ();
 sg13g2_fill_1 FILLER_58_2804 ();
 sg13g2_fill_2 FILLER_58_2815 ();
 sg13g2_decap_4 FILLER_58_2839 ();
 sg13g2_fill_2 FILLER_58_2843 ();
 sg13g2_fill_1 FILLER_58_2867 ();
 sg13g2_decap_8 FILLER_58_2894 ();
 sg13g2_fill_2 FILLER_58_2901 ();
 sg13g2_fill_1 FILLER_58_2903 ();
 sg13g2_fill_2 FILLER_58_2939 ();
 sg13g2_fill_1 FILLER_58_2941 ();
 sg13g2_decap_8 FILLER_58_2947 ();
 sg13g2_fill_2 FILLER_58_2954 ();
 sg13g2_fill_1 FILLER_58_2956 ();
 sg13g2_fill_2 FILLER_58_2967 ();
 sg13g2_fill_1 FILLER_58_2978 ();
 sg13g2_decap_8 FILLER_58_3012 ();
 sg13g2_decap_8 FILLER_58_3019 ();
 sg13g2_decap_8 FILLER_58_3026 ();
 sg13g2_decap_8 FILLER_58_3033 ();
 sg13g2_decap_8 FILLER_58_3040 ();
 sg13g2_decap_8 FILLER_58_3047 ();
 sg13g2_decap_8 FILLER_58_3054 ();
 sg13g2_decap_8 FILLER_58_3061 ();
 sg13g2_decap_8 FILLER_58_3068 ();
 sg13g2_decap_8 FILLER_58_3075 ();
 sg13g2_decap_8 FILLER_58_3082 ();
 sg13g2_decap_8 FILLER_58_3089 ();
 sg13g2_decap_8 FILLER_58_3096 ();
 sg13g2_decap_8 FILLER_58_3103 ();
 sg13g2_decap_8 FILLER_58_3110 ();
 sg13g2_decap_8 FILLER_58_3117 ();
 sg13g2_decap_8 FILLER_58_3124 ();
 sg13g2_decap_8 FILLER_58_3131 ();
 sg13g2_decap_8 FILLER_58_3138 ();
 sg13g2_decap_8 FILLER_58_3145 ();
 sg13g2_decap_8 FILLER_58_3152 ();
 sg13g2_decap_8 FILLER_58_3159 ();
 sg13g2_decap_8 FILLER_58_3166 ();
 sg13g2_decap_8 FILLER_58_3173 ();
 sg13g2_decap_8 FILLER_58_3180 ();
 sg13g2_decap_8 FILLER_58_3187 ();
 sg13g2_decap_8 FILLER_58_3194 ();
 sg13g2_decap_8 FILLER_58_3201 ();
 sg13g2_decap_8 FILLER_58_3208 ();
 sg13g2_decap_8 FILLER_58_3215 ();
 sg13g2_decap_8 FILLER_58_3222 ();
 sg13g2_decap_8 FILLER_58_3229 ();
 sg13g2_decap_8 FILLER_58_3236 ();
 sg13g2_decap_8 FILLER_58_3243 ();
 sg13g2_decap_8 FILLER_58_3250 ();
 sg13g2_decap_8 FILLER_58_3257 ();
 sg13g2_decap_8 FILLER_58_3264 ();
 sg13g2_decap_8 FILLER_58_3271 ();
 sg13g2_decap_8 FILLER_58_3278 ();
 sg13g2_decap_8 FILLER_58_3285 ();
 sg13g2_decap_8 FILLER_58_3292 ();
 sg13g2_decap_8 FILLER_58_3299 ();
 sg13g2_decap_8 FILLER_58_3306 ();
 sg13g2_decap_8 FILLER_58_3313 ();
 sg13g2_decap_8 FILLER_58_3320 ();
 sg13g2_decap_8 FILLER_58_3327 ();
 sg13g2_decap_8 FILLER_58_3334 ();
 sg13g2_decap_8 FILLER_58_3341 ();
 sg13g2_decap_8 FILLER_58_3348 ();
 sg13g2_decap_8 FILLER_58_3355 ();
 sg13g2_decap_8 FILLER_58_3362 ();
 sg13g2_decap_8 FILLER_58_3369 ();
 sg13g2_decap_8 FILLER_58_3376 ();
 sg13g2_decap_8 FILLER_58_3383 ();
 sg13g2_decap_8 FILLER_58_3390 ();
 sg13g2_decap_8 FILLER_58_3397 ();
 sg13g2_decap_8 FILLER_58_3404 ();
 sg13g2_decap_8 FILLER_58_3411 ();
 sg13g2_decap_8 FILLER_58_3418 ();
 sg13g2_decap_8 FILLER_58_3425 ();
 sg13g2_decap_8 FILLER_58_3432 ();
 sg13g2_decap_8 FILLER_58_3439 ();
 sg13g2_decap_8 FILLER_58_3446 ();
 sg13g2_decap_8 FILLER_58_3453 ();
 sg13g2_decap_8 FILLER_58_3460 ();
 sg13g2_decap_8 FILLER_58_3467 ();
 sg13g2_decap_8 FILLER_58_3474 ();
 sg13g2_decap_8 FILLER_58_3481 ();
 sg13g2_decap_8 FILLER_58_3488 ();
 sg13g2_decap_8 FILLER_58_3495 ();
 sg13g2_decap_8 FILLER_58_3502 ();
 sg13g2_decap_8 FILLER_58_3509 ();
 sg13g2_decap_8 FILLER_58_3516 ();
 sg13g2_decap_8 FILLER_58_3523 ();
 sg13g2_decap_8 FILLER_58_3530 ();
 sg13g2_decap_8 FILLER_58_3537 ();
 sg13g2_decap_8 FILLER_58_3544 ();
 sg13g2_decap_8 FILLER_58_3551 ();
 sg13g2_decap_8 FILLER_58_3558 ();
 sg13g2_decap_8 FILLER_58_3565 ();
 sg13g2_decap_8 FILLER_58_3572 ();
 sg13g2_fill_1 FILLER_58_3579 ();
 sg13g2_decap_4 FILLER_59_56 ();
 sg13g2_fill_1 FILLER_59_83 ();
 sg13g2_decap_4 FILLER_59_113 ();
 sg13g2_fill_1 FILLER_59_117 ();
 sg13g2_fill_2 FILLER_59_122 ();
 sg13g2_fill_1 FILLER_59_129 ();
 sg13g2_decap_8 FILLER_59_140 ();
 sg13g2_decap_8 FILLER_59_147 ();
 sg13g2_fill_2 FILLER_59_172 ();
 sg13g2_fill_1 FILLER_59_183 ();
 sg13g2_fill_1 FILLER_59_194 ();
 sg13g2_fill_2 FILLER_59_214 ();
 sg13g2_decap_4 FILLER_59_243 ();
 sg13g2_fill_2 FILLER_59_247 ();
 sg13g2_fill_1 FILLER_59_262 ();
 sg13g2_decap_4 FILLER_59_281 ();
 sg13g2_fill_1 FILLER_59_306 ();
 sg13g2_decap_8 FILLER_59_312 ();
 sg13g2_decap_8 FILLER_59_319 ();
 sg13g2_fill_1 FILLER_59_326 ();
 sg13g2_fill_2 FILLER_59_336 ();
 sg13g2_decap_8 FILLER_59_356 ();
 sg13g2_fill_2 FILLER_59_363 ();
 sg13g2_decap_8 FILLER_59_370 ();
 sg13g2_fill_1 FILLER_59_377 ();
 sg13g2_decap_8 FILLER_59_413 ();
 sg13g2_fill_2 FILLER_59_420 ();
 sg13g2_fill_2 FILLER_59_438 ();
 sg13g2_decap_8 FILLER_59_444 ();
 sg13g2_decap_4 FILLER_59_451 ();
 sg13g2_fill_1 FILLER_59_455 ();
 sg13g2_fill_1 FILLER_59_469 ();
 sg13g2_fill_2 FILLER_59_484 ();
 sg13g2_fill_2 FILLER_59_496 ();
 sg13g2_fill_1 FILLER_59_498 ();
 sg13g2_fill_1 FILLER_59_507 ();
 sg13g2_decap_4 FILLER_59_553 ();
 sg13g2_fill_1 FILLER_59_557 ();
 sg13g2_decap_8 FILLER_59_568 ();
 sg13g2_fill_1 FILLER_59_575 ();
 sg13g2_fill_2 FILLER_59_587 ();
 sg13g2_fill_1 FILLER_59_589 ();
 sg13g2_fill_1 FILLER_59_598 ();
 sg13g2_fill_2 FILLER_59_613 ();
 sg13g2_fill_2 FILLER_59_619 ();
 sg13g2_decap_8 FILLER_59_627 ();
 sg13g2_decap_4 FILLER_59_634 ();
 sg13g2_decap_4 FILLER_59_644 ();
 sg13g2_fill_2 FILLER_59_648 ();
 sg13g2_fill_2 FILLER_59_661 ();
 sg13g2_fill_1 FILLER_59_674 ();
 sg13g2_fill_1 FILLER_59_683 ();
 sg13g2_fill_2 FILLER_59_693 ();
 sg13g2_fill_1 FILLER_59_711 ();
 sg13g2_fill_1 FILLER_59_723 ();
 sg13g2_decap_8 FILLER_59_775 ();
 sg13g2_fill_2 FILLER_59_782 ();
 sg13g2_fill_2 FILLER_59_789 ();
 sg13g2_fill_1 FILLER_59_791 ();
 sg13g2_decap_4 FILLER_59_824 ();
 sg13g2_fill_2 FILLER_59_868 ();
 sg13g2_fill_1 FILLER_59_878 ();
 sg13g2_fill_2 FILLER_59_896 ();
 sg13g2_fill_2 FILLER_59_931 ();
 sg13g2_fill_1 FILLER_59_933 ();
 sg13g2_decap_8 FILLER_59_954 ();
 sg13g2_decap_8 FILLER_59_961 ();
 sg13g2_decap_8 FILLER_59_968 ();
 sg13g2_decap_8 FILLER_59_975 ();
 sg13g2_decap_4 FILLER_59_982 ();
 sg13g2_fill_1 FILLER_59_986 ();
 sg13g2_fill_1 FILLER_59_1001 ();
 sg13g2_fill_1 FILLER_59_1013 ();
 sg13g2_decap_4 FILLER_59_1018 ();
 sg13g2_decap_4 FILLER_59_1031 ();
 sg13g2_decap_4 FILLER_59_1039 ();
 sg13g2_fill_2 FILLER_59_1043 ();
 sg13g2_fill_2 FILLER_59_1049 ();
 sg13g2_fill_2 FILLER_59_1066 ();
 sg13g2_decap_4 FILLER_59_1076 ();
 sg13g2_decap_4 FILLER_59_1135 ();
 sg13g2_fill_1 FILLER_59_1139 ();
 sg13g2_decap_4 FILLER_59_1179 ();
 sg13g2_fill_1 FILLER_59_1183 ();
 sg13g2_fill_2 FILLER_59_1213 ();
 sg13g2_decap_4 FILLER_59_1250 ();
 sg13g2_fill_2 FILLER_59_1285 ();
 sg13g2_fill_2 FILLER_59_1302 ();
 sg13g2_fill_1 FILLER_59_1304 ();
 sg13g2_fill_2 FILLER_59_1367 ();
 sg13g2_fill_1 FILLER_59_1403 ();
 sg13g2_fill_2 FILLER_59_1439 ();
 sg13g2_fill_1 FILLER_59_1441 ();
 sg13g2_decap_4 FILLER_59_1455 ();
 sg13g2_fill_1 FILLER_59_1459 ();
 sg13g2_fill_2 FILLER_59_1468 ();
 sg13g2_fill_2 FILLER_59_1493 ();
 sg13g2_decap_8 FILLER_59_1500 ();
 sg13g2_fill_2 FILLER_59_1507 ();
 sg13g2_decap_8 FILLER_59_1537 ();
 sg13g2_decap_8 FILLER_59_1544 ();
 sg13g2_decap_8 FILLER_59_1551 ();
 sg13g2_decap_8 FILLER_59_1558 ();
 sg13g2_fill_1 FILLER_59_1565 ();
 sg13g2_fill_1 FILLER_59_1571 ();
 sg13g2_decap_8 FILLER_59_1581 ();
 sg13g2_decap_4 FILLER_59_1588 ();
 sg13g2_decap_4 FILLER_59_1627 ();
 sg13g2_fill_2 FILLER_59_1631 ();
 sg13g2_decap_8 FILLER_59_1641 ();
 sg13g2_decap_8 FILLER_59_1648 ();
 sg13g2_decap_8 FILLER_59_1659 ();
 sg13g2_decap_8 FILLER_59_1666 ();
 sg13g2_fill_2 FILLER_59_1673 ();
 sg13g2_fill_1 FILLER_59_1675 ();
 sg13g2_decap_4 FILLER_59_1692 ();
 sg13g2_fill_1 FILLER_59_1696 ();
 sg13g2_decap_8 FILLER_59_1708 ();
 sg13g2_decap_4 FILLER_59_1715 ();
 sg13g2_decap_8 FILLER_59_1729 ();
 sg13g2_fill_2 FILLER_59_1736 ();
 sg13g2_fill_1 FILLER_59_1738 ();
 sg13g2_decap_8 FILLER_59_1744 ();
 sg13g2_fill_1 FILLER_59_1767 ();
 sg13g2_decap_8 FILLER_59_1803 ();
 sg13g2_decap_8 FILLER_59_1810 ();
 sg13g2_fill_2 FILLER_59_1817 ();
 sg13g2_fill_1 FILLER_59_1819 ();
 sg13g2_fill_2 FILLER_59_1829 ();
 sg13g2_fill_1 FILLER_59_1831 ();
 sg13g2_decap_4 FILLER_59_1863 ();
 sg13g2_decap_8 FILLER_59_1893 ();
 sg13g2_fill_1 FILLER_59_1900 ();
 sg13g2_decap_4 FILLER_59_1914 ();
 sg13g2_fill_2 FILLER_59_1918 ();
 sg13g2_fill_2 FILLER_59_1956 ();
 sg13g2_decap_8 FILLER_59_1971 ();
 sg13g2_decap_4 FILLER_59_1978 ();
 sg13g2_fill_1 FILLER_59_1982 ();
 sg13g2_decap_4 FILLER_59_1997 ();
 sg13g2_fill_2 FILLER_59_2006 ();
 sg13g2_fill_1 FILLER_59_2008 ();
 sg13g2_decap_4 FILLER_59_2016 ();
 sg13g2_fill_2 FILLER_59_2020 ();
 sg13g2_decap_4 FILLER_59_2027 ();
 sg13g2_fill_2 FILLER_59_2031 ();
 sg13g2_fill_2 FILLER_59_2045 ();
 sg13g2_fill_1 FILLER_59_2047 ();
 sg13g2_fill_2 FILLER_59_2068 ();
 sg13g2_fill_1 FILLER_59_2070 ();
 sg13g2_decap_4 FILLER_59_2074 ();
 sg13g2_fill_2 FILLER_59_2078 ();
 sg13g2_decap_8 FILLER_59_2085 ();
 sg13g2_fill_2 FILLER_59_2092 ();
 sg13g2_decap_8 FILLER_59_2100 ();
 sg13g2_decap_4 FILLER_59_2127 ();
 sg13g2_fill_2 FILLER_59_2131 ();
 sg13g2_fill_2 FILLER_59_2137 ();
 sg13g2_fill_2 FILLER_59_2159 ();
 sg13g2_fill_1 FILLER_59_2161 ();
 sg13g2_fill_1 FILLER_59_2167 ();
 sg13g2_decap_8 FILLER_59_2194 ();
 sg13g2_decap_4 FILLER_59_2201 ();
 sg13g2_decap_4 FILLER_59_2210 ();
 sg13g2_fill_1 FILLER_59_2223 ();
 sg13g2_fill_2 FILLER_59_2233 ();
 sg13g2_fill_1 FILLER_59_2245 ();
 sg13g2_fill_2 FILLER_59_2254 ();
 sg13g2_fill_2 FILLER_59_2264 ();
 sg13g2_fill_1 FILLER_59_2266 ();
 sg13g2_fill_2 FILLER_59_2277 ();
 sg13g2_fill_1 FILLER_59_2279 ();
 sg13g2_decap_4 FILLER_59_2285 ();
 sg13g2_fill_1 FILLER_59_2289 ();
 sg13g2_decap_8 FILLER_59_2295 ();
 sg13g2_fill_1 FILLER_59_2302 ();
 sg13g2_decap_8 FILLER_59_2312 ();
 sg13g2_decap_8 FILLER_59_2322 ();
 sg13g2_decap_4 FILLER_59_2329 ();
 sg13g2_fill_1 FILLER_59_2337 ();
 sg13g2_decap_4 FILLER_59_2342 ();
 sg13g2_decap_8 FILLER_59_2350 ();
 sg13g2_decap_8 FILLER_59_2357 ();
 sg13g2_decap_8 FILLER_59_2364 ();
 sg13g2_decap_4 FILLER_59_2371 ();
 sg13g2_fill_2 FILLER_59_2375 ();
 sg13g2_decap_8 FILLER_59_2381 ();
 sg13g2_fill_2 FILLER_59_2417 ();
 sg13g2_fill_1 FILLER_59_2419 ();
 sg13g2_fill_2 FILLER_59_2440 ();
 sg13g2_fill_2 FILLER_59_2448 ();
 sg13g2_decap_8 FILLER_59_2493 ();
 sg13g2_fill_2 FILLER_59_2500 ();
 sg13g2_fill_1 FILLER_59_2508 ();
 sg13g2_fill_1 FILLER_59_2533 ();
 sg13g2_fill_2 FILLER_59_2540 ();
 sg13g2_fill_1 FILLER_59_2551 ();
 sg13g2_fill_2 FILLER_59_2556 ();
 sg13g2_fill_1 FILLER_59_2558 ();
 sg13g2_fill_1 FILLER_59_2596 ();
 sg13g2_decap_4 FILLER_59_2611 ();
 sg13g2_decap_4 FILLER_59_2638 ();
 sg13g2_decap_4 FILLER_59_2669 ();
 sg13g2_fill_1 FILLER_59_2673 ();
 sg13g2_fill_2 FILLER_59_2679 ();
 sg13g2_fill_2 FILLER_59_2685 ();
 sg13g2_fill_1 FILLER_59_2687 ();
 sg13g2_fill_1 FILLER_59_2699 ();
 sg13g2_fill_2 FILLER_59_2710 ();
 sg13g2_fill_2 FILLER_59_2716 ();
 sg13g2_fill_1 FILLER_59_2718 ();
 sg13g2_fill_1 FILLER_59_2724 ();
 sg13g2_fill_1 FILLER_59_2730 ();
 sg13g2_fill_2 FILLER_59_2743 ();
 sg13g2_fill_2 FILLER_59_2780 ();
 sg13g2_fill_1 FILLER_59_2782 ();
 sg13g2_fill_2 FILLER_59_2838 ();
 sg13g2_decap_4 FILLER_59_2852 ();
 sg13g2_fill_1 FILLER_59_2861 ();
 sg13g2_fill_1 FILLER_59_2878 ();
 sg13g2_decap_8 FILLER_59_2883 ();
 sg13g2_decap_8 FILLER_59_2890 ();
 sg13g2_decap_8 FILLER_59_2897 ();
 sg13g2_decap_4 FILLER_59_2932 ();
 sg13g2_fill_2 FILLER_59_2936 ();
 sg13g2_fill_2 FILLER_59_2943 ();
 sg13g2_fill_1 FILLER_59_2945 ();
 sg13g2_fill_2 FILLER_59_2954 ();
 sg13g2_fill_1 FILLER_59_2956 ();
 sg13g2_fill_2 FILLER_59_2963 ();
 sg13g2_decap_8 FILLER_59_3002 ();
 sg13g2_decap_8 FILLER_59_3009 ();
 sg13g2_decap_8 FILLER_59_3016 ();
 sg13g2_decap_8 FILLER_59_3023 ();
 sg13g2_decap_8 FILLER_59_3030 ();
 sg13g2_decap_8 FILLER_59_3037 ();
 sg13g2_decap_8 FILLER_59_3044 ();
 sg13g2_decap_8 FILLER_59_3051 ();
 sg13g2_decap_8 FILLER_59_3058 ();
 sg13g2_decap_8 FILLER_59_3065 ();
 sg13g2_decap_8 FILLER_59_3072 ();
 sg13g2_decap_8 FILLER_59_3079 ();
 sg13g2_decap_8 FILLER_59_3086 ();
 sg13g2_decap_8 FILLER_59_3093 ();
 sg13g2_decap_8 FILLER_59_3100 ();
 sg13g2_decap_8 FILLER_59_3107 ();
 sg13g2_decap_8 FILLER_59_3114 ();
 sg13g2_decap_8 FILLER_59_3121 ();
 sg13g2_decap_8 FILLER_59_3128 ();
 sg13g2_decap_8 FILLER_59_3135 ();
 sg13g2_decap_8 FILLER_59_3142 ();
 sg13g2_decap_8 FILLER_59_3149 ();
 sg13g2_decap_8 FILLER_59_3156 ();
 sg13g2_decap_8 FILLER_59_3163 ();
 sg13g2_decap_8 FILLER_59_3170 ();
 sg13g2_decap_8 FILLER_59_3177 ();
 sg13g2_decap_8 FILLER_59_3184 ();
 sg13g2_decap_8 FILLER_59_3191 ();
 sg13g2_decap_8 FILLER_59_3198 ();
 sg13g2_decap_8 FILLER_59_3205 ();
 sg13g2_decap_8 FILLER_59_3212 ();
 sg13g2_decap_8 FILLER_59_3219 ();
 sg13g2_decap_8 FILLER_59_3226 ();
 sg13g2_decap_8 FILLER_59_3233 ();
 sg13g2_decap_8 FILLER_59_3240 ();
 sg13g2_decap_8 FILLER_59_3247 ();
 sg13g2_decap_8 FILLER_59_3254 ();
 sg13g2_decap_8 FILLER_59_3261 ();
 sg13g2_decap_8 FILLER_59_3268 ();
 sg13g2_decap_8 FILLER_59_3275 ();
 sg13g2_decap_8 FILLER_59_3282 ();
 sg13g2_decap_8 FILLER_59_3289 ();
 sg13g2_decap_8 FILLER_59_3296 ();
 sg13g2_decap_8 FILLER_59_3303 ();
 sg13g2_decap_8 FILLER_59_3310 ();
 sg13g2_decap_8 FILLER_59_3317 ();
 sg13g2_decap_8 FILLER_59_3324 ();
 sg13g2_decap_8 FILLER_59_3331 ();
 sg13g2_decap_8 FILLER_59_3338 ();
 sg13g2_decap_8 FILLER_59_3345 ();
 sg13g2_decap_8 FILLER_59_3352 ();
 sg13g2_decap_8 FILLER_59_3359 ();
 sg13g2_decap_8 FILLER_59_3366 ();
 sg13g2_decap_8 FILLER_59_3373 ();
 sg13g2_decap_8 FILLER_59_3380 ();
 sg13g2_decap_8 FILLER_59_3387 ();
 sg13g2_decap_8 FILLER_59_3394 ();
 sg13g2_decap_8 FILLER_59_3401 ();
 sg13g2_decap_8 FILLER_59_3408 ();
 sg13g2_decap_8 FILLER_59_3415 ();
 sg13g2_decap_8 FILLER_59_3422 ();
 sg13g2_decap_8 FILLER_59_3429 ();
 sg13g2_decap_8 FILLER_59_3436 ();
 sg13g2_decap_8 FILLER_59_3443 ();
 sg13g2_decap_8 FILLER_59_3450 ();
 sg13g2_decap_8 FILLER_59_3457 ();
 sg13g2_decap_8 FILLER_59_3464 ();
 sg13g2_decap_8 FILLER_59_3471 ();
 sg13g2_decap_8 FILLER_59_3478 ();
 sg13g2_decap_8 FILLER_59_3485 ();
 sg13g2_decap_8 FILLER_59_3492 ();
 sg13g2_decap_8 FILLER_59_3499 ();
 sg13g2_decap_8 FILLER_59_3506 ();
 sg13g2_decap_8 FILLER_59_3513 ();
 sg13g2_decap_8 FILLER_59_3520 ();
 sg13g2_decap_8 FILLER_59_3527 ();
 sg13g2_decap_8 FILLER_59_3534 ();
 sg13g2_decap_8 FILLER_59_3541 ();
 sg13g2_decap_8 FILLER_59_3548 ();
 sg13g2_decap_8 FILLER_59_3555 ();
 sg13g2_decap_8 FILLER_59_3562 ();
 sg13g2_decap_8 FILLER_59_3569 ();
 sg13g2_decap_4 FILLER_59_3576 ();
 sg13g2_fill_2 FILLER_60_68 ();
 sg13g2_decap_4 FILLER_60_82 ();
 sg13g2_decap_8 FILLER_60_91 ();
 sg13g2_decap_4 FILLER_60_98 ();
 sg13g2_fill_1 FILLER_60_102 ();
 sg13g2_decap_8 FILLER_60_107 ();
 sg13g2_fill_2 FILLER_60_114 ();
 sg13g2_decap_8 FILLER_60_144 ();
 sg13g2_fill_1 FILLER_60_151 ();
 sg13g2_decap_8 FILLER_60_156 ();
 sg13g2_fill_1 FILLER_60_189 ();
 sg13g2_fill_2 FILLER_60_221 ();
 sg13g2_decap_8 FILLER_60_253 ();
 sg13g2_fill_1 FILLER_60_274 ();
 sg13g2_fill_2 FILLER_60_297 ();
 sg13g2_fill_2 FILLER_60_328 ();
 sg13g2_fill_1 FILLER_60_330 ();
 sg13g2_fill_2 FILLER_60_400 ();
 sg13g2_decap_4 FILLER_60_434 ();
 sg13g2_fill_2 FILLER_60_438 ();
 sg13g2_decap_8 FILLER_60_448 ();
 sg13g2_decap_4 FILLER_60_455 ();
 sg13g2_fill_2 FILLER_60_459 ();
 sg13g2_decap_4 FILLER_60_466 ();
 sg13g2_fill_2 FILLER_60_470 ();
 sg13g2_decap_4 FILLER_60_477 ();
 sg13g2_decap_8 FILLER_60_486 ();
 sg13g2_fill_2 FILLER_60_493 ();
 sg13g2_fill_1 FILLER_60_495 ();
 sg13g2_decap_4 FILLER_60_541 ();
 sg13g2_fill_2 FILLER_60_591 ();
 sg13g2_fill_1 FILLER_60_593 ();
 sg13g2_decap_4 FILLER_60_600 ();
 sg13g2_fill_2 FILLER_60_648 ();
 sg13g2_fill_2 FILLER_60_658 ();
 sg13g2_fill_2 FILLER_60_666 ();
 sg13g2_fill_2 FILLER_60_691 ();
 sg13g2_fill_1 FILLER_60_722 ();
 sg13g2_fill_1 FILLER_60_763 ();
 sg13g2_fill_2 FILLER_60_821 ();
 sg13g2_fill_1 FILLER_60_823 ();
 sg13g2_fill_2 FILLER_60_829 ();
 sg13g2_fill_1 FILLER_60_831 ();
 sg13g2_decap_8 FILLER_60_843 ();
 sg13g2_decap_4 FILLER_60_850 ();
 sg13g2_fill_1 FILLER_60_854 ();
 sg13g2_fill_2 FILLER_60_877 ();
 sg13g2_fill_1 FILLER_60_879 ();
 sg13g2_fill_1 FILLER_60_888 ();
 sg13g2_fill_2 FILLER_60_893 ();
 sg13g2_decap_8 FILLER_60_901 ();
 sg13g2_decap_8 FILLER_60_908 ();
 sg13g2_decap_4 FILLER_60_915 ();
 sg13g2_fill_1 FILLER_60_919 ();
 sg13g2_fill_2 FILLER_60_982 ();
 sg13g2_fill_1 FILLER_60_984 ();
 sg13g2_fill_1 FILLER_60_989 ();
 sg13g2_decap_4 FILLER_60_1000 ();
 sg13g2_fill_2 FILLER_60_1030 ();
 sg13g2_fill_1 FILLER_60_1042 ();
 sg13g2_fill_2 FILLER_60_1066 ();
 sg13g2_decap_8 FILLER_60_1076 ();
 sg13g2_decap_8 FILLER_60_1083 ();
 sg13g2_fill_1 FILLER_60_1096 ();
 sg13g2_decap_8 FILLER_60_1118 ();
 sg13g2_decap_8 FILLER_60_1125 ();
 sg13g2_fill_1 FILLER_60_1132 ();
 sg13g2_decap_4 FILLER_60_1174 ();
 sg13g2_fill_2 FILLER_60_1178 ();
 sg13g2_decap_4 FILLER_60_1188 ();
 sg13g2_fill_2 FILLER_60_1192 ();
 sg13g2_fill_1 FILLER_60_1220 ();
 sg13g2_fill_1 FILLER_60_1239 ();
 sg13g2_fill_2 FILLER_60_1253 ();
 sg13g2_fill_1 FILLER_60_1279 ();
 sg13g2_fill_2 FILLER_60_1320 ();
 sg13g2_fill_2 FILLER_60_1345 ();
 sg13g2_fill_1 FILLER_60_1352 ();
 sg13g2_decap_4 FILLER_60_1357 ();
 sg13g2_decap_4 FILLER_60_1373 ();
 sg13g2_fill_2 FILLER_60_1377 ();
 sg13g2_fill_2 FILLER_60_1392 ();
 sg13g2_fill_1 FILLER_60_1394 ();
 sg13g2_fill_1 FILLER_60_1400 ();
 sg13g2_decap_8 FILLER_60_1406 ();
 sg13g2_fill_2 FILLER_60_1413 ();
 sg13g2_decap_4 FILLER_60_1423 ();
 sg13g2_fill_1 FILLER_60_1427 ();
 sg13g2_fill_2 FILLER_60_1433 ();
 sg13g2_fill_1 FILLER_60_1435 ();
 sg13g2_fill_2 FILLER_60_1442 ();
 sg13g2_decap_8 FILLER_60_1449 ();
 sg13g2_decap_4 FILLER_60_1456 ();
 sg13g2_fill_2 FILLER_60_1491 ();
 sg13g2_fill_2 FILLER_60_1519 ();
 sg13g2_fill_1 FILLER_60_1521 ();
 sg13g2_fill_2 FILLER_60_1527 ();
 sg13g2_fill_1 FILLER_60_1529 ();
 sg13g2_fill_1 FILLER_60_1540 ();
 sg13g2_decap_8 FILLER_60_1586 ();
 sg13g2_fill_2 FILLER_60_1593 ();
 sg13g2_fill_1 FILLER_60_1595 ();
 sg13g2_fill_2 FILLER_60_1601 ();
 sg13g2_decap_8 FILLER_60_1607 ();
 sg13g2_decap_8 FILLER_60_1614 ();
 sg13g2_fill_2 FILLER_60_1621 ();
 sg13g2_fill_1 FILLER_60_1623 ();
 sg13g2_fill_2 FILLER_60_1663 ();
 sg13g2_decap_8 FILLER_60_1695 ();
 sg13g2_decap_4 FILLER_60_1714 ();
 sg13g2_decap_4 FILLER_60_1734 ();
 sg13g2_decap_4 FILLER_60_1759 ();
 sg13g2_fill_1 FILLER_60_1763 ();
 sg13g2_decap_8 FILLER_60_1772 ();
 sg13g2_fill_1 FILLER_60_1779 ();
 sg13g2_fill_2 FILLER_60_1801 ();
 sg13g2_fill_2 FILLER_60_1824 ();
 sg13g2_fill_1 FILLER_60_1826 ();
 sg13g2_fill_2 FILLER_60_1848 ();
 sg13g2_fill_1 FILLER_60_1850 ();
 sg13g2_fill_2 FILLER_60_1874 ();
 sg13g2_decap_8 FILLER_60_1902 ();
 sg13g2_decap_8 FILLER_60_1909 ();
 sg13g2_decap_4 FILLER_60_1916 ();
 sg13g2_fill_2 FILLER_60_1928 ();
 sg13g2_fill_1 FILLER_60_1930 ();
 sg13g2_fill_2 FILLER_60_1944 ();
 sg13g2_decap_8 FILLER_60_1959 ();
 sg13g2_fill_2 FILLER_60_1966 ();
 sg13g2_fill_2 FILLER_60_1984 ();
 sg13g2_fill_1 FILLER_60_1986 ();
 sg13g2_fill_2 FILLER_60_2003 ();
 sg13g2_decap_4 FILLER_60_2013 ();
 sg13g2_fill_2 FILLER_60_2017 ();
 sg13g2_decap_8 FILLER_60_2035 ();
 sg13g2_decap_8 FILLER_60_2042 ();
 sg13g2_fill_1 FILLER_60_2049 ();
 sg13g2_decap_8 FILLER_60_2054 ();
 sg13g2_fill_2 FILLER_60_2061 ();
 sg13g2_fill_2 FILLER_60_2081 ();
 sg13g2_decap_4 FILLER_60_2088 ();
 sg13g2_fill_1 FILLER_60_2092 ();
 sg13g2_decap_8 FILLER_60_2115 ();
 sg13g2_decap_8 FILLER_60_2122 ();
 sg13g2_decap_8 FILLER_60_2129 ();
 sg13g2_fill_1 FILLER_60_2136 ();
 sg13g2_decap_8 FILLER_60_2149 ();
 sg13g2_decap_8 FILLER_60_2156 ();
 sg13g2_decap_4 FILLER_60_2163 ();
 sg13g2_fill_2 FILLER_60_2167 ();
 sg13g2_fill_1 FILLER_60_2173 ();
 sg13g2_decap_4 FILLER_60_2189 ();
 sg13g2_fill_1 FILLER_60_2193 ();
 sg13g2_fill_2 FILLER_60_2236 ();
 sg13g2_decap_8 FILLER_60_2248 ();
 sg13g2_fill_1 FILLER_60_2272 ();
 sg13g2_decap_4 FILLER_60_2278 ();
 sg13g2_decap_4 FILLER_60_2292 ();
 sg13g2_fill_2 FILLER_60_2304 ();
 sg13g2_decap_4 FILLER_60_2322 ();
 sg13g2_fill_1 FILLER_60_2326 ();
 sg13g2_fill_2 FILLER_60_2385 ();
 sg13g2_fill_1 FILLER_60_2387 ();
 sg13g2_decap_8 FILLER_60_2434 ();
 sg13g2_fill_2 FILLER_60_2441 ();
 sg13g2_fill_1 FILLER_60_2443 ();
 sg13g2_decap_4 FILLER_60_2448 ();
 sg13g2_fill_2 FILLER_60_2465 ();
 sg13g2_decap_4 FILLER_60_2567 ();
 sg13g2_fill_1 FILLER_60_2571 ();
 sg13g2_decap_4 FILLER_60_2590 ();
 sg13g2_decap_4 FILLER_60_2604 ();
 sg13g2_fill_1 FILLER_60_2608 ();
 sg13g2_fill_1 FILLER_60_2626 ();
 sg13g2_decap_8 FILLER_60_2641 ();
 sg13g2_decap_4 FILLER_60_2648 ();
 sg13g2_fill_2 FILLER_60_2662 ();
 sg13g2_fill_1 FILLER_60_2664 ();
 sg13g2_fill_1 FILLER_60_2673 ();
 sg13g2_decap_8 FILLER_60_2682 ();
 sg13g2_decap_8 FILLER_60_2689 ();
 sg13g2_decap_8 FILLER_60_2706 ();
 sg13g2_decap_4 FILLER_60_2713 ();
 sg13g2_fill_1 FILLER_60_2717 ();
 sg13g2_decap_8 FILLER_60_2728 ();
 sg13g2_decap_8 FILLER_60_2735 ();
 sg13g2_fill_2 FILLER_60_2742 ();
 sg13g2_decap_4 FILLER_60_2754 ();
 sg13g2_fill_1 FILLER_60_2758 ();
 sg13g2_decap_8 FILLER_60_2774 ();
 sg13g2_decap_8 FILLER_60_2781 ();
 sg13g2_decap_8 FILLER_60_2788 ();
 sg13g2_decap_4 FILLER_60_2808 ();
 sg13g2_fill_1 FILLER_60_2812 ();
 sg13g2_fill_2 FILLER_60_2818 ();
 sg13g2_fill_2 FILLER_60_2825 ();
 sg13g2_fill_1 FILLER_60_2827 ();
 sg13g2_decap_8 FILLER_60_2838 ();
 sg13g2_fill_2 FILLER_60_2845 ();
 sg13g2_fill_1 FILLER_60_2860 ();
 sg13g2_fill_2 FILLER_60_2871 ();
 sg13g2_fill_1 FILLER_60_2873 ();
 sg13g2_decap_8 FILLER_60_2887 ();
 sg13g2_fill_1 FILLER_60_2894 ();
 sg13g2_fill_1 FILLER_60_2908 ();
 sg13g2_fill_1 FILLER_60_2914 ();
 sg13g2_fill_2 FILLER_60_2920 ();
 sg13g2_fill_2 FILLER_60_2926 ();
 sg13g2_decap_4 FILLER_60_2951 ();
 sg13g2_fill_1 FILLER_60_2955 ();
 sg13g2_decap_4 FILLER_60_2966 ();
 sg13g2_decap_8 FILLER_60_2992 ();
 sg13g2_decap_8 FILLER_60_2999 ();
 sg13g2_decap_8 FILLER_60_3006 ();
 sg13g2_decap_8 FILLER_60_3013 ();
 sg13g2_decap_8 FILLER_60_3020 ();
 sg13g2_decap_8 FILLER_60_3027 ();
 sg13g2_decap_8 FILLER_60_3034 ();
 sg13g2_decap_8 FILLER_60_3041 ();
 sg13g2_decap_8 FILLER_60_3048 ();
 sg13g2_decap_8 FILLER_60_3055 ();
 sg13g2_decap_8 FILLER_60_3062 ();
 sg13g2_decap_8 FILLER_60_3069 ();
 sg13g2_decap_8 FILLER_60_3076 ();
 sg13g2_decap_8 FILLER_60_3083 ();
 sg13g2_decap_8 FILLER_60_3090 ();
 sg13g2_decap_8 FILLER_60_3097 ();
 sg13g2_decap_8 FILLER_60_3104 ();
 sg13g2_decap_8 FILLER_60_3111 ();
 sg13g2_decap_8 FILLER_60_3118 ();
 sg13g2_decap_8 FILLER_60_3125 ();
 sg13g2_decap_8 FILLER_60_3132 ();
 sg13g2_decap_8 FILLER_60_3139 ();
 sg13g2_decap_8 FILLER_60_3146 ();
 sg13g2_decap_8 FILLER_60_3153 ();
 sg13g2_decap_8 FILLER_60_3160 ();
 sg13g2_decap_8 FILLER_60_3167 ();
 sg13g2_decap_8 FILLER_60_3174 ();
 sg13g2_decap_8 FILLER_60_3181 ();
 sg13g2_decap_8 FILLER_60_3188 ();
 sg13g2_decap_8 FILLER_60_3195 ();
 sg13g2_decap_8 FILLER_60_3202 ();
 sg13g2_decap_8 FILLER_60_3209 ();
 sg13g2_decap_8 FILLER_60_3216 ();
 sg13g2_decap_8 FILLER_60_3223 ();
 sg13g2_decap_8 FILLER_60_3230 ();
 sg13g2_decap_8 FILLER_60_3237 ();
 sg13g2_decap_8 FILLER_60_3244 ();
 sg13g2_decap_8 FILLER_60_3251 ();
 sg13g2_decap_8 FILLER_60_3258 ();
 sg13g2_decap_8 FILLER_60_3265 ();
 sg13g2_decap_8 FILLER_60_3272 ();
 sg13g2_decap_8 FILLER_60_3279 ();
 sg13g2_decap_8 FILLER_60_3286 ();
 sg13g2_decap_8 FILLER_60_3293 ();
 sg13g2_decap_8 FILLER_60_3300 ();
 sg13g2_decap_8 FILLER_60_3307 ();
 sg13g2_decap_8 FILLER_60_3314 ();
 sg13g2_decap_8 FILLER_60_3321 ();
 sg13g2_decap_8 FILLER_60_3328 ();
 sg13g2_decap_8 FILLER_60_3335 ();
 sg13g2_decap_8 FILLER_60_3342 ();
 sg13g2_decap_8 FILLER_60_3349 ();
 sg13g2_decap_8 FILLER_60_3356 ();
 sg13g2_decap_8 FILLER_60_3363 ();
 sg13g2_decap_8 FILLER_60_3370 ();
 sg13g2_decap_8 FILLER_60_3377 ();
 sg13g2_decap_8 FILLER_60_3384 ();
 sg13g2_decap_8 FILLER_60_3391 ();
 sg13g2_decap_8 FILLER_60_3398 ();
 sg13g2_decap_8 FILLER_60_3405 ();
 sg13g2_decap_8 FILLER_60_3412 ();
 sg13g2_decap_8 FILLER_60_3419 ();
 sg13g2_decap_8 FILLER_60_3426 ();
 sg13g2_decap_8 FILLER_60_3433 ();
 sg13g2_decap_8 FILLER_60_3440 ();
 sg13g2_decap_8 FILLER_60_3447 ();
 sg13g2_decap_8 FILLER_60_3454 ();
 sg13g2_decap_8 FILLER_60_3461 ();
 sg13g2_decap_8 FILLER_60_3468 ();
 sg13g2_decap_8 FILLER_60_3475 ();
 sg13g2_decap_8 FILLER_60_3482 ();
 sg13g2_decap_8 FILLER_60_3489 ();
 sg13g2_decap_8 FILLER_60_3496 ();
 sg13g2_decap_8 FILLER_60_3503 ();
 sg13g2_decap_8 FILLER_60_3510 ();
 sg13g2_decap_8 FILLER_60_3517 ();
 sg13g2_decap_8 FILLER_60_3524 ();
 sg13g2_decap_8 FILLER_60_3531 ();
 sg13g2_decap_8 FILLER_60_3538 ();
 sg13g2_decap_8 FILLER_60_3545 ();
 sg13g2_decap_8 FILLER_60_3552 ();
 sg13g2_decap_8 FILLER_60_3559 ();
 sg13g2_decap_8 FILLER_60_3566 ();
 sg13g2_decap_8 FILLER_60_3573 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_fill_2 FILLER_61_7 ();
 sg13g2_fill_1 FILLER_61_26 ();
 sg13g2_fill_2 FILLER_61_48 ();
 sg13g2_fill_1 FILLER_61_50 ();
 sg13g2_decap_8 FILLER_61_82 ();
 sg13g2_decap_8 FILLER_61_89 ();
 sg13g2_fill_1 FILLER_61_96 ();
 sg13g2_decap_8 FILLER_61_111 ();
 sg13g2_fill_2 FILLER_61_118 ();
 sg13g2_fill_1 FILLER_61_120 ();
 sg13g2_fill_2 FILLER_61_137 ();
 sg13g2_fill_1 FILLER_61_139 ();
 sg13g2_decap_8 FILLER_61_166 ();
 sg13g2_decap_8 FILLER_61_177 ();
 sg13g2_fill_2 FILLER_61_184 ();
 sg13g2_decap_8 FILLER_61_196 ();
 sg13g2_fill_2 FILLER_61_203 ();
 sg13g2_fill_1 FILLER_61_205 ();
 sg13g2_fill_2 FILLER_61_210 ();
 sg13g2_fill_2 FILLER_61_238 ();
 sg13g2_fill_1 FILLER_61_240 ();
 sg13g2_decap_4 FILLER_61_267 ();
 sg13g2_fill_1 FILLER_61_271 ();
 sg13g2_decap_8 FILLER_61_307 ();
 sg13g2_decap_4 FILLER_61_314 ();
 sg13g2_fill_2 FILLER_61_318 ();
 sg13g2_decap_8 FILLER_61_325 ();
 sg13g2_decap_8 FILLER_61_332 ();
 sg13g2_fill_2 FILLER_61_339 ();
 sg13g2_decap_8 FILLER_61_354 ();
 sg13g2_decap_8 FILLER_61_361 ();
 sg13g2_fill_2 FILLER_61_368 ();
 sg13g2_decap_8 FILLER_61_374 ();
 sg13g2_fill_2 FILLER_61_395 ();
 sg13g2_fill_1 FILLER_61_433 ();
 sg13g2_fill_2 FILLER_61_454 ();
 sg13g2_decap_4 FILLER_61_469 ();
 sg13g2_fill_2 FILLER_61_473 ();
 sg13g2_decap_8 FILLER_61_487 ();
 sg13g2_decap_4 FILLER_61_504 ();
 sg13g2_fill_1 FILLER_61_508 ();
 sg13g2_fill_2 FILLER_61_523 ();
 sg13g2_fill_2 FILLER_61_544 ();
 sg13g2_fill_1 FILLER_61_546 ();
 sg13g2_fill_1 FILLER_61_561 ();
 sg13g2_fill_2 FILLER_61_610 ();
 sg13g2_decap_4 FILLER_61_674 ();
 sg13g2_fill_1 FILLER_61_678 ();
 sg13g2_fill_2 FILLER_61_758 ();
 sg13g2_fill_1 FILLER_61_793 ();
 sg13g2_fill_2 FILLER_61_829 ();
 sg13g2_fill_1 FILLER_61_831 ();
 sg13g2_decap_8 FILLER_61_850 ();
 sg13g2_fill_1 FILLER_61_857 ();
 sg13g2_fill_2 FILLER_61_884 ();
 sg13g2_decap_4 FILLER_61_912 ();
 sg13g2_fill_1 FILLER_61_916 ();
 sg13g2_fill_1 FILLER_61_930 ();
 sg13g2_fill_1 FILLER_61_944 ();
 sg13g2_decap_4 FILLER_61_958 ();
 sg13g2_fill_1 FILLER_61_971 ();
 sg13g2_fill_2 FILLER_61_977 ();
 sg13g2_fill_1 FILLER_61_979 ();
 sg13g2_fill_2 FILLER_61_994 ();
 sg13g2_fill_1 FILLER_61_996 ();
 sg13g2_fill_2 FILLER_61_1005 ();
 sg13g2_fill_1 FILLER_61_1007 ();
 sg13g2_fill_2 FILLER_61_1022 ();
 sg13g2_decap_8 FILLER_61_1122 ();
 sg13g2_fill_1 FILLER_61_1134 ();
 sg13g2_decap_8 FILLER_61_1143 ();
 sg13g2_decap_8 FILLER_61_1150 ();
 sg13g2_fill_2 FILLER_61_1157 ();
 sg13g2_fill_2 FILLER_61_1164 ();
 sg13g2_fill_1 FILLER_61_1166 ();
 sg13g2_fill_1 FILLER_61_1171 ();
 sg13g2_decap_4 FILLER_61_1189 ();
 sg13g2_fill_1 FILLER_61_1193 ();
 sg13g2_fill_2 FILLER_61_1206 ();
 sg13g2_fill_2 FILLER_61_1217 ();
 sg13g2_fill_1 FILLER_61_1219 ();
 sg13g2_fill_1 FILLER_61_1248 ();
 sg13g2_decap_8 FILLER_61_1266 ();
 sg13g2_decap_8 FILLER_61_1273 ();
 sg13g2_fill_1 FILLER_61_1280 ();
 sg13g2_fill_1 FILLER_61_1290 ();
 sg13g2_fill_2 FILLER_61_1310 ();
 sg13g2_fill_2 FILLER_61_1355 ();
 sg13g2_fill_1 FILLER_61_1357 ();
 sg13g2_fill_2 FILLER_61_1376 ();
 sg13g2_fill_1 FILLER_61_1378 ();
 sg13g2_decap_8 FILLER_61_1387 ();
 sg13g2_fill_2 FILLER_61_1403 ();
 sg13g2_fill_2 FILLER_61_1442 ();
 sg13g2_fill_1 FILLER_61_1444 ();
 sg13g2_decap_8 FILLER_61_1453 ();
 sg13g2_decap_8 FILLER_61_1460 ();
 sg13g2_decap_8 FILLER_61_1467 ();
 sg13g2_decap_4 FILLER_61_1474 ();
 sg13g2_fill_2 FILLER_61_1486 ();
 sg13g2_fill_2 FILLER_61_1502 ();
 sg13g2_decap_8 FILLER_61_1508 ();
 sg13g2_decap_4 FILLER_61_1515 ();
 sg13g2_fill_1 FILLER_61_1519 ();
 sg13g2_fill_2 FILLER_61_1561 ();
 sg13g2_fill_1 FILLER_61_1563 ();
 sg13g2_fill_1 FILLER_61_1604 ();
 sg13g2_fill_2 FILLER_61_1618 ();
 sg13g2_fill_2 FILLER_61_1626 ();
 sg13g2_decap_8 FILLER_61_1636 ();
 sg13g2_decap_8 FILLER_61_1647 ();
 sg13g2_decap_8 FILLER_61_1654 ();
 sg13g2_decap_8 FILLER_61_1671 ();
 sg13g2_decap_8 FILLER_61_1678 ();
 sg13g2_decap_8 FILLER_61_1685 ();
 sg13g2_decap_4 FILLER_61_1692 ();
 sg13g2_fill_1 FILLER_61_1701 ();
 sg13g2_decap_4 FILLER_61_1714 ();
 sg13g2_decap_4 FILLER_61_1723 ();
 sg13g2_decap_4 FILLER_61_1732 ();
 sg13g2_fill_2 FILLER_61_1736 ();
 sg13g2_decap_8 FILLER_61_1751 ();
 sg13g2_fill_2 FILLER_61_1758 ();
 sg13g2_fill_1 FILLER_61_1760 ();
 sg13g2_fill_1 FILLER_61_1771 ();
 sg13g2_fill_2 FILLER_61_1785 ();
 sg13g2_fill_1 FILLER_61_1787 ();
 sg13g2_fill_2 FILLER_61_1801 ();
 sg13g2_fill_2 FILLER_61_1807 ();
 sg13g2_fill_1 FILLER_61_1809 ();
 sg13g2_decap_4 FILLER_61_1818 ();
 sg13g2_decap_4 FILLER_61_1843 ();
 sg13g2_fill_1 FILLER_61_1847 ();
 sg13g2_decap_4 FILLER_61_1872 ();
 sg13g2_fill_1 FILLER_61_1876 ();
 sg13g2_decap_8 FILLER_61_1894 ();
 sg13g2_fill_1 FILLER_61_1901 ();
 sg13g2_decap_8 FILLER_61_1906 ();
 sg13g2_fill_2 FILLER_61_1913 ();
 sg13g2_fill_1 FILLER_61_1915 ();
 sg13g2_decap_4 FILLER_61_1924 ();
 sg13g2_fill_2 FILLER_61_1936 ();
 sg13g2_fill_1 FILLER_61_1955 ();
 sg13g2_fill_2 FILLER_61_1969 ();
 sg13g2_fill_1 FILLER_61_1975 ();
 sg13g2_decap_8 FILLER_61_1993 ();
 sg13g2_fill_2 FILLER_61_2000 ();
 sg13g2_fill_1 FILLER_61_2002 ();
 sg13g2_decap_8 FILLER_61_2011 ();
 sg13g2_decap_4 FILLER_61_2018 ();
 sg13g2_fill_1 FILLER_61_2022 ();
 sg13g2_decap_8 FILLER_61_2043 ();
 sg13g2_decap_8 FILLER_61_2050 ();
 sg13g2_decap_4 FILLER_61_2057 ();
 sg13g2_fill_1 FILLER_61_2061 ();
 sg13g2_decap_8 FILLER_61_2069 ();
 sg13g2_fill_2 FILLER_61_2076 ();
 sg13g2_fill_1 FILLER_61_2078 ();
 sg13g2_fill_2 FILLER_61_2103 ();
 sg13g2_decap_8 FILLER_61_2122 ();
 sg13g2_fill_1 FILLER_61_2129 ();
 sg13g2_fill_2 FILLER_61_2134 ();
 sg13g2_fill_2 FILLER_61_2140 ();
 sg13g2_decap_4 FILLER_61_2157 ();
 sg13g2_fill_1 FILLER_61_2174 ();
 sg13g2_decap_4 FILLER_61_2188 ();
 sg13g2_fill_1 FILLER_61_2192 ();
 sg13g2_fill_1 FILLER_61_2206 ();
 sg13g2_decap_8 FILLER_61_2215 ();
 sg13g2_decap_4 FILLER_61_2231 ();
 sg13g2_fill_2 FILLER_61_2235 ();
 sg13g2_fill_2 FILLER_61_2241 ();
 sg13g2_fill_1 FILLER_61_2243 ();
 sg13g2_fill_1 FILLER_61_2259 ();
 sg13g2_decap_8 FILLER_61_2270 ();
 sg13g2_decap_8 FILLER_61_2277 ();
 sg13g2_decap_8 FILLER_61_2284 ();
 sg13g2_fill_2 FILLER_61_2291 ();
 sg13g2_decap_8 FILLER_61_2313 ();
 sg13g2_decap_8 FILLER_61_2320 ();
 sg13g2_fill_2 FILLER_61_2340 ();
 sg13g2_fill_1 FILLER_61_2342 ();
 sg13g2_fill_1 FILLER_61_2352 ();
 sg13g2_fill_2 FILLER_61_2373 ();
 sg13g2_fill_1 FILLER_61_2375 ();
 sg13g2_fill_1 FILLER_61_2395 ();
 sg13g2_fill_1 FILLER_61_2409 ();
 sg13g2_fill_2 FILLER_61_2436 ();
 sg13g2_fill_2 FILLER_61_2442 ();
 sg13g2_fill_1 FILLER_61_2444 ();
 sg13g2_fill_1 FILLER_61_2449 ();
 sg13g2_fill_2 FILLER_61_2488 ();
 sg13g2_decap_8 FILLER_61_2499 ();
 sg13g2_fill_2 FILLER_61_2506 ();
 sg13g2_fill_1 FILLER_61_2515 ();
 sg13g2_fill_2 FILLER_61_2532 ();
 sg13g2_decap_8 FILLER_61_2565 ();
 sg13g2_decap_8 FILLER_61_2572 ();
 sg13g2_fill_1 FILLER_61_2579 ();
 sg13g2_decap_8 FILLER_61_2600 ();
 sg13g2_fill_1 FILLER_61_2607 ();
 sg13g2_fill_1 FILLER_61_2622 ();
 sg13g2_decap_8 FILLER_61_2637 ();
 sg13g2_fill_2 FILLER_61_2644 ();
 sg13g2_fill_1 FILLER_61_2673 ();
 sg13g2_decap_8 FILLER_61_2684 ();
 sg13g2_fill_2 FILLER_61_2691 ();
 sg13g2_fill_2 FILLER_61_2697 ();
 sg13g2_fill_1 FILLER_61_2699 ();
 sg13g2_fill_1 FILLER_61_2709 ();
 sg13g2_decap_4 FILLER_61_2754 ();
 sg13g2_fill_2 FILLER_61_2758 ();
 sg13g2_decap_8 FILLER_61_2771 ();
 sg13g2_decap_8 FILLER_61_2778 ();
 sg13g2_fill_1 FILLER_61_2785 ();
 sg13g2_fill_1 FILLER_61_2791 ();
 sg13g2_decap_8 FILLER_61_2805 ();
 sg13g2_decap_8 FILLER_61_2812 ();
 sg13g2_decap_4 FILLER_61_2819 ();
 sg13g2_decap_8 FILLER_61_2833 ();
 sg13g2_decap_8 FILLER_61_2840 ();
 sg13g2_fill_1 FILLER_61_2847 ();
 sg13g2_fill_1 FILLER_61_2868 ();
 sg13g2_decap_8 FILLER_61_2874 ();
 sg13g2_decap_8 FILLER_61_2881 ();
 sg13g2_decap_8 FILLER_61_2888 ();
 sg13g2_decap_4 FILLER_61_2895 ();
 sg13g2_decap_4 FILLER_61_2952 ();
 sg13g2_fill_1 FILLER_61_2974 ();
 sg13g2_decap_8 FILLER_61_3001 ();
 sg13g2_decap_8 FILLER_61_3008 ();
 sg13g2_decap_8 FILLER_61_3015 ();
 sg13g2_decap_8 FILLER_61_3022 ();
 sg13g2_decap_8 FILLER_61_3029 ();
 sg13g2_decap_8 FILLER_61_3036 ();
 sg13g2_decap_8 FILLER_61_3043 ();
 sg13g2_decap_8 FILLER_61_3050 ();
 sg13g2_decap_8 FILLER_61_3057 ();
 sg13g2_decap_8 FILLER_61_3064 ();
 sg13g2_decap_8 FILLER_61_3071 ();
 sg13g2_decap_8 FILLER_61_3078 ();
 sg13g2_decap_8 FILLER_61_3085 ();
 sg13g2_decap_8 FILLER_61_3092 ();
 sg13g2_decap_8 FILLER_61_3099 ();
 sg13g2_decap_8 FILLER_61_3106 ();
 sg13g2_decap_8 FILLER_61_3113 ();
 sg13g2_decap_8 FILLER_61_3120 ();
 sg13g2_decap_8 FILLER_61_3127 ();
 sg13g2_decap_8 FILLER_61_3134 ();
 sg13g2_decap_8 FILLER_61_3141 ();
 sg13g2_decap_8 FILLER_61_3148 ();
 sg13g2_decap_8 FILLER_61_3155 ();
 sg13g2_decap_8 FILLER_61_3162 ();
 sg13g2_decap_8 FILLER_61_3169 ();
 sg13g2_decap_8 FILLER_61_3176 ();
 sg13g2_decap_8 FILLER_61_3183 ();
 sg13g2_decap_8 FILLER_61_3190 ();
 sg13g2_decap_8 FILLER_61_3197 ();
 sg13g2_decap_8 FILLER_61_3204 ();
 sg13g2_decap_8 FILLER_61_3211 ();
 sg13g2_decap_8 FILLER_61_3218 ();
 sg13g2_decap_8 FILLER_61_3225 ();
 sg13g2_decap_8 FILLER_61_3232 ();
 sg13g2_decap_8 FILLER_61_3239 ();
 sg13g2_decap_8 FILLER_61_3246 ();
 sg13g2_decap_8 FILLER_61_3253 ();
 sg13g2_decap_8 FILLER_61_3260 ();
 sg13g2_decap_8 FILLER_61_3267 ();
 sg13g2_decap_8 FILLER_61_3274 ();
 sg13g2_decap_8 FILLER_61_3281 ();
 sg13g2_decap_8 FILLER_61_3288 ();
 sg13g2_decap_8 FILLER_61_3295 ();
 sg13g2_decap_8 FILLER_61_3302 ();
 sg13g2_decap_8 FILLER_61_3309 ();
 sg13g2_decap_8 FILLER_61_3316 ();
 sg13g2_decap_8 FILLER_61_3323 ();
 sg13g2_decap_8 FILLER_61_3330 ();
 sg13g2_decap_8 FILLER_61_3337 ();
 sg13g2_decap_8 FILLER_61_3344 ();
 sg13g2_decap_8 FILLER_61_3351 ();
 sg13g2_decap_8 FILLER_61_3358 ();
 sg13g2_decap_8 FILLER_61_3365 ();
 sg13g2_decap_8 FILLER_61_3372 ();
 sg13g2_decap_8 FILLER_61_3379 ();
 sg13g2_decap_8 FILLER_61_3386 ();
 sg13g2_decap_8 FILLER_61_3393 ();
 sg13g2_decap_8 FILLER_61_3400 ();
 sg13g2_decap_8 FILLER_61_3407 ();
 sg13g2_decap_8 FILLER_61_3414 ();
 sg13g2_decap_8 FILLER_61_3421 ();
 sg13g2_decap_8 FILLER_61_3428 ();
 sg13g2_decap_8 FILLER_61_3435 ();
 sg13g2_decap_8 FILLER_61_3442 ();
 sg13g2_decap_8 FILLER_61_3449 ();
 sg13g2_decap_8 FILLER_61_3456 ();
 sg13g2_decap_8 FILLER_61_3463 ();
 sg13g2_decap_8 FILLER_61_3470 ();
 sg13g2_decap_8 FILLER_61_3477 ();
 sg13g2_decap_8 FILLER_61_3484 ();
 sg13g2_decap_8 FILLER_61_3491 ();
 sg13g2_decap_8 FILLER_61_3498 ();
 sg13g2_decap_8 FILLER_61_3505 ();
 sg13g2_decap_8 FILLER_61_3512 ();
 sg13g2_decap_8 FILLER_61_3519 ();
 sg13g2_decap_8 FILLER_61_3526 ();
 sg13g2_decap_8 FILLER_61_3533 ();
 sg13g2_decap_8 FILLER_61_3540 ();
 sg13g2_decap_8 FILLER_61_3547 ();
 sg13g2_decap_8 FILLER_61_3554 ();
 sg13g2_decap_8 FILLER_61_3561 ();
 sg13g2_decap_8 FILLER_61_3568 ();
 sg13g2_decap_4 FILLER_61_3575 ();
 sg13g2_fill_1 FILLER_61_3579 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_7 ();
 sg13g2_fill_1 FILLER_62_11 ();
 sg13g2_decap_8 FILLER_62_16 ();
 sg13g2_fill_1 FILLER_62_73 ();
 sg13g2_fill_2 FILLER_62_95 ();
 sg13g2_fill_1 FILLER_62_97 ();
 sg13g2_fill_1 FILLER_62_106 ();
 sg13g2_fill_2 FILLER_62_117 ();
 sg13g2_fill_1 FILLER_62_119 ();
 sg13g2_fill_1 FILLER_62_138 ();
 sg13g2_fill_1 FILLER_62_148 ();
 sg13g2_fill_2 FILLER_62_190 ();
 sg13g2_fill_1 FILLER_62_192 ();
 sg13g2_fill_1 FILLER_62_198 ();
 sg13g2_fill_1 FILLER_62_204 ();
 sg13g2_decap_8 FILLER_62_231 ();
 sg13g2_decap_4 FILLER_62_238 ();
 sg13g2_fill_2 FILLER_62_242 ();
 sg13g2_decap_4 FILLER_62_248 ();
 sg13g2_decap_8 FILLER_62_256 ();
 sg13g2_fill_1 FILLER_62_263 ();
 sg13g2_decap_8 FILLER_62_274 ();
 sg13g2_fill_1 FILLER_62_286 ();
 sg13g2_decap_8 FILLER_62_296 ();
 sg13g2_fill_1 FILLER_62_303 ();
 sg13g2_fill_1 FILLER_62_335 ();
 sg13g2_fill_1 FILLER_62_373 ();
 sg13g2_decap_8 FILLER_62_395 ();
 sg13g2_fill_2 FILLER_62_402 ();
 sg13g2_decap_8 FILLER_62_433 ();
 sg13g2_fill_2 FILLER_62_440 ();
 sg13g2_fill_1 FILLER_62_448 ();
 sg13g2_fill_2 FILLER_62_461 ();
 sg13g2_fill_1 FILLER_62_463 ();
 sg13g2_fill_1 FILLER_62_499 ();
 sg13g2_decap_4 FILLER_62_510 ();
 sg13g2_decap_4 FILLER_62_526 ();
 sg13g2_fill_1 FILLER_62_579 ();
 sg13g2_decap_8 FILLER_62_589 ();
 sg13g2_fill_1 FILLER_62_596 ();
 sg13g2_decap_4 FILLER_62_607 ();
 sg13g2_fill_1 FILLER_62_611 ();
 sg13g2_fill_2 FILLER_62_619 ();
 sg13g2_fill_1 FILLER_62_621 ();
 sg13g2_fill_2 FILLER_62_627 ();
 sg13g2_fill_2 FILLER_62_633 ();
 sg13g2_fill_2 FILLER_62_663 ();
 sg13g2_fill_1 FILLER_62_746 ();
 sg13g2_fill_1 FILLER_62_803 ();
 sg13g2_fill_1 FILLER_62_808 ();
 sg13g2_decap_4 FILLER_62_824 ();
 sg13g2_fill_2 FILLER_62_828 ();
 sg13g2_fill_2 FILLER_62_835 ();
 sg13g2_fill_1 FILLER_62_837 ();
 sg13g2_decap_4 FILLER_62_851 ();
 sg13g2_fill_1 FILLER_62_869 ();
 sg13g2_fill_2 FILLER_62_887 ();
 sg13g2_fill_2 FILLER_62_920 ();
 sg13g2_fill_1 FILLER_62_922 ();
 sg13g2_fill_2 FILLER_62_949 ();
 sg13g2_fill_2 FILLER_62_956 ();
 sg13g2_fill_1 FILLER_62_958 ();
 sg13g2_fill_2 FILLER_62_1065 ();
 sg13g2_fill_1 FILLER_62_1067 ();
 sg13g2_decap_4 FILLER_62_1115 ();
 sg13g2_fill_1 FILLER_62_1119 ();
 sg13g2_fill_1 FILLER_62_1150 ();
 sg13g2_fill_2 FILLER_62_1188 ();
 sg13g2_fill_1 FILLER_62_1190 ();
 sg13g2_fill_2 FILLER_62_1217 ();
 sg13g2_fill_1 FILLER_62_1219 ();
 sg13g2_fill_2 FILLER_62_1225 ();
 sg13g2_fill_1 FILLER_62_1227 ();
 sg13g2_fill_1 FILLER_62_1238 ();
 sg13g2_decap_4 FILLER_62_1244 ();
 sg13g2_fill_1 FILLER_62_1248 ();
 sg13g2_fill_2 FILLER_62_1289 ();
 sg13g2_fill_1 FILLER_62_1291 ();
 sg13g2_decap_4 FILLER_62_1300 ();
 sg13g2_decap_4 FILLER_62_1336 ();
 sg13g2_decap_8 FILLER_62_1344 ();
 sg13g2_decap_8 FILLER_62_1351 ();
 sg13g2_fill_2 FILLER_62_1358 ();
 sg13g2_decap_8 FILLER_62_1365 ();
 sg13g2_decap_4 FILLER_62_1372 ();
 sg13g2_decap_8 FILLER_62_1420 ();
 sg13g2_fill_2 FILLER_62_1431 ();
 sg13g2_fill_1 FILLER_62_1433 ();
 sg13g2_decap_4 FILLER_62_1460 ();
 sg13g2_fill_1 FILLER_62_1464 ();
 sg13g2_fill_2 FILLER_62_1486 ();
 sg13g2_fill_1 FILLER_62_1488 ();
 sg13g2_decap_8 FILLER_62_1504 ();
 sg13g2_fill_2 FILLER_62_1511 ();
 sg13g2_fill_1 FILLER_62_1513 ();
 sg13g2_fill_2 FILLER_62_1526 ();
 sg13g2_fill_1 FILLER_62_1528 ();
 sg13g2_fill_2 FILLER_62_1534 ();
 sg13g2_decap_4 FILLER_62_1548 ();
 sg13g2_fill_2 FILLER_62_1552 ();
 sg13g2_fill_2 FILLER_62_1572 ();
 sg13g2_fill_1 FILLER_62_1588 ();
 sg13g2_decap_4 FILLER_62_1597 ();
 sg13g2_fill_2 FILLER_62_1601 ();
 sg13g2_decap_4 FILLER_62_1608 ();
 sg13g2_fill_1 FILLER_62_1612 ();
 sg13g2_decap_8 FILLER_62_1639 ();
 sg13g2_decap_8 FILLER_62_1646 ();
 sg13g2_fill_1 FILLER_62_1653 ();
 sg13g2_fill_2 FILLER_62_1658 ();
 sg13g2_fill_1 FILLER_62_1660 ();
 sg13g2_fill_2 FILLER_62_1666 ();
 sg13g2_fill_1 FILLER_62_1673 ();
 sg13g2_decap_8 FILLER_62_1716 ();
 sg13g2_fill_1 FILLER_62_1723 ();
 sg13g2_decap_8 FILLER_62_1737 ();
 sg13g2_fill_2 FILLER_62_1744 ();
 sg13g2_decap_4 FILLER_62_1751 ();
 sg13g2_fill_2 FILLER_62_1755 ();
 sg13g2_fill_2 FILLER_62_1765 ();
 sg13g2_decap_4 FILLER_62_1780 ();
 sg13g2_fill_1 FILLER_62_1784 ();
 sg13g2_decap_4 FILLER_62_1796 ();
 sg13g2_fill_1 FILLER_62_1800 ();
 sg13g2_decap_8 FILLER_62_1805 ();
 sg13g2_decap_8 FILLER_62_1812 ();
 sg13g2_decap_8 FILLER_62_1819 ();
 sg13g2_decap_4 FILLER_62_1826 ();
 sg13g2_fill_2 FILLER_62_1830 ();
 sg13g2_decap_8 FILLER_62_1836 ();
 sg13g2_fill_1 FILLER_62_1843 ();
 sg13g2_decap_8 FILLER_62_1870 ();
 sg13g2_decap_8 FILLER_62_1877 ();
 sg13g2_decap_8 FILLER_62_1884 ();
 sg13g2_decap_8 FILLER_62_1917 ();
 sg13g2_decap_8 FILLER_62_1924 ();
 sg13g2_decap_4 FILLER_62_1931 ();
 sg13g2_fill_2 FILLER_62_1935 ();
 sg13g2_decap_8 FILLER_62_1957 ();
 sg13g2_decap_8 FILLER_62_1964 ();
 sg13g2_decap_4 FILLER_62_1971 ();
 sg13g2_decap_8 FILLER_62_1991 ();
 sg13g2_decap_8 FILLER_62_1998 ();
 sg13g2_decap_4 FILLER_62_2018 ();
 sg13g2_fill_2 FILLER_62_2053 ();
 sg13g2_fill_1 FILLER_62_2063 ();
 sg13g2_decap_8 FILLER_62_2072 ();
 sg13g2_fill_2 FILLER_62_2079 ();
 sg13g2_decap_8 FILLER_62_2094 ();
 sg13g2_fill_1 FILLER_62_2101 ();
 sg13g2_decap_8 FILLER_62_2110 ();
 sg13g2_decap_8 FILLER_62_2117 ();
 sg13g2_decap_8 FILLER_62_2124 ();
 sg13g2_fill_1 FILLER_62_2131 ();
 sg13g2_fill_2 FILLER_62_2141 ();
 sg13g2_fill_1 FILLER_62_2143 ();
 sg13g2_decap_8 FILLER_62_2159 ();
 sg13g2_decap_4 FILLER_62_2166 ();
 sg13g2_fill_2 FILLER_62_2170 ();
 sg13g2_fill_1 FILLER_62_2181 ();
 sg13g2_decap_4 FILLER_62_2191 ();
 sg13g2_fill_1 FILLER_62_2195 ();
 sg13g2_fill_2 FILLER_62_2211 ();
 sg13g2_fill_1 FILLER_62_2213 ();
 sg13g2_fill_2 FILLER_62_2218 ();
 sg13g2_fill_1 FILLER_62_2220 ();
 sg13g2_decap_8 FILLER_62_2237 ();
 sg13g2_fill_2 FILLER_62_2244 ();
 sg13g2_fill_1 FILLER_62_2246 ();
 sg13g2_decap_8 FILLER_62_2260 ();
 sg13g2_decap_8 FILLER_62_2267 ();
 sg13g2_fill_2 FILLER_62_2274 ();
 sg13g2_fill_1 FILLER_62_2276 ();
 sg13g2_fill_1 FILLER_62_2295 ();
 sg13g2_fill_1 FILLER_62_2309 ();
 sg13g2_fill_1 FILLER_62_2319 ();
 sg13g2_fill_2 FILLER_62_2365 ();
 sg13g2_fill_2 FILLER_62_2376 ();
 sg13g2_fill_2 FILLER_62_2404 ();
 sg13g2_fill_2 FILLER_62_2465 ();
 sg13g2_decap_8 FILLER_62_2508 ();
 sg13g2_fill_2 FILLER_62_2515 ();
 sg13g2_fill_2 FILLER_62_2530 ();
 sg13g2_decap_8 FILLER_62_2573 ();
 sg13g2_decap_8 FILLER_62_2600 ();
 sg13g2_fill_1 FILLER_62_2607 ();
 sg13g2_decap_4 FILLER_62_2631 ();
 sg13g2_fill_2 FILLER_62_2635 ();
 sg13g2_decap_8 FILLER_62_2671 ();
 sg13g2_fill_2 FILLER_62_2678 ();
 sg13g2_fill_1 FILLER_62_2680 ();
 sg13g2_fill_2 FILLER_62_2693 ();
 sg13g2_fill_1 FILLER_62_2707 ();
 sg13g2_fill_2 FILLER_62_2713 ();
 sg13g2_fill_1 FILLER_62_2715 ();
 sg13g2_fill_1 FILLER_62_2725 ();
 sg13g2_decap_8 FILLER_62_2734 ();
 sg13g2_decap_8 FILLER_62_2754 ();
 sg13g2_decap_4 FILLER_62_2761 ();
 sg13g2_fill_1 FILLER_62_2765 ();
 sg13g2_fill_2 FILLER_62_2782 ();
 sg13g2_fill_1 FILLER_62_2801 ();
 sg13g2_fill_1 FILLER_62_2815 ();
 sg13g2_fill_2 FILLER_62_2819 ();
 sg13g2_fill_1 FILLER_62_2826 ();
 sg13g2_fill_2 FILLER_62_2852 ();
 sg13g2_fill_1 FILLER_62_2854 ();
 sg13g2_fill_2 FILLER_62_2895 ();
 sg13g2_fill_2 FILLER_62_2907 ();
 sg13g2_fill_1 FILLER_62_2909 ();
 sg13g2_decap_8 FILLER_62_2915 ();
 sg13g2_decap_8 FILLER_62_2922 ();
 sg13g2_fill_1 FILLER_62_2929 ();
 sg13g2_decap_8 FILLER_62_2935 ();
 sg13g2_decap_8 FILLER_62_2942 ();
 sg13g2_fill_1 FILLER_62_2949 ();
 sg13g2_fill_2 FILLER_62_2967 ();
 sg13g2_fill_1 FILLER_62_2969 ();
 sg13g2_decap_8 FILLER_62_2977 ();
 sg13g2_fill_2 FILLER_62_2984 ();
 sg13g2_decap_8 FILLER_62_2999 ();
 sg13g2_decap_8 FILLER_62_3006 ();
 sg13g2_decap_8 FILLER_62_3013 ();
 sg13g2_decap_8 FILLER_62_3020 ();
 sg13g2_decap_8 FILLER_62_3027 ();
 sg13g2_decap_8 FILLER_62_3034 ();
 sg13g2_decap_8 FILLER_62_3041 ();
 sg13g2_decap_8 FILLER_62_3048 ();
 sg13g2_decap_8 FILLER_62_3055 ();
 sg13g2_decap_8 FILLER_62_3062 ();
 sg13g2_decap_8 FILLER_62_3069 ();
 sg13g2_decap_8 FILLER_62_3076 ();
 sg13g2_decap_8 FILLER_62_3083 ();
 sg13g2_decap_8 FILLER_62_3090 ();
 sg13g2_decap_8 FILLER_62_3097 ();
 sg13g2_decap_8 FILLER_62_3104 ();
 sg13g2_decap_8 FILLER_62_3111 ();
 sg13g2_decap_8 FILLER_62_3118 ();
 sg13g2_decap_8 FILLER_62_3125 ();
 sg13g2_decap_8 FILLER_62_3132 ();
 sg13g2_decap_8 FILLER_62_3139 ();
 sg13g2_decap_8 FILLER_62_3146 ();
 sg13g2_decap_8 FILLER_62_3153 ();
 sg13g2_decap_8 FILLER_62_3160 ();
 sg13g2_decap_8 FILLER_62_3167 ();
 sg13g2_decap_8 FILLER_62_3174 ();
 sg13g2_decap_8 FILLER_62_3181 ();
 sg13g2_decap_8 FILLER_62_3188 ();
 sg13g2_decap_8 FILLER_62_3195 ();
 sg13g2_decap_8 FILLER_62_3202 ();
 sg13g2_decap_8 FILLER_62_3209 ();
 sg13g2_decap_8 FILLER_62_3216 ();
 sg13g2_decap_8 FILLER_62_3223 ();
 sg13g2_decap_8 FILLER_62_3230 ();
 sg13g2_decap_8 FILLER_62_3237 ();
 sg13g2_decap_8 FILLER_62_3244 ();
 sg13g2_decap_8 FILLER_62_3251 ();
 sg13g2_decap_8 FILLER_62_3258 ();
 sg13g2_decap_8 FILLER_62_3265 ();
 sg13g2_decap_8 FILLER_62_3272 ();
 sg13g2_decap_8 FILLER_62_3279 ();
 sg13g2_decap_8 FILLER_62_3286 ();
 sg13g2_decap_8 FILLER_62_3293 ();
 sg13g2_decap_8 FILLER_62_3300 ();
 sg13g2_decap_8 FILLER_62_3307 ();
 sg13g2_decap_8 FILLER_62_3314 ();
 sg13g2_decap_8 FILLER_62_3321 ();
 sg13g2_decap_8 FILLER_62_3328 ();
 sg13g2_decap_8 FILLER_62_3335 ();
 sg13g2_decap_8 FILLER_62_3342 ();
 sg13g2_decap_8 FILLER_62_3349 ();
 sg13g2_decap_8 FILLER_62_3356 ();
 sg13g2_decap_8 FILLER_62_3363 ();
 sg13g2_decap_8 FILLER_62_3370 ();
 sg13g2_decap_8 FILLER_62_3377 ();
 sg13g2_decap_8 FILLER_62_3384 ();
 sg13g2_decap_8 FILLER_62_3391 ();
 sg13g2_decap_8 FILLER_62_3398 ();
 sg13g2_decap_8 FILLER_62_3405 ();
 sg13g2_decap_8 FILLER_62_3412 ();
 sg13g2_decap_8 FILLER_62_3419 ();
 sg13g2_decap_8 FILLER_62_3426 ();
 sg13g2_decap_8 FILLER_62_3433 ();
 sg13g2_decap_8 FILLER_62_3440 ();
 sg13g2_decap_8 FILLER_62_3447 ();
 sg13g2_decap_8 FILLER_62_3454 ();
 sg13g2_decap_8 FILLER_62_3461 ();
 sg13g2_decap_8 FILLER_62_3468 ();
 sg13g2_decap_8 FILLER_62_3475 ();
 sg13g2_decap_8 FILLER_62_3482 ();
 sg13g2_decap_8 FILLER_62_3489 ();
 sg13g2_decap_8 FILLER_62_3496 ();
 sg13g2_decap_8 FILLER_62_3503 ();
 sg13g2_decap_8 FILLER_62_3510 ();
 sg13g2_decap_8 FILLER_62_3517 ();
 sg13g2_decap_8 FILLER_62_3524 ();
 sg13g2_decap_8 FILLER_62_3531 ();
 sg13g2_decap_8 FILLER_62_3538 ();
 sg13g2_decap_8 FILLER_62_3545 ();
 sg13g2_decap_8 FILLER_62_3552 ();
 sg13g2_decap_8 FILLER_62_3559 ();
 sg13g2_decap_8 FILLER_62_3566 ();
 sg13g2_decap_8 FILLER_62_3573 ();
 sg13g2_fill_1 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_27 ();
 sg13g2_fill_1 FILLER_63_83 ();
 sg13g2_decap_4 FILLER_63_96 ();
 sg13g2_decap_4 FILLER_63_105 ();
 sg13g2_fill_2 FILLER_63_109 ();
 sg13g2_fill_1 FILLER_63_128 ();
 sg13g2_decap_4 FILLER_63_135 ();
 sg13g2_decap_4 FILLER_63_165 ();
 sg13g2_fill_1 FILLER_63_187 ();
 sg13g2_fill_1 FILLER_63_193 ();
 sg13g2_decap_8 FILLER_63_204 ();
 sg13g2_fill_1 FILLER_63_211 ();
 sg13g2_fill_2 FILLER_63_230 ();
 sg13g2_fill_1 FILLER_63_232 ();
 sg13g2_fill_2 FILLER_63_259 ();
 sg13g2_fill_2 FILLER_63_270 ();
 sg13g2_fill_2 FILLER_63_307 ();
 sg13g2_decap_8 FILLER_63_332 ();
 sg13g2_decap_4 FILLER_63_339 ();
 sg13g2_fill_2 FILLER_63_343 ();
 sg13g2_fill_1 FILLER_63_376 ();
 sg13g2_decap_8 FILLER_63_401 ();
 sg13g2_decap_4 FILLER_63_408 ();
 sg13g2_fill_1 FILLER_63_412 ();
 sg13g2_decap_8 FILLER_63_418 ();
 sg13g2_decap_8 FILLER_63_425 ();
 sg13g2_decap_8 FILLER_63_439 ();
 sg13g2_decap_4 FILLER_63_446 ();
 sg13g2_fill_2 FILLER_63_450 ();
 sg13g2_decap_8 FILLER_63_461 ();
 sg13g2_fill_2 FILLER_63_468 ();
 sg13g2_decap_8 FILLER_63_477 ();
 sg13g2_fill_2 FILLER_63_492 ();
 sg13g2_fill_2 FILLER_63_514 ();
 sg13g2_fill_2 FILLER_63_521 ();
 sg13g2_fill_2 FILLER_63_538 ();
 sg13g2_fill_1 FILLER_63_540 ();
 sg13g2_fill_2 FILLER_63_545 ();
 sg13g2_fill_2 FILLER_63_581 ();
 sg13g2_fill_1 FILLER_63_583 ();
 sg13g2_decap_4 FILLER_63_610 ();
 sg13g2_fill_1 FILLER_63_645 ();
 sg13g2_fill_1 FILLER_63_675 ();
 sg13g2_fill_2 FILLER_63_760 ();
 sg13g2_fill_2 FILLER_63_768 ();
 sg13g2_fill_2 FILLER_63_796 ();
 sg13g2_fill_1 FILLER_63_803 ();
 sg13g2_decap_8 FILLER_63_824 ();
 sg13g2_fill_1 FILLER_63_831 ();
 sg13g2_fill_1 FILLER_63_851 ();
 sg13g2_fill_1 FILLER_63_883 ();
 sg13g2_fill_2 FILLER_63_888 ();
 sg13g2_fill_1 FILLER_63_890 ();
 sg13g2_fill_2 FILLER_63_909 ();
 sg13g2_fill_1 FILLER_63_942 ();
 sg13g2_fill_1 FILLER_63_958 ();
 sg13g2_decap_8 FILLER_63_964 ();
 sg13g2_decap_4 FILLER_63_971 ();
 sg13g2_fill_1 FILLER_63_975 ();
 sg13g2_fill_1 FILLER_63_985 ();
 sg13g2_decap_4 FILLER_63_995 ();
 sg13g2_fill_1 FILLER_63_999 ();
 sg13g2_fill_2 FILLER_63_1035 ();
 sg13g2_decap_8 FILLER_63_1055 ();
 sg13g2_decap_4 FILLER_63_1076 ();
 sg13g2_fill_1 FILLER_63_1106 ();
 sg13g2_decap_8 FILLER_63_1112 ();
 sg13g2_decap_8 FILLER_63_1119 ();
 sg13g2_decap_4 FILLER_63_1126 ();
 sg13g2_fill_1 FILLER_63_1130 ();
 sg13g2_decap_4 FILLER_63_1141 ();
 sg13g2_fill_1 FILLER_63_1145 ();
 sg13g2_fill_2 FILLER_63_1150 ();
 sg13g2_fill_1 FILLER_63_1152 ();
 sg13g2_fill_1 FILLER_63_1158 ();
 sg13g2_decap_4 FILLER_63_1163 ();
 sg13g2_decap_8 FILLER_63_1185 ();
 sg13g2_decap_8 FILLER_63_1192 ();
 sg13g2_fill_2 FILLER_63_1199 ();
 sg13g2_fill_2 FILLER_63_1205 ();
 sg13g2_fill_1 FILLER_63_1207 ();
 sg13g2_decap_8 FILLER_63_1236 ();
 sg13g2_decap_4 FILLER_63_1247 ();
 sg13g2_fill_1 FILLER_63_1262 ();
 sg13g2_decap_4 FILLER_63_1284 ();
 sg13g2_fill_1 FILLER_63_1288 ();
 sg13g2_decap_8 FILLER_63_1294 ();
 sg13g2_decap_8 FILLER_63_1301 ();
 sg13g2_decap_8 FILLER_63_1308 ();
 sg13g2_decap_4 FILLER_63_1315 ();
 sg13g2_fill_2 FILLER_63_1319 ();
 sg13g2_fill_2 FILLER_63_1325 ();
 sg13g2_fill_1 FILLER_63_1327 ();
 sg13g2_fill_1 FILLER_63_1336 ();
 sg13g2_decap_8 FILLER_63_1371 ();
 sg13g2_decap_8 FILLER_63_1378 ();
 sg13g2_decap_4 FILLER_63_1421 ();
 sg13g2_fill_2 FILLER_63_1425 ();
 sg13g2_fill_2 FILLER_63_1430 ();
 sg13g2_fill_1 FILLER_63_1432 ();
 sg13g2_decap_4 FILLER_63_1438 ();
 sg13g2_fill_2 FILLER_63_1442 ();
 sg13g2_fill_2 FILLER_63_1453 ();
 sg13g2_decap_8 FILLER_63_1467 ();
 sg13g2_decap_4 FILLER_63_1474 ();
 sg13g2_fill_2 FILLER_63_1478 ();
 sg13g2_decap_4 FILLER_63_1484 ();
 sg13g2_decap_8 FILLER_63_1493 ();
 sg13g2_fill_2 FILLER_63_1500 ();
 sg13g2_fill_1 FILLER_63_1502 ();
 sg13g2_fill_2 FILLER_63_1538 ();
 sg13g2_fill_1 FILLER_63_1540 ();
 sg13g2_decap_4 FILLER_63_1572 ();
 sg13g2_decap_4 FILLER_63_1580 ();
 sg13g2_fill_2 FILLER_63_1584 ();
 sg13g2_decap_4 FILLER_63_1595 ();
 sg13g2_fill_1 FILLER_63_1599 ();
 sg13g2_decap_8 FILLER_63_1608 ();
 sg13g2_fill_1 FILLER_63_1615 ();
 sg13g2_fill_1 FILLER_63_1620 ();
 sg13g2_fill_2 FILLER_63_1625 ();
 sg13g2_fill_1 FILLER_63_1627 ();
 sg13g2_fill_2 FILLER_63_1640 ();
 sg13g2_fill_1 FILLER_63_1642 ();
 sg13g2_decap_4 FILLER_63_1678 ();
 sg13g2_fill_1 FILLER_63_1682 ();
 sg13g2_fill_2 FILLER_63_1691 ();
 sg13g2_decap_8 FILLER_63_1697 ();
 sg13g2_decap_8 FILLER_63_1704 ();
 sg13g2_decap_4 FILLER_63_1711 ();
 sg13g2_fill_1 FILLER_63_1715 ();
 sg13g2_fill_2 FILLER_63_1729 ();
 sg13g2_fill_1 FILLER_63_1731 ();
 sg13g2_fill_2 FILLER_63_1758 ();
 sg13g2_fill_2 FILLER_63_1765 ();
 sg13g2_fill_1 FILLER_63_1767 ();
 sg13g2_decap_8 FILLER_63_1772 ();
 sg13g2_decap_8 FILLER_63_1779 ();
 sg13g2_decap_4 FILLER_63_1786 ();
 sg13g2_decap_4 FILLER_63_1816 ();
 sg13g2_fill_1 FILLER_63_1820 ();
 sg13g2_decap_8 FILLER_63_1847 ();
 sg13g2_fill_1 FILLER_63_1854 ();
 sg13g2_fill_1 FILLER_63_1859 ();
 sg13g2_decap_4 FILLER_63_1869 ();
 sg13g2_fill_1 FILLER_63_1873 ();
 sg13g2_decap_4 FILLER_63_1900 ();
 sg13g2_fill_2 FILLER_63_1909 ();
 sg13g2_fill_1 FILLER_63_1911 ();
 sg13g2_decap_8 FILLER_63_1938 ();
 sg13g2_fill_2 FILLER_63_1945 ();
 sg13g2_decap_8 FILLER_63_1953 ();
 sg13g2_decap_4 FILLER_63_1960 ();
 sg13g2_fill_2 FILLER_63_1964 ();
 sg13g2_fill_2 FILLER_63_1974 ();
 sg13g2_fill_1 FILLER_63_1976 ();
 sg13g2_decap_8 FILLER_63_1998 ();
 sg13g2_fill_2 FILLER_63_2005 ();
 sg13g2_decap_8 FILLER_63_2018 ();
 sg13g2_fill_1 FILLER_63_2025 ();
 sg13g2_fill_2 FILLER_63_2039 ();
 sg13g2_fill_1 FILLER_63_2041 ();
 sg13g2_fill_2 FILLER_63_2053 ();
 sg13g2_fill_1 FILLER_63_2055 ();
 sg13g2_decap_8 FILLER_63_2069 ();
 sg13g2_decap_4 FILLER_63_2076 ();
 sg13g2_fill_1 FILLER_63_2080 ();
 sg13g2_decap_8 FILLER_63_2101 ();
 sg13g2_decap_4 FILLER_63_2108 ();
 sg13g2_fill_1 FILLER_63_2112 ();
 sg13g2_decap_4 FILLER_63_2136 ();
 sg13g2_fill_1 FILLER_63_2140 ();
 sg13g2_fill_1 FILLER_63_2145 ();
 sg13g2_decap_4 FILLER_63_2156 ();
 sg13g2_fill_1 FILLER_63_2160 ();
 sg13g2_decap_4 FILLER_63_2174 ();
 sg13g2_decap_4 FILLER_63_2188 ();
 sg13g2_fill_2 FILLER_63_2192 ();
 sg13g2_decap_8 FILLER_63_2207 ();
 sg13g2_fill_2 FILLER_63_2214 ();
 sg13g2_fill_1 FILLER_63_2216 ();
 sg13g2_decap_4 FILLER_63_2245 ();
 sg13g2_fill_2 FILLER_63_2249 ();
 sg13g2_fill_1 FILLER_63_2271 ();
 sg13g2_fill_2 FILLER_63_2286 ();
 sg13g2_fill_1 FILLER_63_2288 ();
 sg13g2_decap_8 FILLER_63_2298 ();
 sg13g2_decap_4 FILLER_63_2305 ();
 sg13g2_fill_2 FILLER_63_2309 ();
 sg13g2_decap_8 FILLER_63_2321 ();
 sg13g2_fill_2 FILLER_63_2328 ();
 sg13g2_fill_1 FILLER_63_2330 ();
 sg13g2_decap_4 FILLER_63_2337 ();
 sg13g2_fill_1 FILLER_63_2341 ();
 sg13g2_decap_4 FILLER_63_2345 ();
 sg13g2_fill_1 FILLER_63_2349 ();
 sg13g2_fill_2 FILLER_63_2379 ();
 sg13g2_fill_2 FILLER_63_2385 ();
 sg13g2_fill_1 FILLER_63_2387 ();
 sg13g2_fill_2 FILLER_63_2403 ();
 sg13g2_fill_1 FILLER_63_2405 ();
 sg13g2_decap_4 FILLER_63_2419 ();
 sg13g2_fill_1 FILLER_63_2423 ();
 sg13g2_decap_8 FILLER_63_2428 ();
 sg13g2_decap_8 FILLER_63_2435 ();
 sg13g2_decap_8 FILLER_63_2442 ();
 sg13g2_fill_2 FILLER_63_2449 ();
 sg13g2_fill_2 FILLER_63_2499 ();
 sg13g2_fill_1 FILLER_63_2501 ();
 sg13g2_decap_8 FILLER_63_2509 ();
 sg13g2_fill_1 FILLER_63_2544 ();
 sg13g2_fill_2 FILLER_63_2558 ();
 sg13g2_decap_8 FILLER_63_2569 ();
 sg13g2_decap_4 FILLER_63_2576 ();
 sg13g2_decap_4 FILLER_63_2595 ();
 sg13g2_decap_8 FILLER_63_2604 ();
 sg13g2_fill_2 FILLER_63_2611 ();
 sg13g2_fill_1 FILLER_63_2613 ();
 sg13g2_fill_1 FILLER_63_2619 ();
 sg13g2_decap_8 FILLER_63_2625 ();
 sg13g2_decap_8 FILLER_63_2632 ();
 sg13g2_decap_8 FILLER_63_2639 ();
 sg13g2_decap_8 FILLER_63_2646 ();
 sg13g2_fill_2 FILLER_63_2653 ();
 sg13g2_fill_1 FILLER_63_2684 ();
 sg13g2_fill_2 FILLER_63_2690 ();
 sg13g2_decap_8 FILLER_63_2697 ();
 sg13g2_decap_8 FILLER_63_2704 ();
 sg13g2_fill_2 FILLER_63_2715 ();
 sg13g2_fill_1 FILLER_63_2717 ();
 sg13g2_decap_4 FILLER_63_2726 ();
 sg13g2_fill_1 FILLER_63_2730 ();
 sg13g2_fill_2 FILLER_63_2735 ();
 sg13g2_fill_1 FILLER_63_2737 ();
 sg13g2_decap_8 FILLER_63_2743 ();
 sg13g2_decap_8 FILLER_63_2750 ();
 sg13g2_decap_8 FILLER_63_2757 ();
 sg13g2_decap_4 FILLER_63_2764 ();
 sg13g2_fill_1 FILLER_63_2768 ();
 sg13g2_decap_4 FILLER_63_2781 ();
 sg13g2_fill_1 FILLER_63_2785 ();
 sg13g2_decap_8 FILLER_63_2794 ();
 sg13g2_decap_8 FILLER_63_2801 ();
 sg13g2_fill_1 FILLER_63_2808 ();
 sg13g2_fill_2 FILLER_63_2832 ();
 sg13g2_decap_8 FILLER_63_2846 ();
 sg13g2_decap_4 FILLER_63_2853 ();
 sg13g2_fill_1 FILLER_63_2857 ();
 sg13g2_decap_8 FILLER_63_2881 ();
 sg13g2_fill_2 FILLER_63_2888 ();
 sg13g2_fill_2 FILLER_63_2902 ();
 sg13g2_decap_4 FILLER_63_2909 ();
 sg13g2_fill_1 FILLER_63_2913 ();
 sg13g2_decap_4 FILLER_63_2946 ();
 sg13g2_fill_1 FILLER_63_2950 ();
 sg13g2_fill_1 FILLER_63_2956 ();
 sg13g2_fill_2 FILLER_63_2967 ();
 sg13g2_fill_1 FILLER_63_2969 ();
 sg13g2_decap_8 FILLER_63_3003 ();
 sg13g2_decap_8 FILLER_63_3010 ();
 sg13g2_decap_8 FILLER_63_3017 ();
 sg13g2_decap_8 FILLER_63_3024 ();
 sg13g2_decap_8 FILLER_63_3031 ();
 sg13g2_decap_8 FILLER_63_3038 ();
 sg13g2_decap_8 FILLER_63_3045 ();
 sg13g2_decap_8 FILLER_63_3052 ();
 sg13g2_decap_8 FILLER_63_3059 ();
 sg13g2_decap_8 FILLER_63_3066 ();
 sg13g2_decap_8 FILLER_63_3073 ();
 sg13g2_decap_8 FILLER_63_3080 ();
 sg13g2_decap_8 FILLER_63_3087 ();
 sg13g2_decap_8 FILLER_63_3094 ();
 sg13g2_decap_8 FILLER_63_3101 ();
 sg13g2_decap_8 FILLER_63_3108 ();
 sg13g2_decap_8 FILLER_63_3115 ();
 sg13g2_decap_8 FILLER_63_3122 ();
 sg13g2_decap_8 FILLER_63_3129 ();
 sg13g2_decap_8 FILLER_63_3136 ();
 sg13g2_decap_8 FILLER_63_3143 ();
 sg13g2_decap_8 FILLER_63_3150 ();
 sg13g2_decap_8 FILLER_63_3157 ();
 sg13g2_decap_8 FILLER_63_3164 ();
 sg13g2_decap_8 FILLER_63_3171 ();
 sg13g2_decap_8 FILLER_63_3178 ();
 sg13g2_decap_8 FILLER_63_3185 ();
 sg13g2_decap_8 FILLER_63_3192 ();
 sg13g2_decap_8 FILLER_63_3199 ();
 sg13g2_decap_8 FILLER_63_3206 ();
 sg13g2_decap_8 FILLER_63_3213 ();
 sg13g2_decap_8 FILLER_63_3220 ();
 sg13g2_decap_8 FILLER_63_3227 ();
 sg13g2_decap_8 FILLER_63_3234 ();
 sg13g2_decap_8 FILLER_63_3241 ();
 sg13g2_decap_8 FILLER_63_3248 ();
 sg13g2_decap_8 FILLER_63_3255 ();
 sg13g2_decap_8 FILLER_63_3262 ();
 sg13g2_decap_8 FILLER_63_3269 ();
 sg13g2_decap_8 FILLER_63_3276 ();
 sg13g2_decap_8 FILLER_63_3283 ();
 sg13g2_decap_8 FILLER_63_3290 ();
 sg13g2_decap_8 FILLER_63_3297 ();
 sg13g2_decap_8 FILLER_63_3304 ();
 sg13g2_decap_8 FILLER_63_3311 ();
 sg13g2_decap_8 FILLER_63_3318 ();
 sg13g2_decap_8 FILLER_63_3325 ();
 sg13g2_decap_8 FILLER_63_3332 ();
 sg13g2_decap_8 FILLER_63_3339 ();
 sg13g2_decap_8 FILLER_63_3346 ();
 sg13g2_decap_8 FILLER_63_3353 ();
 sg13g2_decap_8 FILLER_63_3360 ();
 sg13g2_decap_8 FILLER_63_3367 ();
 sg13g2_decap_8 FILLER_63_3374 ();
 sg13g2_decap_8 FILLER_63_3381 ();
 sg13g2_decap_8 FILLER_63_3388 ();
 sg13g2_decap_8 FILLER_63_3395 ();
 sg13g2_decap_8 FILLER_63_3402 ();
 sg13g2_decap_8 FILLER_63_3409 ();
 sg13g2_decap_8 FILLER_63_3416 ();
 sg13g2_decap_8 FILLER_63_3423 ();
 sg13g2_decap_8 FILLER_63_3430 ();
 sg13g2_decap_8 FILLER_63_3437 ();
 sg13g2_decap_8 FILLER_63_3444 ();
 sg13g2_decap_8 FILLER_63_3451 ();
 sg13g2_decap_8 FILLER_63_3458 ();
 sg13g2_decap_8 FILLER_63_3465 ();
 sg13g2_decap_8 FILLER_63_3472 ();
 sg13g2_decap_8 FILLER_63_3479 ();
 sg13g2_decap_8 FILLER_63_3486 ();
 sg13g2_decap_8 FILLER_63_3493 ();
 sg13g2_decap_8 FILLER_63_3500 ();
 sg13g2_decap_8 FILLER_63_3507 ();
 sg13g2_decap_8 FILLER_63_3514 ();
 sg13g2_decap_8 FILLER_63_3521 ();
 sg13g2_decap_8 FILLER_63_3528 ();
 sg13g2_decap_8 FILLER_63_3535 ();
 sg13g2_decap_8 FILLER_63_3542 ();
 sg13g2_decap_8 FILLER_63_3549 ();
 sg13g2_decap_8 FILLER_63_3556 ();
 sg13g2_decap_8 FILLER_63_3563 ();
 sg13g2_decap_8 FILLER_63_3570 ();
 sg13g2_fill_2 FILLER_63_3577 ();
 sg13g2_fill_1 FILLER_63_3579 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_4 FILLER_64_7 ();
 sg13g2_decap_4 FILLER_64_15 ();
 sg13g2_fill_1 FILLER_64_19 ();
 sg13g2_fill_2 FILLER_64_51 ();
 sg13g2_fill_1 FILLER_64_53 ();
 sg13g2_decap_4 FILLER_64_60 ();
 sg13g2_fill_2 FILLER_64_64 ();
 sg13g2_fill_2 FILLER_64_76 ();
 sg13g2_fill_1 FILLER_64_78 ();
 sg13g2_fill_2 FILLER_64_84 ();
 sg13g2_fill_1 FILLER_64_86 ();
 sg13g2_decap_8 FILLER_64_103 ();
 sg13g2_fill_2 FILLER_64_110 ();
 sg13g2_fill_1 FILLER_64_112 ();
 sg13g2_decap_8 FILLER_64_136 ();
 sg13g2_fill_2 FILLER_64_143 ();
 sg13g2_fill_1 FILLER_64_145 ();
 sg13g2_fill_2 FILLER_64_165 ();
 sg13g2_fill_1 FILLER_64_167 ();
 sg13g2_decap_8 FILLER_64_234 ();
 sg13g2_fill_2 FILLER_64_241 ();
 sg13g2_decap_4 FILLER_64_269 ();
 sg13g2_fill_1 FILLER_64_273 ();
 sg13g2_decap_4 FILLER_64_296 ();
 sg13g2_fill_2 FILLER_64_300 ();
 sg13g2_fill_2 FILLER_64_328 ();
 sg13g2_fill_1 FILLER_64_330 ();
 sg13g2_fill_1 FILLER_64_384 ();
 sg13g2_fill_2 FILLER_64_391 ();
 sg13g2_fill_1 FILLER_64_445 ();
 sg13g2_fill_2 FILLER_64_454 ();
 sg13g2_fill_2 FILLER_64_467 ();
 sg13g2_fill_1 FILLER_64_469 ();
 sg13g2_fill_2 FILLER_64_485 ();
 sg13g2_fill_1 FILLER_64_487 ();
 sg13g2_decap_4 FILLER_64_513 ();
 sg13g2_decap_8 FILLER_64_540 ();
 sg13g2_decap_8 FILLER_64_547 ();
 sg13g2_decap_4 FILLER_64_554 ();
 sg13g2_fill_2 FILLER_64_558 ();
 sg13g2_fill_1 FILLER_64_565 ();
 sg13g2_decap_8 FILLER_64_575 ();
 sg13g2_fill_2 FILLER_64_591 ();
 sg13g2_fill_1 FILLER_64_738 ();
 sg13g2_fill_2 FILLER_64_763 ();
 sg13g2_fill_2 FILLER_64_770 ();
 sg13g2_fill_2 FILLER_64_791 ();
 sg13g2_fill_2 FILLER_64_810 ();
 sg13g2_decap_4 FILLER_64_827 ();
 sg13g2_fill_2 FILLER_64_831 ();
 sg13g2_decap_4 FILLER_64_839 ();
 sg13g2_fill_1 FILLER_64_854 ();
 sg13g2_decap_4 FILLER_64_873 ();
 sg13g2_fill_2 FILLER_64_877 ();
 sg13g2_fill_2 FILLER_64_893 ();
 sg13g2_fill_1 FILLER_64_895 ();
 sg13g2_fill_1 FILLER_64_927 ();
 sg13g2_fill_2 FILLER_64_968 ();
 sg13g2_fill_2 FILLER_64_996 ();
 sg13g2_decap_4 FILLER_64_1004 ();
 sg13g2_fill_1 FILLER_64_1013 ();
 sg13g2_decap_8 FILLER_64_1019 ();
 sg13g2_fill_2 FILLER_64_1026 ();
 sg13g2_fill_1 FILLER_64_1028 ();
 sg13g2_decap_8 FILLER_64_1055 ();
 sg13g2_decap_8 FILLER_64_1062 ();
 sg13g2_fill_1 FILLER_64_1069 ();
 sg13g2_fill_1 FILLER_64_1096 ();
 sg13g2_decap_8 FILLER_64_1120 ();
 sg13g2_decap_4 FILLER_64_1127 ();
 sg13g2_decap_8 FILLER_64_1145 ();
 sg13g2_decap_4 FILLER_64_1152 ();
 sg13g2_fill_1 FILLER_64_1156 ();
 sg13g2_decap_4 FILLER_64_1193 ();
 sg13g2_fill_2 FILLER_64_1197 ();
 sg13g2_fill_2 FILLER_64_1225 ();
 sg13g2_fill_2 FILLER_64_1258 ();
 sg13g2_decap_4 FILLER_64_1264 ();
 sg13g2_fill_1 FILLER_64_1268 ();
 sg13g2_decap_4 FILLER_64_1275 ();
 sg13g2_fill_2 FILLER_64_1292 ();
 sg13g2_fill_1 FILLER_64_1294 ();
 sg13g2_decap_8 FILLER_64_1325 ();
 sg13g2_fill_2 FILLER_64_1332 ();
 sg13g2_decap_4 FILLER_64_1350 ();
 sg13g2_fill_1 FILLER_64_1354 ();
 sg13g2_decap_4 FILLER_64_1359 ();
 sg13g2_fill_2 FILLER_64_1363 ();
 sg13g2_fill_2 FILLER_64_1391 ();
 sg13g2_fill_1 FILLER_64_1393 ();
 sg13g2_fill_1 FILLER_64_1408 ();
 sg13g2_fill_2 FILLER_64_1433 ();
 sg13g2_fill_1 FILLER_64_1448 ();
 sg13g2_fill_2 FILLER_64_1506 ();
 sg13g2_fill_1 FILLER_64_1508 ();
 sg13g2_fill_2 FILLER_64_1518 ();
 sg13g2_fill_1 FILLER_64_1520 ();
 sg13g2_fill_2 FILLER_64_1537 ();
 sg13g2_fill_2 FILLER_64_1562 ();
 sg13g2_fill_1 FILLER_64_1564 ();
 sg13g2_fill_2 FILLER_64_1580 ();
 sg13g2_fill_2 FILLER_64_1629 ();
 sg13g2_fill_1 FILLER_64_1631 ();
 sg13g2_decap_8 FILLER_64_1658 ();
 sg13g2_decap_4 FILLER_64_1665 ();
 sg13g2_decap_8 FILLER_64_1681 ();
 sg13g2_decap_4 FILLER_64_1688 ();
 sg13g2_decap_8 FILLER_64_1732 ();
 sg13g2_fill_1 FILLER_64_1739 ();
 sg13g2_decap_8 FILLER_64_1792 ();
 sg13g2_fill_2 FILLER_64_1799 ();
 sg13g2_fill_2 FILLER_64_1810 ();
 sg13g2_fill_1 FILLER_64_1812 ();
 sg13g2_fill_2 FILLER_64_1840 ();
 sg13g2_fill_2 FILLER_64_1847 ();
 sg13g2_fill_1 FILLER_64_1849 ();
 sg13g2_decap_8 FILLER_64_1889 ();
 sg13g2_fill_1 FILLER_64_1896 ();
 sg13g2_fill_2 FILLER_64_1912 ();
 sg13g2_fill_1 FILLER_64_1914 ();
 sg13g2_fill_2 FILLER_64_1929 ();
 sg13g2_decap_8 FILLER_64_1936 ();
 sg13g2_fill_1 FILLER_64_1943 ();
 sg13g2_fill_1 FILLER_64_1952 ();
 sg13g2_decap_4 FILLER_64_1961 ();
 sg13g2_fill_1 FILLER_64_1965 ();
 sg13g2_fill_2 FILLER_64_1977 ();
 sg13g2_fill_2 FILLER_64_2009 ();
 sg13g2_fill_1 FILLER_64_2011 ();
 sg13g2_decap_4 FILLER_64_2023 ();
 sg13g2_fill_2 FILLER_64_2049 ();
 sg13g2_fill_1 FILLER_64_2103 ();
 sg13g2_decap_4 FILLER_64_2113 ();
 sg13g2_decap_8 FILLER_64_2122 ();
 sg13g2_fill_2 FILLER_64_2133 ();
 sg13g2_fill_1 FILLER_64_2152 ();
 sg13g2_fill_2 FILLER_64_2161 ();
 sg13g2_fill_1 FILLER_64_2176 ();
 sg13g2_decap_8 FILLER_64_2197 ();
 sg13g2_decap_4 FILLER_64_2212 ();
 sg13g2_decap_4 FILLER_64_2220 ();
 sg13g2_fill_1 FILLER_64_2224 ();
 sg13g2_decap_4 FILLER_64_2230 ();
 sg13g2_fill_1 FILLER_64_2234 ();
 sg13g2_fill_2 FILLER_64_2244 ();
 sg13g2_fill_1 FILLER_64_2246 ();
 sg13g2_decap_8 FILLER_64_2255 ();
 sg13g2_decap_8 FILLER_64_2262 ();
 sg13g2_fill_1 FILLER_64_2269 ();
 sg13g2_decap_8 FILLER_64_2301 ();
 sg13g2_decap_4 FILLER_64_2347 ();
 sg13g2_decap_8 FILLER_64_2422 ();
 sg13g2_decap_8 FILLER_64_2429 ();
 sg13g2_decap_4 FILLER_64_2436 ();
 sg13g2_fill_2 FILLER_64_2440 ();
 sg13g2_decap_8 FILLER_64_2469 ();
 sg13g2_decap_8 FILLER_64_2476 ();
 sg13g2_decap_4 FILLER_64_2483 ();
 sg13g2_fill_2 FILLER_64_2498 ();
 sg13g2_fill_1 FILLER_64_2500 ();
 sg13g2_fill_2 FILLER_64_2553 ();
 sg13g2_fill_1 FILLER_64_2555 ();
 sg13g2_fill_2 FILLER_64_2576 ();
 sg13g2_decap_8 FILLER_64_2602 ();
 sg13g2_fill_2 FILLER_64_2609 ();
 sg13g2_decap_8 FILLER_64_2639 ();
 sg13g2_fill_2 FILLER_64_2646 ();
 sg13g2_fill_1 FILLER_64_2648 ();
 sg13g2_fill_1 FILLER_64_2667 ();
 sg13g2_decap_4 FILLER_64_2677 ();
 sg13g2_fill_1 FILLER_64_2681 ();
 sg13g2_fill_1 FILLER_64_2706 ();
 sg13g2_fill_2 FILLER_64_2721 ();
 sg13g2_decap_4 FILLER_64_2727 ();
 sg13g2_fill_1 FILLER_64_2767 ();
 sg13g2_fill_1 FILLER_64_2784 ();
 sg13g2_decap_4 FILLER_64_2798 ();
 sg13g2_fill_2 FILLER_64_2802 ();
 sg13g2_decap_4 FILLER_64_2808 ();
 sg13g2_decap_8 FILLER_64_2827 ();
 sg13g2_fill_2 FILLER_64_2834 ();
 sg13g2_decap_4 FILLER_64_2841 ();
 sg13g2_fill_2 FILLER_64_2845 ();
 sg13g2_decap_4 FILLER_64_2862 ();
 sg13g2_fill_2 FILLER_64_2866 ();
 sg13g2_decap_8 FILLER_64_2872 ();
 sg13g2_decap_8 FILLER_64_2879 ();
 sg13g2_fill_2 FILLER_64_2886 ();
 sg13g2_fill_1 FILLER_64_2888 ();
 sg13g2_decap_4 FILLER_64_2925 ();
 sg13g2_decap_4 FILLER_64_2933 ();
 sg13g2_fill_2 FILLER_64_2937 ();
 sg13g2_decap_4 FILLER_64_2947 ();
 sg13g2_fill_1 FILLER_64_2951 ();
 sg13g2_fill_2 FILLER_64_2965 ();
 sg13g2_fill_1 FILLER_64_2967 ();
 sg13g2_decap_8 FILLER_64_2975 ();
 sg13g2_fill_1 FILLER_64_2986 ();
 sg13g2_decap_8 FILLER_64_3000 ();
 sg13g2_decap_8 FILLER_64_3007 ();
 sg13g2_decap_8 FILLER_64_3014 ();
 sg13g2_decap_8 FILLER_64_3021 ();
 sg13g2_decap_8 FILLER_64_3028 ();
 sg13g2_decap_8 FILLER_64_3035 ();
 sg13g2_decap_8 FILLER_64_3042 ();
 sg13g2_decap_8 FILLER_64_3049 ();
 sg13g2_decap_8 FILLER_64_3056 ();
 sg13g2_decap_8 FILLER_64_3063 ();
 sg13g2_decap_8 FILLER_64_3070 ();
 sg13g2_decap_8 FILLER_64_3077 ();
 sg13g2_decap_8 FILLER_64_3084 ();
 sg13g2_decap_8 FILLER_64_3091 ();
 sg13g2_decap_8 FILLER_64_3098 ();
 sg13g2_decap_8 FILLER_64_3105 ();
 sg13g2_decap_8 FILLER_64_3112 ();
 sg13g2_decap_8 FILLER_64_3119 ();
 sg13g2_decap_8 FILLER_64_3126 ();
 sg13g2_decap_8 FILLER_64_3133 ();
 sg13g2_decap_8 FILLER_64_3140 ();
 sg13g2_decap_8 FILLER_64_3147 ();
 sg13g2_decap_8 FILLER_64_3154 ();
 sg13g2_decap_8 FILLER_64_3161 ();
 sg13g2_decap_8 FILLER_64_3168 ();
 sg13g2_decap_8 FILLER_64_3175 ();
 sg13g2_decap_8 FILLER_64_3182 ();
 sg13g2_decap_8 FILLER_64_3189 ();
 sg13g2_decap_8 FILLER_64_3196 ();
 sg13g2_decap_8 FILLER_64_3203 ();
 sg13g2_decap_8 FILLER_64_3210 ();
 sg13g2_decap_8 FILLER_64_3217 ();
 sg13g2_decap_8 FILLER_64_3224 ();
 sg13g2_decap_8 FILLER_64_3231 ();
 sg13g2_decap_8 FILLER_64_3238 ();
 sg13g2_decap_8 FILLER_64_3245 ();
 sg13g2_decap_8 FILLER_64_3252 ();
 sg13g2_decap_8 FILLER_64_3259 ();
 sg13g2_decap_8 FILLER_64_3266 ();
 sg13g2_decap_8 FILLER_64_3273 ();
 sg13g2_decap_8 FILLER_64_3280 ();
 sg13g2_decap_8 FILLER_64_3287 ();
 sg13g2_decap_8 FILLER_64_3294 ();
 sg13g2_decap_8 FILLER_64_3301 ();
 sg13g2_decap_8 FILLER_64_3308 ();
 sg13g2_decap_8 FILLER_64_3315 ();
 sg13g2_decap_8 FILLER_64_3322 ();
 sg13g2_decap_8 FILLER_64_3329 ();
 sg13g2_decap_8 FILLER_64_3336 ();
 sg13g2_decap_8 FILLER_64_3343 ();
 sg13g2_decap_8 FILLER_64_3350 ();
 sg13g2_decap_8 FILLER_64_3357 ();
 sg13g2_decap_8 FILLER_64_3364 ();
 sg13g2_decap_8 FILLER_64_3371 ();
 sg13g2_decap_8 FILLER_64_3378 ();
 sg13g2_decap_8 FILLER_64_3385 ();
 sg13g2_decap_8 FILLER_64_3392 ();
 sg13g2_decap_8 FILLER_64_3399 ();
 sg13g2_decap_8 FILLER_64_3406 ();
 sg13g2_decap_8 FILLER_64_3413 ();
 sg13g2_decap_8 FILLER_64_3420 ();
 sg13g2_decap_8 FILLER_64_3427 ();
 sg13g2_decap_8 FILLER_64_3434 ();
 sg13g2_decap_8 FILLER_64_3441 ();
 sg13g2_decap_8 FILLER_64_3448 ();
 sg13g2_decap_8 FILLER_64_3455 ();
 sg13g2_decap_8 FILLER_64_3462 ();
 sg13g2_decap_8 FILLER_64_3469 ();
 sg13g2_decap_8 FILLER_64_3476 ();
 sg13g2_decap_8 FILLER_64_3483 ();
 sg13g2_decap_8 FILLER_64_3490 ();
 sg13g2_decap_8 FILLER_64_3497 ();
 sg13g2_decap_8 FILLER_64_3504 ();
 sg13g2_decap_8 FILLER_64_3511 ();
 sg13g2_decap_8 FILLER_64_3518 ();
 sg13g2_decap_8 FILLER_64_3525 ();
 sg13g2_decap_8 FILLER_64_3532 ();
 sg13g2_decap_8 FILLER_64_3539 ();
 sg13g2_decap_8 FILLER_64_3546 ();
 sg13g2_decap_8 FILLER_64_3553 ();
 sg13g2_decap_8 FILLER_64_3560 ();
 sg13g2_decap_8 FILLER_64_3567 ();
 sg13g2_decap_4 FILLER_64_3574 ();
 sg13g2_fill_2 FILLER_64_3578 ();
 sg13g2_fill_2 FILLER_65_26 ();
 sg13g2_fill_1 FILLER_65_28 ();
 sg13g2_decap_4 FILLER_65_51 ();
 sg13g2_decap_4 FILLER_65_73 ();
 sg13g2_fill_1 FILLER_65_77 ();
 sg13g2_decap_4 FILLER_65_86 ();
 sg13g2_decap_8 FILLER_65_100 ();
 sg13g2_decap_4 FILLER_65_111 ();
 sg13g2_fill_1 FILLER_65_152 ();
 sg13g2_fill_2 FILLER_65_175 ();
 sg13g2_fill_1 FILLER_65_177 ();
 sg13g2_decap_8 FILLER_65_206 ();
 sg13g2_decap_4 FILLER_65_213 ();
 sg13g2_fill_1 FILLER_65_217 ();
 sg13g2_decap_8 FILLER_65_235 ();
 sg13g2_decap_8 FILLER_65_242 ();
 sg13g2_fill_1 FILLER_65_249 ();
 sg13g2_fill_2 FILLER_65_257 ();
 sg13g2_fill_1 FILLER_65_259 ();
 sg13g2_decap_8 FILLER_65_272 ();
 sg13g2_decap_4 FILLER_65_279 ();
 sg13g2_fill_2 FILLER_65_283 ();
 sg13g2_decap_4 FILLER_65_298 ();
 sg13g2_fill_2 FILLER_65_302 ();
 sg13g2_decap_8 FILLER_65_327 ();
 sg13g2_fill_1 FILLER_65_360 ();
 sg13g2_decap_8 FILLER_65_429 ();
 sg13g2_decap_8 FILLER_65_436 ();
 sg13g2_decap_4 FILLER_65_443 ();
 sg13g2_fill_1 FILLER_65_447 ();
 sg13g2_decap_4 FILLER_65_456 ();
 sg13g2_decap_8 FILLER_65_465 ();
 sg13g2_fill_2 FILLER_65_472 ();
 sg13g2_decap_4 FILLER_65_480 ();
 sg13g2_fill_1 FILLER_65_484 ();
 sg13g2_fill_2 FILLER_65_494 ();
 sg13g2_fill_2 FILLER_65_502 ();
 sg13g2_decap_4 FILLER_65_520 ();
 sg13g2_fill_1 FILLER_65_524 ();
 sg13g2_decap_8 FILLER_65_533 ();
 sg13g2_decap_8 FILLER_65_540 ();
 sg13g2_fill_1 FILLER_65_560 ();
 sg13g2_fill_1 FILLER_65_599 ();
 sg13g2_fill_1 FILLER_65_608 ();
 sg13g2_fill_2 FILLER_65_666 ();
 sg13g2_fill_2 FILLER_65_685 ();
 sg13g2_decap_4 FILLER_65_691 ();
 sg13g2_fill_1 FILLER_65_695 ();
 sg13g2_decap_4 FILLER_65_700 ();
 sg13g2_fill_1 FILLER_65_713 ();
 sg13g2_fill_2 FILLER_65_731 ();
 sg13g2_fill_1 FILLER_65_742 ();
 sg13g2_decap_4 FILLER_65_755 ();
 sg13g2_decap_4 FILLER_65_763 ();
 sg13g2_fill_1 FILLER_65_793 ();
 sg13g2_decap_8 FILLER_65_822 ();
 sg13g2_fill_2 FILLER_65_829 ();
 sg13g2_fill_2 FILLER_65_852 ();
 sg13g2_fill_1 FILLER_65_854 ();
 sg13g2_fill_1 FILLER_65_907 ();
 sg13g2_decap_4 FILLER_65_917 ();
 sg13g2_decap_8 FILLER_65_930 ();
 sg13g2_fill_1 FILLER_65_937 ();
 sg13g2_decap_4 FILLER_65_942 ();
 sg13g2_fill_1 FILLER_65_962 ();
 sg13g2_decap_8 FILLER_65_972 ();
 sg13g2_fill_2 FILLER_65_979 ();
 sg13g2_fill_2 FILLER_65_985 ();
 sg13g2_decap_4 FILLER_65_1019 ();
 sg13g2_fill_1 FILLER_65_1023 ();
 sg13g2_fill_2 FILLER_65_1093 ();
 sg13g2_fill_2 FILLER_65_1124 ();
 sg13g2_decap_8 FILLER_65_1152 ();
 sg13g2_decap_4 FILLER_65_1190 ();
 sg13g2_fill_2 FILLER_65_1194 ();
 sg13g2_fill_2 FILLER_65_1201 ();
 sg13g2_fill_1 FILLER_65_1203 ();
 sg13g2_fill_1 FILLER_65_1209 ();
 sg13g2_decap_4 FILLER_65_1214 ();
 sg13g2_fill_1 FILLER_65_1218 ();
 sg13g2_fill_2 FILLER_65_1233 ();
 sg13g2_decap_8 FILLER_65_1240 ();
 sg13g2_fill_1 FILLER_65_1247 ();
 sg13g2_fill_1 FILLER_65_1269 ();
 sg13g2_fill_2 FILLER_65_1292 ();
 sg13g2_decap_4 FILLER_65_1334 ();
 sg13g2_fill_1 FILLER_65_1338 ();
 sg13g2_decap_8 FILLER_65_1343 ();
 sg13g2_decap_4 FILLER_65_1368 ();
 sg13g2_fill_2 FILLER_65_1421 ();
 sg13g2_fill_1 FILLER_65_1423 ();
 sg13g2_fill_2 FILLER_65_1454 ();
 sg13g2_fill_1 FILLER_65_1456 ();
 sg13g2_fill_2 FILLER_65_1462 ();
 sg13g2_fill_1 FILLER_65_1469 ();
 sg13g2_decap_8 FILLER_65_1483 ();
 sg13g2_fill_1 FILLER_65_1490 ();
 sg13g2_decap_8 FILLER_65_1495 ();
 sg13g2_fill_2 FILLER_65_1502 ();
 sg13g2_fill_1 FILLER_65_1504 ();
 sg13g2_fill_1 FILLER_65_1536 ();
 sg13g2_fill_2 FILLER_65_1547 ();
 sg13g2_decap_8 FILLER_65_1575 ();
 sg13g2_decap_8 FILLER_65_1582 ();
 sg13g2_decap_4 FILLER_65_1589 ();
 sg13g2_decap_8 FILLER_65_1605 ();
 sg13g2_decap_4 FILLER_65_1612 ();
 sg13g2_fill_2 FILLER_65_1616 ();
 sg13g2_fill_2 FILLER_65_1631 ();
 sg13g2_fill_1 FILLER_65_1642 ();
 sg13g2_decap_8 FILLER_65_1655 ();
 sg13g2_decap_4 FILLER_65_1662 ();
 sg13g2_fill_2 FILLER_65_1705 ();
 sg13g2_fill_1 FILLER_65_1733 ();
 sg13g2_decap_4 FILLER_65_1749 ();
 sg13g2_fill_2 FILLER_65_1795 ();
 sg13g2_decap_8 FILLER_65_1815 ();
 sg13g2_fill_2 FILLER_65_1865 ();
 sg13g2_fill_1 FILLER_65_1867 ();
 sg13g2_fill_2 FILLER_65_1873 ();
 sg13g2_decap_8 FILLER_65_1879 ();
 sg13g2_decap_4 FILLER_65_1899 ();
 sg13g2_fill_1 FILLER_65_1911 ();
 sg13g2_decap_4 FILLER_65_1917 ();
 sg13g2_fill_2 FILLER_65_1921 ();
 sg13g2_fill_1 FILLER_65_1927 ();
 sg13g2_decap_4 FILLER_65_1933 ();
 sg13g2_fill_1 FILLER_65_1937 ();
 sg13g2_decap_8 FILLER_65_1957 ();
 sg13g2_decap_8 FILLER_65_1964 ();
 sg13g2_fill_2 FILLER_65_1971 ();
 sg13g2_fill_1 FILLER_65_1973 ();
 sg13g2_fill_2 FILLER_65_2001 ();
 sg13g2_fill_2 FILLER_65_2010 ();
 sg13g2_fill_1 FILLER_65_2012 ();
 sg13g2_decap_8 FILLER_65_2018 ();
 sg13g2_decap_8 FILLER_65_2025 ();
 sg13g2_decap_4 FILLER_65_2032 ();
 sg13g2_fill_1 FILLER_65_2036 ();
 sg13g2_fill_2 FILLER_65_2042 ();
 sg13g2_decap_8 FILLER_65_2069 ();
 sg13g2_fill_2 FILLER_65_2076 ();
 sg13g2_fill_1 FILLER_65_2078 ();
 sg13g2_decap_8 FILLER_65_2112 ();
 sg13g2_decap_4 FILLER_65_2119 ();
 sg13g2_decap_8 FILLER_65_2131 ();
 sg13g2_fill_2 FILLER_65_2142 ();
 sg13g2_fill_1 FILLER_65_2144 ();
 sg13g2_decap_8 FILLER_65_2157 ();
 sg13g2_decap_8 FILLER_65_2164 ();
 sg13g2_decap_8 FILLER_65_2171 ();
 sg13g2_decap_8 FILLER_65_2178 ();
 sg13g2_fill_1 FILLER_65_2185 ();
 sg13g2_fill_2 FILLER_65_2199 ();
 sg13g2_decap_4 FILLER_65_2206 ();
 sg13g2_fill_2 FILLER_65_2224 ();
 sg13g2_fill_1 FILLER_65_2226 ();
 sg13g2_fill_2 FILLER_65_2240 ();
 sg13g2_decap_4 FILLER_65_2260 ();
 sg13g2_fill_1 FILLER_65_2264 ();
 sg13g2_fill_1 FILLER_65_2270 ();
 sg13g2_fill_2 FILLER_65_2290 ();
 sg13g2_fill_2 FILLER_65_2297 ();
 sg13g2_fill_1 FILLER_65_2308 ();
 sg13g2_decap_8 FILLER_65_2315 ();
 sg13g2_decap_8 FILLER_65_2322 ();
 sg13g2_fill_2 FILLER_65_2368 ();
 sg13g2_decap_8 FILLER_65_2396 ();
 sg13g2_decap_4 FILLER_65_2403 ();
 sg13g2_fill_1 FILLER_65_2407 ();
 sg13g2_decap_4 FILLER_65_2439 ();
 sg13g2_fill_1 FILLER_65_2443 ();
 sg13g2_fill_1 FILLER_65_2468 ();
 sg13g2_decap_4 FILLER_65_2495 ();
 sg13g2_fill_1 FILLER_65_2499 ();
 sg13g2_fill_2 FILLER_65_2507 ();
 sg13g2_decap_8 FILLER_65_2522 ();
 sg13g2_decap_8 FILLER_65_2529 ();
 sg13g2_fill_2 FILLER_65_2540 ();
 sg13g2_decap_4 FILLER_65_2551 ();
 sg13g2_fill_2 FILLER_65_2559 ();
 sg13g2_fill_2 FILLER_65_2571 ();
 sg13g2_fill_1 FILLER_65_2578 ();
 sg13g2_fill_2 FILLER_65_2593 ();
 sg13g2_fill_1 FILLER_65_2595 ();
 sg13g2_decap_8 FILLER_65_2606 ();
 sg13g2_decap_8 FILLER_65_2613 ();
 sg13g2_decap_8 FILLER_65_2639 ();
 sg13g2_decap_4 FILLER_65_2646 ();
 sg13g2_fill_1 FILLER_65_2662 ();
 sg13g2_fill_2 FILLER_65_2682 ();
 sg13g2_fill_1 FILLER_65_2684 ();
 sg13g2_fill_1 FILLER_65_2693 ();
 sg13g2_fill_2 FILLER_65_2698 ();
 sg13g2_decap_4 FILLER_65_2714 ();
 sg13g2_fill_1 FILLER_65_2718 ();
 sg13g2_decap_8 FILLER_65_2723 ();
 sg13g2_decap_8 FILLER_65_2730 ();
 sg13g2_decap_8 FILLER_65_2737 ();
 sg13g2_fill_2 FILLER_65_2744 ();
 sg13g2_decap_4 FILLER_65_2758 ();
 sg13g2_fill_2 FILLER_65_2762 ();
 sg13g2_fill_2 FILLER_65_2774 ();
 sg13g2_fill_2 FILLER_65_2781 ();
 sg13g2_fill_2 FILLER_65_2794 ();
 sg13g2_fill_2 FILLER_65_2804 ();
 sg13g2_fill_2 FILLER_65_2822 ();
 sg13g2_fill_1 FILLER_65_2832 ();
 sg13g2_fill_2 FILLER_65_2846 ();
 sg13g2_fill_1 FILLER_65_2848 ();
 sg13g2_decap_8 FILLER_65_2883 ();
 sg13g2_decap_4 FILLER_65_2895 ();
 sg13g2_fill_2 FILLER_65_2902 ();
 sg13g2_fill_1 FILLER_65_2904 ();
 sg13g2_decap_8 FILLER_65_2914 ();
 sg13g2_fill_2 FILLER_65_2921 ();
 sg13g2_fill_1 FILLER_65_2923 ();
 sg13g2_decap_4 FILLER_65_2967 ();
 sg13g2_decap_8 FILLER_65_2997 ();
 sg13g2_decap_8 FILLER_65_3004 ();
 sg13g2_decap_8 FILLER_65_3011 ();
 sg13g2_decap_8 FILLER_65_3018 ();
 sg13g2_decap_8 FILLER_65_3025 ();
 sg13g2_decap_8 FILLER_65_3032 ();
 sg13g2_decap_8 FILLER_65_3039 ();
 sg13g2_decap_8 FILLER_65_3046 ();
 sg13g2_decap_8 FILLER_65_3053 ();
 sg13g2_decap_8 FILLER_65_3060 ();
 sg13g2_decap_8 FILLER_65_3067 ();
 sg13g2_decap_8 FILLER_65_3074 ();
 sg13g2_decap_8 FILLER_65_3081 ();
 sg13g2_decap_8 FILLER_65_3088 ();
 sg13g2_decap_8 FILLER_65_3095 ();
 sg13g2_decap_8 FILLER_65_3102 ();
 sg13g2_decap_8 FILLER_65_3109 ();
 sg13g2_decap_8 FILLER_65_3116 ();
 sg13g2_decap_8 FILLER_65_3123 ();
 sg13g2_decap_8 FILLER_65_3130 ();
 sg13g2_decap_8 FILLER_65_3137 ();
 sg13g2_decap_8 FILLER_65_3144 ();
 sg13g2_decap_8 FILLER_65_3151 ();
 sg13g2_decap_8 FILLER_65_3158 ();
 sg13g2_decap_8 FILLER_65_3165 ();
 sg13g2_decap_8 FILLER_65_3172 ();
 sg13g2_decap_8 FILLER_65_3179 ();
 sg13g2_decap_8 FILLER_65_3186 ();
 sg13g2_decap_8 FILLER_65_3193 ();
 sg13g2_decap_8 FILLER_65_3200 ();
 sg13g2_decap_8 FILLER_65_3207 ();
 sg13g2_decap_8 FILLER_65_3214 ();
 sg13g2_decap_8 FILLER_65_3221 ();
 sg13g2_decap_8 FILLER_65_3228 ();
 sg13g2_decap_8 FILLER_65_3235 ();
 sg13g2_decap_8 FILLER_65_3242 ();
 sg13g2_decap_8 FILLER_65_3249 ();
 sg13g2_decap_8 FILLER_65_3256 ();
 sg13g2_decap_8 FILLER_65_3263 ();
 sg13g2_decap_8 FILLER_65_3270 ();
 sg13g2_decap_8 FILLER_65_3277 ();
 sg13g2_decap_8 FILLER_65_3284 ();
 sg13g2_decap_8 FILLER_65_3291 ();
 sg13g2_decap_8 FILLER_65_3298 ();
 sg13g2_decap_8 FILLER_65_3305 ();
 sg13g2_decap_8 FILLER_65_3312 ();
 sg13g2_decap_8 FILLER_65_3319 ();
 sg13g2_decap_8 FILLER_65_3326 ();
 sg13g2_decap_8 FILLER_65_3333 ();
 sg13g2_decap_8 FILLER_65_3340 ();
 sg13g2_decap_8 FILLER_65_3347 ();
 sg13g2_decap_8 FILLER_65_3354 ();
 sg13g2_decap_8 FILLER_65_3361 ();
 sg13g2_decap_8 FILLER_65_3368 ();
 sg13g2_decap_8 FILLER_65_3375 ();
 sg13g2_decap_8 FILLER_65_3382 ();
 sg13g2_decap_8 FILLER_65_3389 ();
 sg13g2_decap_8 FILLER_65_3396 ();
 sg13g2_decap_8 FILLER_65_3403 ();
 sg13g2_decap_8 FILLER_65_3410 ();
 sg13g2_decap_8 FILLER_65_3417 ();
 sg13g2_decap_8 FILLER_65_3424 ();
 sg13g2_decap_8 FILLER_65_3431 ();
 sg13g2_decap_8 FILLER_65_3438 ();
 sg13g2_decap_8 FILLER_65_3445 ();
 sg13g2_decap_8 FILLER_65_3452 ();
 sg13g2_decap_8 FILLER_65_3459 ();
 sg13g2_decap_8 FILLER_65_3466 ();
 sg13g2_decap_8 FILLER_65_3473 ();
 sg13g2_decap_8 FILLER_65_3480 ();
 sg13g2_decap_8 FILLER_65_3487 ();
 sg13g2_decap_8 FILLER_65_3494 ();
 sg13g2_decap_8 FILLER_65_3501 ();
 sg13g2_decap_8 FILLER_65_3508 ();
 sg13g2_decap_8 FILLER_65_3515 ();
 sg13g2_decap_8 FILLER_65_3522 ();
 sg13g2_decap_8 FILLER_65_3529 ();
 sg13g2_decap_8 FILLER_65_3536 ();
 sg13g2_decap_8 FILLER_65_3543 ();
 sg13g2_decap_8 FILLER_65_3550 ();
 sg13g2_decap_8 FILLER_65_3557 ();
 sg13g2_decap_8 FILLER_65_3564 ();
 sg13g2_decap_8 FILLER_65_3571 ();
 sg13g2_fill_2 FILLER_65_3578 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_54 ();
 sg13g2_fill_2 FILLER_66_61 ();
 sg13g2_fill_1 FILLER_66_63 ();
 sg13g2_decap_4 FILLER_66_94 ();
 sg13g2_fill_1 FILLER_66_108 ();
 sg13g2_fill_2 FILLER_66_114 ();
 sg13g2_decap_8 FILLER_66_124 ();
 sg13g2_decap_4 FILLER_66_131 ();
 sg13g2_fill_2 FILLER_66_135 ();
 sg13g2_decap_8 FILLER_66_141 ();
 sg13g2_fill_1 FILLER_66_148 ();
 sg13g2_decap_4 FILLER_66_180 ();
 sg13g2_fill_2 FILLER_66_184 ();
 sg13g2_decap_8 FILLER_66_212 ();
 sg13g2_fill_2 FILLER_66_219 ();
 sg13g2_fill_1 FILLER_66_221 ();
 sg13g2_fill_2 FILLER_66_248 ();
 sg13g2_fill_2 FILLER_66_263 ();
 sg13g2_fill_1 FILLER_66_265 ();
 sg13g2_decap_4 FILLER_66_276 ();
 sg13g2_fill_2 FILLER_66_303 ();
 sg13g2_decap_8 FILLER_66_313 ();
 sg13g2_decap_4 FILLER_66_320 ();
 sg13g2_fill_2 FILLER_66_324 ();
 sg13g2_fill_1 FILLER_66_370 ();
 sg13g2_fill_2 FILLER_66_402 ();
 sg13g2_fill_1 FILLER_66_404 ();
 sg13g2_decap_4 FILLER_66_440 ();
 sg13g2_fill_1 FILLER_66_444 ();
 sg13g2_fill_2 FILLER_66_511 ();
 sg13g2_fill_1 FILLER_66_520 ();
 sg13g2_fill_2 FILLER_66_533 ();
 sg13g2_fill_1 FILLER_66_535 ();
 sg13g2_fill_1 FILLER_66_549 ();
 sg13g2_decap_8 FILLER_66_562 ();
 sg13g2_decap_8 FILLER_66_569 ();
 sg13g2_decap_4 FILLER_66_580 ();
 sg13g2_decap_8 FILLER_66_588 ();
 sg13g2_decap_8 FILLER_66_595 ();
 sg13g2_decap_4 FILLER_66_602 ();
 sg13g2_fill_2 FILLER_66_606 ();
 sg13g2_fill_1 FILLER_66_634 ();
 sg13g2_fill_2 FILLER_66_725 ();
 sg13g2_fill_1 FILLER_66_727 ();
 sg13g2_fill_2 FILLER_66_733 ();
 sg13g2_fill_1 FILLER_66_735 ();
 sg13g2_fill_1 FILLER_66_755 ();
 sg13g2_decap_8 FILLER_66_762 ();
 sg13g2_decap_4 FILLER_66_769 ();
 sg13g2_fill_2 FILLER_66_786 ();
 sg13g2_decap_8 FILLER_66_875 ();
 sg13g2_decap_8 FILLER_66_882 ();
 sg13g2_fill_2 FILLER_66_889 ();
 sg13g2_fill_1 FILLER_66_891 ();
 sg13g2_decap_4 FILLER_66_896 ();
 sg13g2_fill_1 FILLER_66_900 ();
 sg13g2_fill_2 FILLER_66_932 ();
 sg13g2_decap_4 FILLER_66_942 ();
 sg13g2_fill_1 FILLER_66_977 ();
 sg13g2_fill_2 FILLER_66_1030 ();
 sg13g2_fill_2 FILLER_66_1116 ();
 sg13g2_fill_1 FILLER_66_1135 ();
 sg13g2_decap_4 FILLER_66_1164 ();
 sg13g2_fill_2 FILLER_66_1168 ();
 sg13g2_fill_2 FILLER_66_1189 ();
 sg13g2_fill_1 FILLER_66_1191 ();
 sg13g2_decap_4 FILLER_66_1223 ();
 sg13g2_fill_1 FILLER_66_1236 ();
 sg13g2_fill_2 FILLER_66_1261 ();
 sg13g2_fill_1 FILLER_66_1263 ();
 sg13g2_fill_1 FILLER_66_1269 ();
 sg13g2_fill_2 FILLER_66_1302 ();
 sg13g2_fill_2 FILLER_66_1313 ();
 sg13g2_fill_1 FILLER_66_1315 ();
 sg13g2_decap_4 FILLER_66_1372 ();
 sg13g2_fill_1 FILLER_66_1393 ();
 sg13g2_fill_2 FILLER_66_1433 ();
 sg13g2_decap_8 FILLER_66_1439 ();
 sg13g2_decap_8 FILLER_66_1446 ();
 sg13g2_fill_2 FILLER_66_1466 ();
 sg13g2_decap_4 FILLER_66_1481 ();
 sg13g2_fill_2 FILLER_66_1485 ();
 sg13g2_decap_8 FILLER_66_1491 ();
 sg13g2_decap_4 FILLER_66_1511 ();
 sg13g2_fill_1 FILLER_66_1527 ();
 sg13g2_fill_1 FILLER_66_1556 ();
 sg13g2_fill_1 FILLER_66_1565 ();
 sg13g2_fill_2 FILLER_66_1602 ();
 sg13g2_fill_1 FILLER_66_1604 ();
 sg13g2_fill_1 FILLER_66_1640 ();
 sg13g2_fill_2 FILLER_66_1646 ();
 sg13g2_decap_4 FILLER_66_1674 ();
 sg13g2_fill_1 FILLER_66_1678 ();
 sg13g2_fill_1 FILLER_66_1687 ();
 sg13g2_fill_1 FILLER_66_1697 ();
 sg13g2_decap_8 FILLER_66_1703 ();
 sg13g2_fill_1 FILLER_66_1710 ();
 sg13g2_fill_2 FILLER_66_1715 ();
 sg13g2_decap_8 FILLER_66_1730 ();
 sg13g2_fill_1 FILLER_66_1737 ();
 sg13g2_fill_2 FILLER_66_1746 ();
 sg13g2_fill_1 FILLER_66_1756 ();
 sg13g2_decap_4 FILLER_66_1788 ();
 sg13g2_fill_1 FILLER_66_1792 ();
 sg13g2_decap_8 FILLER_66_1824 ();
 sg13g2_decap_4 FILLER_66_1831 ();
 sg13g2_fill_1 FILLER_66_1835 ();
 sg13g2_decap_8 FILLER_66_1849 ();
 sg13g2_decap_8 FILLER_66_1856 ();
 sg13g2_decap_4 FILLER_66_1873 ();
 sg13g2_fill_2 FILLER_66_1877 ();
 sg13g2_decap_8 FILLER_66_1885 ();
 sg13g2_decap_8 FILLER_66_1892 ();
 sg13g2_fill_1 FILLER_66_1899 ();
 sg13g2_fill_1 FILLER_66_1908 ();
 sg13g2_fill_2 FILLER_66_1919 ();
 sg13g2_fill_1 FILLER_66_1921 ();
 sg13g2_fill_2 FILLER_66_1953 ();
 sg13g2_decap_8 FILLER_66_1968 ();
 sg13g2_decap_8 FILLER_66_1975 ();
 sg13g2_fill_1 FILLER_66_1989 ();
 sg13g2_fill_2 FILLER_66_1999 ();
 sg13g2_decap_8 FILLER_66_2023 ();
 sg13g2_decap_8 FILLER_66_2030 ();
 sg13g2_decap_4 FILLER_66_2037 ();
 sg13g2_fill_2 FILLER_66_2041 ();
 sg13g2_fill_2 FILLER_66_2061 ();
 sg13g2_fill_1 FILLER_66_2063 ();
 sg13g2_fill_2 FILLER_66_2069 ();
 sg13g2_fill_1 FILLER_66_2071 ();
 sg13g2_fill_1 FILLER_66_2081 ();
 sg13g2_decap_8 FILLER_66_2109 ();
 sg13g2_decap_8 FILLER_66_2116 ();
 sg13g2_decap_4 FILLER_66_2123 ();
 sg13g2_fill_2 FILLER_66_2137 ();
 sg13g2_fill_1 FILLER_66_2148 ();
 sg13g2_fill_1 FILLER_66_2159 ();
 sg13g2_decap_8 FILLER_66_2173 ();
 sg13g2_decap_4 FILLER_66_2180 ();
 sg13g2_fill_1 FILLER_66_2184 ();
 sg13g2_fill_2 FILLER_66_2196 ();
 sg13g2_fill_1 FILLER_66_2198 ();
 sg13g2_decap_8 FILLER_66_2209 ();
 sg13g2_decap_8 FILLER_66_2216 ();
 sg13g2_decap_4 FILLER_66_2223 ();
 sg13g2_fill_1 FILLER_66_2227 ();
 sg13g2_decap_8 FILLER_66_2236 ();
 sg13g2_fill_1 FILLER_66_2243 ();
 sg13g2_decap_4 FILLER_66_2252 ();
 sg13g2_fill_2 FILLER_66_2256 ();
 sg13g2_decap_4 FILLER_66_2266 ();
 sg13g2_fill_2 FILLER_66_2270 ();
 sg13g2_decap_8 FILLER_66_2287 ();
 sg13g2_fill_2 FILLER_66_2294 ();
 sg13g2_decap_8 FILLER_66_2300 ();
 sg13g2_fill_1 FILLER_66_2307 ();
 sg13g2_decap_4 FILLER_66_2326 ();
 sg13g2_fill_2 FILLER_66_2330 ();
 sg13g2_fill_1 FILLER_66_2346 ();
 sg13g2_fill_2 FILLER_66_2352 ();
 sg13g2_fill_1 FILLER_66_2354 ();
 sg13g2_fill_2 FILLER_66_2376 ();
 sg13g2_decap_4 FILLER_66_2404 ();
 sg13g2_fill_2 FILLER_66_2408 ();
 sg13g2_decap_4 FILLER_66_2418 ();
 sg13g2_fill_1 FILLER_66_2422 ();
 sg13g2_fill_1 FILLER_66_2427 ();
 sg13g2_fill_2 FILLER_66_2437 ();
 sg13g2_fill_1 FILLER_66_2439 ();
 sg13g2_decap_4 FILLER_66_2448 ();
 sg13g2_decap_8 FILLER_66_2490 ();
 sg13g2_fill_1 FILLER_66_2523 ();
 sg13g2_fill_2 FILLER_66_2531 ();
 sg13g2_fill_1 FILLER_66_2537 ();
 sg13g2_fill_2 FILLER_66_2552 ();
 sg13g2_fill_2 FILLER_66_2589 ();
 sg13g2_decap_4 FILLER_66_2611 ();
 sg13g2_fill_1 FILLER_66_2651 ();
 sg13g2_fill_2 FILLER_66_2668 ();
 sg13g2_fill_2 FILLER_66_2699 ();
 sg13g2_fill_1 FILLER_66_2701 ();
 sg13g2_fill_2 FILLER_66_2713 ();
 sg13g2_fill_1 FILLER_66_2715 ();
 sg13g2_decap_4 FILLER_66_2733 ();
 sg13g2_fill_1 FILLER_66_2737 ();
 sg13g2_fill_2 FILLER_66_2755 ();
 sg13g2_fill_1 FILLER_66_2757 ();
 sg13g2_fill_2 FILLER_66_2766 ();
 sg13g2_fill_1 FILLER_66_2768 ();
 sg13g2_decap_8 FILLER_66_2791 ();
 sg13g2_fill_2 FILLER_66_2798 ();
 sg13g2_fill_1 FILLER_66_2800 ();
 sg13g2_decap_4 FILLER_66_2827 ();
 sg13g2_fill_1 FILLER_66_2831 ();
 sg13g2_decap_8 FILLER_66_2837 ();
 sg13g2_fill_2 FILLER_66_2844 ();
 sg13g2_decap_8 FILLER_66_2858 ();
 sg13g2_fill_1 FILLER_66_2865 ();
 sg13g2_fill_2 FILLER_66_2875 ();
 sg13g2_fill_1 FILLER_66_2877 ();
 sg13g2_fill_1 FILLER_66_2901 ();
 sg13g2_decap_8 FILLER_66_2919 ();
 sg13g2_fill_1 FILLER_66_2926 ();
 sg13g2_fill_2 FILLER_66_2946 ();
 sg13g2_fill_1 FILLER_66_2948 ();
 sg13g2_fill_2 FILLER_66_2954 ();
 sg13g2_fill_1 FILLER_66_2956 ();
 sg13g2_decap_8 FILLER_66_2962 ();
 sg13g2_fill_1 FILLER_66_2969 ();
 sg13g2_decap_8 FILLER_66_2974 ();
 sg13g2_fill_2 FILLER_66_2981 ();
 sg13g2_decap_8 FILLER_66_2992 ();
 sg13g2_decap_8 FILLER_66_2999 ();
 sg13g2_decap_8 FILLER_66_3006 ();
 sg13g2_decap_8 FILLER_66_3013 ();
 sg13g2_decap_8 FILLER_66_3020 ();
 sg13g2_decap_8 FILLER_66_3027 ();
 sg13g2_decap_8 FILLER_66_3034 ();
 sg13g2_decap_8 FILLER_66_3041 ();
 sg13g2_decap_8 FILLER_66_3048 ();
 sg13g2_decap_8 FILLER_66_3055 ();
 sg13g2_decap_8 FILLER_66_3062 ();
 sg13g2_decap_8 FILLER_66_3069 ();
 sg13g2_decap_8 FILLER_66_3076 ();
 sg13g2_decap_8 FILLER_66_3083 ();
 sg13g2_decap_8 FILLER_66_3090 ();
 sg13g2_decap_8 FILLER_66_3097 ();
 sg13g2_decap_8 FILLER_66_3104 ();
 sg13g2_decap_8 FILLER_66_3111 ();
 sg13g2_decap_8 FILLER_66_3118 ();
 sg13g2_decap_8 FILLER_66_3125 ();
 sg13g2_decap_8 FILLER_66_3132 ();
 sg13g2_decap_8 FILLER_66_3139 ();
 sg13g2_decap_8 FILLER_66_3146 ();
 sg13g2_decap_8 FILLER_66_3153 ();
 sg13g2_decap_8 FILLER_66_3160 ();
 sg13g2_decap_8 FILLER_66_3167 ();
 sg13g2_decap_8 FILLER_66_3174 ();
 sg13g2_decap_8 FILLER_66_3181 ();
 sg13g2_decap_8 FILLER_66_3188 ();
 sg13g2_decap_8 FILLER_66_3195 ();
 sg13g2_decap_8 FILLER_66_3202 ();
 sg13g2_decap_8 FILLER_66_3209 ();
 sg13g2_decap_8 FILLER_66_3216 ();
 sg13g2_decap_8 FILLER_66_3223 ();
 sg13g2_decap_8 FILLER_66_3230 ();
 sg13g2_decap_8 FILLER_66_3237 ();
 sg13g2_decap_8 FILLER_66_3244 ();
 sg13g2_decap_8 FILLER_66_3251 ();
 sg13g2_decap_8 FILLER_66_3258 ();
 sg13g2_decap_8 FILLER_66_3265 ();
 sg13g2_decap_8 FILLER_66_3272 ();
 sg13g2_decap_8 FILLER_66_3279 ();
 sg13g2_decap_8 FILLER_66_3286 ();
 sg13g2_decap_8 FILLER_66_3293 ();
 sg13g2_decap_8 FILLER_66_3300 ();
 sg13g2_decap_8 FILLER_66_3307 ();
 sg13g2_decap_8 FILLER_66_3314 ();
 sg13g2_decap_8 FILLER_66_3321 ();
 sg13g2_decap_8 FILLER_66_3328 ();
 sg13g2_decap_8 FILLER_66_3335 ();
 sg13g2_decap_8 FILLER_66_3342 ();
 sg13g2_decap_8 FILLER_66_3349 ();
 sg13g2_decap_8 FILLER_66_3356 ();
 sg13g2_decap_8 FILLER_66_3363 ();
 sg13g2_decap_8 FILLER_66_3370 ();
 sg13g2_decap_8 FILLER_66_3377 ();
 sg13g2_decap_8 FILLER_66_3384 ();
 sg13g2_decap_8 FILLER_66_3391 ();
 sg13g2_decap_8 FILLER_66_3398 ();
 sg13g2_decap_8 FILLER_66_3405 ();
 sg13g2_decap_8 FILLER_66_3412 ();
 sg13g2_decap_8 FILLER_66_3419 ();
 sg13g2_decap_8 FILLER_66_3426 ();
 sg13g2_decap_8 FILLER_66_3433 ();
 sg13g2_decap_8 FILLER_66_3440 ();
 sg13g2_decap_8 FILLER_66_3447 ();
 sg13g2_decap_8 FILLER_66_3454 ();
 sg13g2_decap_8 FILLER_66_3461 ();
 sg13g2_decap_8 FILLER_66_3468 ();
 sg13g2_decap_8 FILLER_66_3475 ();
 sg13g2_decap_8 FILLER_66_3482 ();
 sg13g2_decap_8 FILLER_66_3489 ();
 sg13g2_decap_8 FILLER_66_3496 ();
 sg13g2_decap_8 FILLER_66_3503 ();
 sg13g2_decap_8 FILLER_66_3510 ();
 sg13g2_decap_8 FILLER_66_3517 ();
 sg13g2_decap_8 FILLER_66_3524 ();
 sg13g2_decap_8 FILLER_66_3531 ();
 sg13g2_decap_8 FILLER_66_3538 ();
 sg13g2_decap_8 FILLER_66_3545 ();
 sg13g2_decap_8 FILLER_66_3552 ();
 sg13g2_decap_8 FILLER_66_3559 ();
 sg13g2_decap_8 FILLER_66_3566 ();
 sg13g2_decap_8 FILLER_66_3573 ();
 sg13g2_fill_2 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_fill_2 FILLER_67_77 ();
 sg13g2_fill_2 FILLER_67_89 ();
 sg13g2_decap_4 FILLER_67_117 ();
 sg13g2_fill_2 FILLER_67_131 ();
 sg13g2_decap_8 FILLER_67_138 ();
 sg13g2_fill_1 FILLER_67_145 ();
 sg13g2_decap_8 FILLER_67_169 ();
 sg13g2_decap_8 FILLER_67_176 ();
 sg13g2_fill_1 FILLER_67_183 ();
 sg13g2_decap_4 FILLER_67_190 ();
 sg13g2_fill_1 FILLER_67_194 ();
 sg13g2_decap_4 FILLER_67_204 ();
 sg13g2_fill_2 FILLER_67_208 ();
 sg13g2_decap_8 FILLER_67_214 ();
 sg13g2_decap_4 FILLER_67_221 ();
 sg13g2_fill_1 FILLER_67_225 ();
 sg13g2_fill_2 FILLER_67_252 ();
 sg13g2_decap_8 FILLER_67_281 ();
 sg13g2_decap_8 FILLER_67_288 ();
 sg13g2_decap_4 FILLER_67_295 ();
 sg13g2_decap_8 FILLER_67_329 ();
 sg13g2_fill_1 FILLER_67_336 ();
 sg13g2_decap_8 FILLER_67_341 ();
 sg13g2_decap_4 FILLER_67_348 ();
 sg13g2_fill_1 FILLER_67_352 ();
 sg13g2_fill_1 FILLER_67_358 ();
 sg13g2_fill_1 FILLER_67_402 ();
 sg13g2_fill_2 FILLER_67_421 ();
 sg13g2_fill_1 FILLER_67_445 ();
 sg13g2_fill_2 FILLER_67_487 ();
 sg13g2_fill_1 FILLER_67_489 ();
 sg13g2_fill_2 FILLER_67_499 ();
 sg13g2_fill_1 FILLER_67_506 ();
 sg13g2_fill_2 FILLER_67_512 ();
 sg13g2_fill_2 FILLER_67_525 ();
 sg13g2_fill_1 FILLER_67_527 ();
 sg13g2_fill_2 FILLER_67_536 ();
 sg13g2_fill_1 FILLER_67_538 ();
 sg13g2_decap_4 FILLER_67_561 ();
 sg13g2_decap_8 FILLER_67_591 ();
 sg13g2_fill_2 FILLER_67_598 ();
 sg13g2_fill_1 FILLER_67_633 ();
 sg13g2_fill_2 FILLER_67_702 ();
 sg13g2_fill_2 FILLER_67_713 ();
 sg13g2_fill_1 FILLER_67_715 ();
 sg13g2_fill_2 FILLER_67_734 ();
 sg13g2_fill_2 FILLER_67_872 ();
 sg13g2_fill_1 FILLER_67_874 ();
 sg13g2_decap_8 FILLER_67_879 ();
 sg13g2_decap_8 FILLER_67_903 ();
 sg13g2_fill_2 FILLER_67_910 ();
 sg13g2_fill_1 FILLER_67_912 ();
 sg13g2_fill_2 FILLER_67_926 ();
 sg13g2_fill_1 FILLER_67_928 ();
 sg13g2_decap_8 FILLER_67_969 ();
 sg13g2_fill_1 FILLER_67_976 ();
 sg13g2_fill_2 FILLER_67_989 ();
 sg13g2_fill_1 FILLER_67_991 ();
 sg13g2_decap_8 FILLER_67_997 ();
 sg13g2_fill_2 FILLER_67_1004 ();
 sg13g2_fill_2 FILLER_67_1009 ();
 sg13g2_fill_1 FILLER_67_1011 ();
 sg13g2_fill_2 FILLER_67_1043 ();
 sg13g2_fill_1 FILLER_67_1045 ();
 sg13g2_fill_2 FILLER_67_1060 ();
 sg13g2_fill_2 FILLER_67_1071 ();
 sg13g2_fill_2 FILLER_67_1116 ();
 sg13g2_fill_2 FILLER_67_1163 ();
 sg13g2_decap_4 FILLER_67_1178 ();
 sg13g2_fill_1 FILLER_67_1182 ();
 sg13g2_fill_2 FILLER_67_1220 ();
 sg13g2_fill_1 FILLER_67_1227 ();
 sg13g2_fill_2 FILLER_67_1266 ();
 sg13g2_fill_1 FILLER_67_1291 ();
 sg13g2_decap_8 FILLER_67_1346 ();
 sg13g2_decap_8 FILLER_67_1353 ();
 sg13g2_decap_8 FILLER_67_1360 ();
 sg13g2_decap_4 FILLER_67_1367 ();
 sg13g2_decap_4 FILLER_67_1388 ();
 sg13g2_fill_2 FILLER_67_1392 ();
 sg13g2_fill_2 FILLER_67_1413 ();
 sg13g2_fill_1 FILLER_67_1415 ();
 sg13g2_fill_2 FILLER_67_1425 ();
 sg13g2_fill_2 FILLER_67_1517 ();
 sg13g2_fill_1 FILLER_67_1519 ();
 sg13g2_fill_1 FILLER_67_1529 ();
 sg13g2_fill_2 FILLER_67_1560 ();
 sg13g2_fill_2 FILLER_67_1585 ();
 sg13g2_fill_1 FILLER_67_1587 ();
 sg13g2_fill_2 FILLER_67_1597 ();
 sg13g2_fill_1 FILLER_67_1599 ();
 sg13g2_fill_2 FILLER_67_1625 ();
 sg13g2_fill_1 FILLER_67_1636 ();
 sg13g2_decap_8 FILLER_67_1681 ();
 sg13g2_fill_2 FILLER_67_1688 ();
 sg13g2_fill_1 FILLER_67_1690 ();
 sg13g2_fill_1 FILLER_67_1706 ();
 sg13g2_fill_2 FILLER_67_1717 ();
 sg13g2_decap_4 FILLER_67_1745 ();
 sg13g2_fill_1 FILLER_67_1749 ();
 sg13g2_decap_4 FILLER_67_1763 ();
 sg13g2_fill_1 FILLER_67_1767 ();
 sg13g2_fill_2 FILLER_67_1792 ();
 sg13g2_fill_1 FILLER_67_1794 ();
 sg13g2_fill_2 FILLER_67_1833 ();
 sg13g2_fill_1 FILLER_67_1835 ();
 sg13g2_fill_2 FILLER_67_1844 ();
 sg13g2_fill_1 FILLER_67_1846 ();
 sg13g2_fill_1 FILLER_67_1852 ();
 sg13g2_fill_1 FILLER_67_1863 ();
 sg13g2_decap_4 FILLER_67_1875 ();
 sg13g2_decap_4 FILLER_67_1899 ();
 sg13g2_fill_1 FILLER_67_1903 ();
 sg13g2_fill_1 FILLER_67_1915 ();
 sg13g2_decap_4 FILLER_67_1929 ();
 sg13g2_fill_1 FILLER_67_1933 ();
 sg13g2_decap_4 FILLER_67_1940 ();
 sg13g2_fill_1 FILLER_67_1944 ();
 sg13g2_fill_2 FILLER_67_1954 ();
 sg13g2_decap_8 FILLER_67_1979 ();
 sg13g2_fill_2 FILLER_67_1986 ();
 sg13g2_fill_1 FILLER_67_1988 ();
 sg13g2_fill_1 FILLER_67_2012 ();
 sg13g2_decap_8 FILLER_67_2017 ();
 sg13g2_decap_8 FILLER_67_2024 ();
 sg13g2_fill_1 FILLER_67_2035 ();
 sg13g2_decap_8 FILLER_67_2044 ();
 sg13g2_decap_4 FILLER_67_2051 ();
 sg13g2_fill_2 FILLER_67_2064 ();
 sg13g2_fill_1 FILLER_67_2066 ();
 sg13g2_decap_8 FILLER_67_2075 ();
 sg13g2_decap_8 FILLER_67_2082 ();
 sg13g2_decap_4 FILLER_67_2089 ();
 sg13g2_decap_8 FILLER_67_2103 ();
 sg13g2_decap_4 FILLER_67_2110 ();
 sg13g2_fill_1 FILLER_67_2114 ();
 sg13g2_fill_1 FILLER_67_2138 ();
 sg13g2_fill_1 FILLER_67_2152 ();
 sg13g2_fill_2 FILLER_67_2158 ();
 sg13g2_fill_1 FILLER_67_2160 ();
 sg13g2_fill_1 FILLER_67_2204 ();
 sg13g2_fill_2 FILLER_67_2231 ();
 sg13g2_fill_1 FILLER_67_2233 ();
 sg13g2_decap_8 FILLER_67_2256 ();
 sg13g2_decap_4 FILLER_67_2263 ();
 sg13g2_fill_1 FILLER_67_2267 ();
 sg13g2_decap_8 FILLER_67_2286 ();
 sg13g2_fill_1 FILLER_67_2293 ();
 sg13g2_fill_2 FILLER_67_2314 ();
 sg13g2_fill_1 FILLER_67_2316 ();
 sg13g2_fill_1 FILLER_67_2344 ();
 sg13g2_fill_2 FILLER_67_2350 ();
 sg13g2_fill_1 FILLER_67_2352 ();
 sg13g2_decap_4 FILLER_67_2379 ();
 sg13g2_decap_8 FILLER_67_2396 ();
 sg13g2_fill_1 FILLER_67_2403 ();
 sg13g2_fill_2 FILLER_67_2435 ();
 sg13g2_fill_1 FILLER_67_2437 ();
 sg13g2_decap_4 FILLER_67_2444 ();
 sg13g2_fill_2 FILLER_67_2466 ();
 sg13g2_fill_1 FILLER_67_2487 ();
 sg13g2_decap_8 FILLER_67_2492 ();
 sg13g2_decap_8 FILLER_67_2499 ();
 sg13g2_fill_2 FILLER_67_2506 ();
 sg13g2_fill_1 FILLER_67_2508 ();
 sg13g2_fill_1 FILLER_67_2574 ();
 sg13g2_decap_4 FILLER_67_2579 ();
 sg13g2_fill_1 FILLER_67_2583 ();
 sg13g2_fill_2 FILLER_67_2593 ();
 sg13g2_decap_8 FILLER_67_2602 ();
 sg13g2_decap_8 FILLER_67_2609 ();
 sg13g2_decap_8 FILLER_67_2616 ();
 sg13g2_fill_1 FILLER_67_2623 ();
 sg13g2_decap_8 FILLER_67_2637 ();
 sg13g2_decap_8 FILLER_67_2644 ();
 sg13g2_decap_4 FILLER_67_2651 ();
 sg13g2_fill_1 FILLER_67_2655 ();
 sg13g2_decap_8 FILLER_67_2660 ();
 sg13g2_decap_8 FILLER_67_2667 ();
 sg13g2_decap_4 FILLER_67_2674 ();
 sg13g2_fill_2 FILLER_67_2678 ();
 sg13g2_fill_1 FILLER_67_2696 ();
 sg13g2_decap_8 FILLER_67_2701 ();
 sg13g2_decap_8 FILLER_67_2708 ();
 sg13g2_fill_2 FILLER_67_2715 ();
 sg13g2_fill_1 FILLER_67_2717 ();
 sg13g2_decap_8 FILLER_67_2731 ();
 sg13g2_decap_8 FILLER_67_2755 ();
 sg13g2_decap_8 FILLER_67_2762 ();
 sg13g2_decap_4 FILLER_67_2769 ();
 sg13g2_decap_8 FILLER_67_2791 ();
 sg13g2_decap_8 FILLER_67_2798 ();
 sg13g2_decap_8 FILLER_67_2820 ();
 sg13g2_fill_1 FILLER_67_2827 ();
 sg13g2_decap_8 FILLER_67_2833 ();
 sg13g2_fill_1 FILLER_67_2840 ();
 sg13g2_fill_2 FILLER_67_2865 ();
 sg13g2_fill_1 FILLER_67_2867 ();
 sg13g2_decap_4 FILLER_67_2885 ();
 sg13g2_fill_2 FILLER_67_2889 ();
 sg13g2_decap_8 FILLER_67_2895 ();
 sg13g2_decap_8 FILLER_67_2922 ();
 sg13g2_fill_2 FILLER_67_2929 ();
 sg13g2_fill_1 FILLER_67_2931 ();
 sg13g2_decap_4 FILLER_67_2935 ();
 sg13g2_fill_1 FILLER_67_2958 ();
 sg13g2_decap_8 FILLER_67_2985 ();
 sg13g2_decap_8 FILLER_67_2992 ();
 sg13g2_decap_8 FILLER_67_2999 ();
 sg13g2_decap_8 FILLER_67_3006 ();
 sg13g2_decap_8 FILLER_67_3013 ();
 sg13g2_decap_8 FILLER_67_3020 ();
 sg13g2_decap_8 FILLER_67_3027 ();
 sg13g2_decap_8 FILLER_67_3034 ();
 sg13g2_decap_8 FILLER_67_3041 ();
 sg13g2_decap_8 FILLER_67_3048 ();
 sg13g2_decap_8 FILLER_67_3055 ();
 sg13g2_decap_8 FILLER_67_3062 ();
 sg13g2_decap_8 FILLER_67_3069 ();
 sg13g2_decap_8 FILLER_67_3076 ();
 sg13g2_decap_8 FILLER_67_3083 ();
 sg13g2_decap_8 FILLER_67_3090 ();
 sg13g2_decap_8 FILLER_67_3097 ();
 sg13g2_decap_8 FILLER_67_3104 ();
 sg13g2_decap_8 FILLER_67_3111 ();
 sg13g2_decap_8 FILLER_67_3118 ();
 sg13g2_decap_8 FILLER_67_3125 ();
 sg13g2_decap_8 FILLER_67_3132 ();
 sg13g2_decap_8 FILLER_67_3139 ();
 sg13g2_decap_8 FILLER_67_3146 ();
 sg13g2_decap_8 FILLER_67_3153 ();
 sg13g2_decap_8 FILLER_67_3160 ();
 sg13g2_decap_8 FILLER_67_3167 ();
 sg13g2_decap_8 FILLER_67_3174 ();
 sg13g2_decap_8 FILLER_67_3181 ();
 sg13g2_decap_8 FILLER_67_3188 ();
 sg13g2_decap_8 FILLER_67_3195 ();
 sg13g2_decap_8 FILLER_67_3202 ();
 sg13g2_decap_8 FILLER_67_3209 ();
 sg13g2_decap_8 FILLER_67_3216 ();
 sg13g2_decap_8 FILLER_67_3223 ();
 sg13g2_decap_8 FILLER_67_3230 ();
 sg13g2_decap_8 FILLER_67_3237 ();
 sg13g2_decap_8 FILLER_67_3244 ();
 sg13g2_decap_8 FILLER_67_3251 ();
 sg13g2_decap_8 FILLER_67_3258 ();
 sg13g2_decap_8 FILLER_67_3265 ();
 sg13g2_decap_8 FILLER_67_3272 ();
 sg13g2_decap_8 FILLER_67_3279 ();
 sg13g2_decap_8 FILLER_67_3286 ();
 sg13g2_decap_8 FILLER_67_3293 ();
 sg13g2_decap_8 FILLER_67_3300 ();
 sg13g2_decap_8 FILLER_67_3307 ();
 sg13g2_decap_8 FILLER_67_3314 ();
 sg13g2_decap_8 FILLER_67_3321 ();
 sg13g2_decap_8 FILLER_67_3328 ();
 sg13g2_decap_8 FILLER_67_3335 ();
 sg13g2_decap_8 FILLER_67_3342 ();
 sg13g2_decap_8 FILLER_67_3349 ();
 sg13g2_decap_8 FILLER_67_3356 ();
 sg13g2_decap_8 FILLER_67_3363 ();
 sg13g2_decap_8 FILLER_67_3370 ();
 sg13g2_decap_8 FILLER_67_3377 ();
 sg13g2_decap_8 FILLER_67_3384 ();
 sg13g2_decap_8 FILLER_67_3391 ();
 sg13g2_decap_8 FILLER_67_3398 ();
 sg13g2_decap_8 FILLER_67_3405 ();
 sg13g2_decap_8 FILLER_67_3412 ();
 sg13g2_decap_8 FILLER_67_3419 ();
 sg13g2_decap_8 FILLER_67_3426 ();
 sg13g2_decap_8 FILLER_67_3433 ();
 sg13g2_decap_8 FILLER_67_3440 ();
 sg13g2_decap_8 FILLER_67_3447 ();
 sg13g2_decap_8 FILLER_67_3454 ();
 sg13g2_decap_8 FILLER_67_3461 ();
 sg13g2_decap_8 FILLER_67_3468 ();
 sg13g2_decap_8 FILLER_67_3475 ();
 sg13g2_decap_8 FILLER_67_3482 ();
 sg13g2_decap_8 FILLER_67_3489 ();
 sg13g2_decap_8 FILLER_67_3496 ();
 sg13g2_decap_8 FILLER_67_3503 ();
 sg13g2_decap_8 FILLER_67_3510 ();
 sg13g2_decap_8 FILLER_67_3517 ();
 sg13g2_decap_8 FILLER_67_3524 ();
 sg13g2_decap_8 FILLER_67_3531 ();
 sg13g2_decap_8 FILLER_67_3538 ();
 sg13g2_decap_8 FILLER_67_3545 ();
 sg13g2_decap_8 FILLER_67_3552 ();
 sg13g2_decap_8 FILLER_67_3559 ();
 sg13g2_decap_8 FILLER_67_3566 ();
 sg13g2_decap_8 FILLER_67_3573 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_4 FILLER_68_7 ();
 sg13g2_decap_4 FILLER_68_15 ();
 sg13g2_fill_2 FILLER_68_19 ();
 sg13g2_fill_2 FILLER_68_38 ();
 sg13g2_fill_1 FILLER_68_40 ();
 sg13g2_fill_2 FILLER_68_68 ();
 sg13g2_fill_2 FILLER_68_82 ();
 sg13g2_fill_1 FILLER_68_94 ();
 sg13g2_decap_4 FILLER_68_158 ();
 sg13g2_fill_2 FILLER_68_197 ();
 sg13g2_fill_2 FILLER_68_235 ();
 sg13g2_fill_2 FILLER_68_250 ();
 sg13g2_fill_2 FILLER_68_262 ();
 sg13g2_fill_1 FILLER_68_269 ();
 sg13g2_fill_2 FILLER_68_279 ();
 sg13g2_fill_1 FILLER_68_281 ();
 sg13g2_decap_4 FILLER_68_291 ();
 sg13g2_fill_1 FILLER_68_318 ();
 sg13g2_decap_4 FILLER_68_328 ();
 sg13g2_fill_1 FILLER_68_332 ();
 sg13g2_fill_2 FILLER_68_362 ();
 sg13g2_fill_2 FILLER_68_369 ();
 sg13g2_fill_1 FILLER_68_371 ();
 sg13g2_fill_2 FILLER_68_381 ();
 sg13g2_fill_1 FILLER_68_383 ();
 sg13g2_fill_1 FILLER_68_424 ();
 sg13g2_fill_2 FILLER_68_428 ();
 sg13g2_fill_1 FILLER_68_430 ();
 sg13g2_fill_1 FILLER_68_492 ();
 sg13g2_decap_4 FILLER_68_507 ();
 sg13g2_fill_2 FILLER_68_511 ();
 sg13g2_fill_2 FILLER_68_546 ();
 sg13g2_fill_1 FILLER_68_548 ();
 sg13g2_decap_4 FILLER_68_564 ();
 sg13g2_fill_2 FILLER_68_568 ();
 sg13g2_decap_4 FILLER_68_574 ();
 sg13g2_fill_2 FILLER_68_578 ();
 sg13g2_decap_4 FILLER_68_585 ();
 sg13g2_fill_1 FILLER_68_589 ();
 sg13g2_fill_1 FILLER_68_616 ();
 sg13g2_fill_2 FILLER_68_676 ();
 sg13g2_decap_4 FILLER_68_688 ();
 sg13g2_fill_2 FILLER_68_692 ();
 sg13g2_decap_4 FILLER_68_725 ();
 sg13g2_fill_1 FILLER_68_760 ();
 sg13g2_decap_4 FILLER_68_765 ();
 sg13g2_fill_1 FILLER_68_769 ();
 sg13g2_fill_1 FILLER_68_787 ();
 sg13g2_fill_2 FILLER_68_794 ();
 sg13g2_fill_1 FILLER_68_801 ();
 sg13g2_decap_8 FILLER_68_809 ();
 sg13g2_decap_8 FILLER_68_816 ();
 sg13g2_fill_2 FILLER_68_823 ();
 sg13g2_fill_1 FILLER_68_844 ();
 sg13g2_fill_2 FILLER_68_927 ();
 sg13g2_fill_1 FILLER_68_929 ();
 sg13g2_fill_2 FILLER_68_953 ();
 sg13g2_fill_1 FILLER_68_955 ();
 sg13g2_fill_1 FILLER_68_970 ();
 sg13g2_fill_2 FILLER_68_1030 ();
 sg13g2_fill_1 FILLER_68_1032 ();
 sg13g2_fill_2 FILLER_68_1043 ();
 sg13g2_fill_1 FILLER_68_1045 ();
 sg13g2_fill_1 FILLER_68_1070 ();
 sg13g2_decap_4 FILLER_68_1092 ();
 sg13g2_fill_2 FILLER_68_1122 ();
 sg13g2_decap_8 FILLER_68_1152 ();
 sg13g2_fill_1 FILLER_68_1159 ();
 sg13g2_decap_4 FILLER_68_1167 ();
 sg13g2_fill_1 FILLER_68_1204 ();
 sg13g2_fill_2 FILLER_68_1214 ();
 sg13g2_fill_1 FILLER_68_1216 ();
 sg13g2_fill_2 FILLER_68_1222 ();
 sg13g2_fill_1 FILLER_68_1224 ();
 sg13g2_fill_2 FILLER_68_1229 ();
 sg13g2_fill_2 FILLER_68_1236 ();
 sg13g2_fill_1 FILLER_68_1238 ();
 sg13g2_fill_2 FILLER_68_1246 ();
 sg13g2_fill_1 FILLER_68_1248 ();
 sg13g2_decap_4 FILLER_68_1253 ();
 sg13g2_fill_2 FILLER_68_1257 ();
 sg13g2_decap_4 FILLER_68_1291 ();
 sg13g2_fill_1 FILLER_68_1295 ();
 sg13g2_fill_1 FILLER_68_1301 ();
 sg13g2_fill_1 FILLER_68_1311 ();
 sg13g2_decap_8 FILLER_68_1325 ();
 sg13g2_fill_1 FILLER_68_1332 ();
 sg13g2_decap_4 FILLER_68_1360 ();
 sg13g2_fill_1 FILLER_68_1364 ();
 sg13g2_decap_8 FILLER_68_1389 ();
 sg13g2_fill_2 FILLER_68_1396 ();
 sg13g2_fill_1 FILLER_68_1407 ();
 sg13g2_fill_2 FILLER_68_1426 ();
 sg13g2_fill_2 FILLER_68_1459 ();
 sg13g2_decap_4 FILLER_68_1469 ();
 sg13g2_fill_2 FILLER_68_1473 ();
 sg13g2_fill_2 FILLER_68_1488 ();
 sg13g2_fill_2 FILLER_68_1504 ();
 sg13g2_fill_2 FILLER_68_1532 ();
 sg13g2_fill_1 FILLER_68_1534 ();
 sg13g2_fill_1 FILLER_68_1558 ();
 sg13g2_fill_2 FILLER_68_1564 ();
 sg13g2_fill_1 FILLER_68_1566 ();
 sg13g2_fill_2 FILLER_68_1605 ();
 sg13g2_fill_1 FILLER_68_1632 ();
 sg13g2_fill_2 FILLER_68_1642 ();
 sg13g2_fill_1 FILLER_68_1644 ();
 sg13g2_decap_4 FILLER_68_1690 ();
 sg13g2_fill_1 FILLER_68_1694 ();
 sg13g2_decap_4 FILLER_68_1699 ();
 sg13g2_fill_2 FILLER_68_1712 ();
 sg13g2_fill_1 FILLER_68_1714 ();
 sg13g2_decap_4 FILLER_68_1741 ();
 sg13g2_fill_1 FILLER_68_1755 ();
 sg13g2_fill_1 FILLER_68_1774 ();
 sg13g2_decap_8 FILLER_68_1806 ();
 sg13g2_fill_1 FILLER_68_1839 ();
 sg13g2_fill_2 FILLER_68_1849 ();
 sg13g2_fill_2 FILLER_68_1856 ();
 sg13g2_decap_8 FILLER_68_1886 ();
 sg13g2_fill_1 FILLER_68_1893 ();
 sg13g2_fill_2 FILLER_68_1899 ();
 sg13g2_fill_1 FILLER_68_1901 ();
 sg13g2_decap_8 FILLER_68_1925 ();
 sg13g2_fill_1 FILLER_68_1932 ();
 sg13g2_fill_1 FILLER_68_1942 ();
 sg13g2_decap_8 FILLER_68_1965 ();
 sg13g2_decap_4 FILLER_68_1972 ();
 sg13g2_fill_2 FILLER_68_1990 ();
 sg13g2_decap_8 FILLER_68_2005 ();
 sg13g2_decap_4 FILLER_68_2016 ();
 sg13g2_decap_8 FILLER_68_2046 ();
 sg13g2_decap_4 FILLER_68_2053 ();
 sg13g2_fill_1 FILLER_68_2057 ();
 sg13g2_decap_8 FILLER_68_2072 ();
 sg13g2_decap_4 FILLER_68_2079 ();
 sg13g2_fill_2 FILLER_68_2083 ();
 sg13g2_decap_8 FILLER_68_2093 ();
 sg13g2_decap_4 FILLER_68_2100 ();
 sg13g2_fill_2 FILLER_68_2122 ();
 sg13g2_fill_1 FILLER_68_2161 ();
 sg13g2_decap_8 FILLER_68_2196 ();
 sg13g2_decap_4 FILLER_68_2208 ();
 sg13g2_fill_2 FILLER_68_2212 ();
 sg13g2_decap_8 FILLER_68_2237 ();
 sg13g2_fill_2 FILLER_68_2244 ();
 sg13g2_fill_2 FILLER_68_2313 ();
 sg13g2_fill_1 FILLER_68_2319 ();
 sg13g2_fill_2 FILLER_68_2325 ();
 sg13g2_fill_1 FILLER_68_2327 ();
 sg13g2_decap_4 FILLER_68_2338 ();
 sg13g2_fill_2 FILLER_68_2342 ();
 sg13g2_fill_1 FILLER_68_2358 ();
 sg13g2_fill_2 FILLER_68_2372 ();
 sg13g2_fill_1 FILLER_68_2374 ();
 sg13g2_fill_1 FILLER_68_2409 ();
 sg13g2_fill_1 FILLER_68_2419 ();
 sg13g2_decap_8 FILLER_68_2475 ();
 sg13g2_decap_8 FILLER_68_2482 ();
 sg13g2_decap_8 FILLER_68_2494 ();
 sg13g2_decap_4 FILLER_68_2501 ();
 sg13g2_fill_1 FILLER_68_2505 ();
 sg13g2_fill_2 FILLER_68_2511 ();
 sg13g2_decap_8 FILLER_68_2517 ();
 sg13g2_decap_8 FILLER_68_2524 ();
 sg13g2_decap_8 FILLER_68_2531 ();
 sg13g2_fill_2 FILLER_68_2538 ();
 sg13g2_fill_1 FILLER_68_2540 ();
 sg13g2_decap_8 FILLER_68_2544 ();
 sg13g2_fill_2 FILLER_68_2551 ();
 sg13g2_decap_8 FILLER_68_2557 ();
 sg13g2_fill_2 FILLER_68_2564 ();
 sg13g2_fill_2 FILLER_68_2609 ();
 sg13g2_fill_1 FILLER_68_2611 ();
 sg13g2_fill_1 FILLER_68_2647 ();
 sg13g2_fill_1 FILLER_68_2656 ();
 sg13g2_fill_1 FILLER_68_2666 ();
 sg13g2_fill_2 FILLER_68_2672 ();
 sg13g2_fill_1 FILLER_68_2674 ();
 sg13g2_decap_8 FILLER_68_2684 ();
 sg13g2_fill_2 FILLER_68_2691 ();
 sg13g2_fill_1 FILLER_68_2693 ();
 sg13g2_decap_8 FILLER_68_2714 ();
 sg13g2_fill_2 FILLER_68_2721 ();
 sg13g2_fill_1 FILLER_68_2736 ();
 sg13g2_fill_2 FILLER_68_2745 ();
 sg13g2_decap_8 FILLER_68_2763 ();
 sg13g2_fill_2 FILLER_68_2770 ();
 sg13g2_decap_8 FILLER_68_2776 ();
 sg13g2_fill_2 FILLER_68_2783 ();
 sg13g2_decap_4 FILLER_68_2795 ();
 sg13g2_fill_2 FILLER_68_2856 ();
 sg13g2_decap_8 FILLER_68_2863 ();
 sg13g2_fill_2 FILLER_68_2870 ();
 sg13g2_fill_1 FILLER_68_2872 ();
 sg13g2_decap_8 FILLER_68_2889 ();
 sg13g2_decap_8 FILLER_68_2896 ();
 sg13g2_decap_4 FILLER_68_2917 ();
 sg13g2_fill_2 FILLER_68_2921 ();
 sg13g2_decap_8 FILLER_68_2941 ();
 sg13g2_decap_8 FILLER_68_2948 ();
 sg13g2_fill_2 FILLER_68_2955 ();
 sg13g2_decap_8 FILLER_68_2960 ();
 sg13g2_decap_4 FILLER_68_2967 ();
 sg13g2_fill_1 FILLER_68_2971 ();
 sg13g2_decap_8 FILLER_68_2981 ();
 sg13g2_decap_8 FILLER_68_2988 ();
 sg13g2_decap_8 FILLER_68_2995 ();
 sg13g2_decap_8 FILLER_68_3002 ();
 sg13g2_decap_8 FILLER_68_3009 ();
 sg13g2_decap_8 FILLER_68_3016 ();
 sg13g2_decap_8 FILLER_68_3023 ();
 sg13g2_decap_8 FILLER_68_3030 ();
 sg13g2_decap_8 FILLER_68_3037 ();
 sg13g2_decap_8 FILLER_68_3044 ();
 sg13g2_decap_8 FILLER_68_3051 ();
 sg13g2_decap_8 FILLER_68_3058 ();
 sg13g2_decap_8 FILLER_68_3065 ();
 sg13g2_decap_8 FILLER_68_3072 ();
 sg13g2_decap_8 FILLER_68_3079 ();
 sg13g2_decap_8 FILLER_68_3086 ();
 sg13g2_decap_8 FILLER_68_3093 ();
 sg13g2_decap_8 FILLER_68_3100 ();
 sg13g2_decap_8 FILLER_68_3107 ();
 sg13g2_decap_8 FILLER_68_3114 ();
 sg13g2_decap_8 FILLER_68_3121 ();
 sg13g2_decap_8 FILLER_68_3128 ();
 sg13g2_decap_8 FILLER_68_3135 ();
 sg13g2_decap_8 FILLER_68_3142 ();
 sg13g2_decap_8 FILLER_68_3149 ();
 sg13g2_decap_8 FILLER_68_3156 ();
 sg13g2_decap_8 FILLER_68_3163 ();
 sg13g2_decap_8 FILLER_68_3170 ();
 sg13g2_decap_8 FILLER_68_3177 ();
 sg13g2_decap_8 FILLER_68_3184 ();
 sg13g2_decap_8 FILLER_68_3191 ();
 sg13g2_decap_8 FILLER_68_3198 ();
 sg13g2_decap_8 FILLER_68_3205 ();
 sg13g2_decap_8 FILLER_68_3212 ();
 sg13g2_decap_8 FILLER_68_3219 ();
 sg13g2_decap_8 FILLER_68_3226 ();
 sg13g2_decap_8 FILLER_68_3233 ();
 sg13g2_decap_8 FILLER_68_3240 ();
 sg13g2_decap_8 FILLER_68_3247 ();
 sg13g2_decap_8 FILLER_68_3254 ();
 sg13g2_decap_8 FILLER_68_3261 ();
 sg13g2_decap_8 FILLER_68_3268 ();
 sg13g2_decap_8 FILLER_68_3275 ();
 sg13g2_decap_8 FILLER_68_3282 ();
 sg13g2_decap_8 FILLER_68_3289 ();
 sg13g2_decap_8 FILLER_68_3296 ();
 sg13g2_decap_8 FILLER_68_3303 ();
 sg13g2_decap_8 FILLER_68_3310 ();
 sg13g2_decap_8 FILLER_68_3317 ();
 sg13g2_decap_8 FILLER_68_3324 ();
 sg13g2_decap_8 FILLER_68_3331 ();
 sg13g2_decap_8 FILLER_68_3338 ();
 sg13g2_decap_8 FILLER_68_3345 ();
 sg13g2_decap_8 FILLER_68_3352 ();
 sg13g2_decap_8 FILLER_68_3359 ();
 sg13g2_decap_8 FILLER_68_3366 ();
 sg13g2_decap_8 FILLER_68_3373 ();
 sg13g2_decap_8 FILLER_68_3380 ();
 sg13g2_decap_8 FILLER_68_3387 ();
 sg13g2_decap_8 FILLER_68_3394 ();
 sg13g2_decap_8 FILLER_68_3401 ();
 sg13g2_decap_8 FILLER_68_3408 ();
 sg13g2_decap_8 FILLER_68_3415 ();
 sg13g2_decap_8 FILLER_68_3422 ();
 sg13g2_decap_8 FILLER_68_3429 ();
 sg13g2_decap_8 FILLER_68_3436 ();
 sg13g2_decap_8 FILLER_68_3443 ();
 sg13g2_decap_8 FILLER_68_3450 ();
 sg13g2_decap_8 FILLER_68_3457 ();
 sg13g2_decap_8 FILLER_68_3464 ();
 sg13g2_decap_8 FILLER_68_3471 ();
 sg13g2_decap_8 FILLER_68_3478 ();
 sg13g2_decap_8 FILLER_68_3485 ();
 sg13g2_decap_8 FILLER_68_3492 ();
 sg13g2_decap_8 FILLER_68_3499 ();
 sg13g2_decap_8 FILLER_68_3506 ();
 sg13g2_decap_8 FILLER_68_3513 ();
 sg13g2_decap_8 FILLER_68_3520 ();
 sg13g2_decap_8 FILLER_68_3527 ();
 sg13g2_decap_8 FILLER_68_3534 ();
 sg13g2_decap_8 FILLER_68_3541 ();
 sg13g2_decap_8 FILLER_68_3548 ();
 sg13g2_decap_8 FILLER_68_3555 ();
 sg13g2_decap_8 FILLER_68_3562 ();
 sg13g2_decap_8 FILLER_68_3569 ();
 sg13g2_decap_4 FILLER_68_3576 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_fill_1 FILLER_69_14 ();
 sg13g2_fill_2 FILLER_69_113 ();
 sg13g2_fill_1 FILLER_69_115 ();
 sg13g2_fill_2 FILLER_69_121 ();
 sg13g2_decap_8 FILLER_69_140 ();
 sg13g2_decap_4 FILLER_69_147 ();
 sg13g2_fill_1 FILLER_69_151 ();
 sg13g2_decap_4 FILLER_69_167 ();
 sg13g2_fill_2 FILLER_69_171 ();
 sg13g2_decap_4 FILLER_69_177 ();
 sg13g2_decap_8 FILLER_69_191 ();
 sg13g2_decap_8 FILLER_69_198 ();
 sg13g2_fill_1 FILLER_69_205 ();
 sg13g2_fill_2 FILLER_69_237 ();
 sg13g2_fill_1 FILLER_69_239 ();
 sg13g2_fill_2 FILLER_69_258 ();
 sg13g2_fill_2 FILLER_69_295 ();
 sg13g2_decap_8 FILLER_69_341 ();
 sg13g2_fill_2 FILLER_69_376 ();
 sg13g2_fill_2 FILLER_69_383 ();
 sg13g2_fill_1 FILLER_69_385 ();
 sg13g2_decap_4 FILLER_69_431 ();
 sg13g2_fill_2 FILLER_69_440 ();
 sg13g2_decap_8 FILLER_69_451 ();
 sg13g2_decap_4 FILLER_69_458 ();
 sg13g2_fill_1 FILLER_69_462 ();
 sg13g2_decap_8 FILLER_69_468 ();
 sg13g2_fill_1 FILLER_69_475 ();
 sg13g2_fill_2 FILLER_69_493 ();
 sg13g2_fill_1 FILLER_69_495 ();
 sg13g2_fill_2 FILLER_69_529 ();
 sg13g2_fill_2 FILLER_69_557 ();
 sg13g2_decap_8 FILLER_69_598 ();
 sg13g2_decap_4 FILLER_69_605 ();
 sg13g2_fill_2 FILLER_69_639 ();
 sg13g2_decap_4 FILLER_69_746 ();
 sg13g2_fill_2 FILLER_69_785 ();
 sg13g2_fill_2 FILLER_69_807 ();
 sg13g2_fill_1 FILLER_69_809 ();
 sg13g2_fill_1 FILLER_69_832 ();
 sg13g2_fill_1 FILLER_69_869 ();
 sg13g2_fill_1 FILLER_69_884 ();
 sg13g2_fill_1 FILLER_69_894 ();
 sg13g2_fill_1 FILLER_69_937 ();
 sg13g2_fill_2 FILLER_69_951 ();
 sg13g2_fill_1 FILLER_69_953 ();
 sg13g2_fill_2 FILLER_69_959 ();
 sg13g2_fill_2 FILLER_69_965 ();
 sg13g2_decap_4 FILLER_69_971 ();
 sg13g2_fill_2 FILLER_69_998 ();
 sg13g2_fill_2 FILLER_69_1003 ();
 sg13g2_fill_1 FILLER_69_1005 ();
 sg13g2_decap_4 FILLER_69_1010 ();
 sg13g2_fill_2 FILLER_69_1053 ();
 sg13g2_fill_1 FILLER_69_1080 ();
 sg13g2_fill_1 FILLER_69_1088 ();
 sg13g2_fill_1 FILLER_69_1161 ();
 sg13g2_decap_8 FILLER_69_1178 ();
 sg13g2_decap_4 FILLER_69_1185 ();
 sg13g2_decap_8 FILLER_69_1193 ();
 sg13g2_decap_4 FILLER_69_1200 ();
 sg13g2_fill_2 FILLER_69_1204 ();
 sg13g2_fill_2 FILLER_69_1216 ();
 sg13g2_decap_4 FILLER_69_1229 ();
 sg13g2_fill_1 FILLER_69_1233 ();
 sg13g2_fill_2 FILLER_69_1264 ();
 sg13g2_decap_4 FILLER_69_1284 ();
 sg13g2_fill_2 FILLER_69_1328 ();
 sg13g2_fill_2 FILLER_69_1349 ();
 sg13g2_fill_2 FILLER_69_1368 ();
 sg13g2_fill_1 FILLER_69_1370 ();
 sg13g2_decap_8 FILLER_69_1384 ();
 sg13g2_decap_4 FILLER_69_1391 ();
 sg13g2_fill_1 FILLER_69_1395 ();
 sg13g2_fill_2 FILLER_69_1417 ();
 sg13g2_fill_1 FILLER_69_1419 ();
 sg13g2_fill_1 FILLER_69_1459 ();
 sg13g2_fill_1 FILLER_69_1465 ();
 sg13g2_fill_2 FILLER_69_1479 ();
 sg13g2_fill_2 FILLER_69_1524 ();
 sg13g2_fill_1 FILLER_69_1526 ();
 sg13g2_fill_2 FILLER_69_1557 ();
 sg13g2_fill_1 FILLER_69_1572 ();
 sg13g2_fill_2 FILLER_69_1599 ();
 sg13g2_decap_4 FILLER_69_1701 ();
 sg13g2_fill_1 FILLER_69_1705 ();
 sg13g2_fill_2 FILLER_69_1732 ();
 sg13g2_fill_2 FILLER_69_1751 ();
 sg13g2_fill_2 FILLER_69_1788 ();
 sg13g2_fill_1 FILLER_69_1790 ();
 sg13g2_decap_8 FILLER_69_1795 ();
 sg13g2_decap_8 FILLER_69_1802 ();
 sg13g2_fill_2 FILLER_69_1809 ();
 sg13g2_fill_1 FILLER_69_1811 ();
 sg13g2_decap_4 FILLER_69_1821 ();
 sg13g2_decap_4 FILLER_69_1834 ();
 sg13g2_fill_1 FILLER_69_1838 ();
 sg13g2_decap_4 FILLER_69_1842 ();
 sg13g2_fill_1 FILLER_69_1846 ();
 sg13g2_fill_2 FILLER_69_1878 ();
 sg13g2_fill_1 FILLER_69_1880 ();
 sg13g2_fill_1 FILLER_69_1907 ();
 sg13g2_decap_8 FILLER_69_1934 ();
 sg13g2_fill_1 FILLER_69_1946 ();
 sg13g2_decap_8 FILLER_69_1957 ();
 sg13g2_decap_8 FILLER_69_1964 ();
 sg13g2_fill_2 FILLER_69_1971 ();
 sg13g2_fill_2 FILLER_69_1999 ();
 sg13g2_fill_2 FILLER_69_2053 ();
 sg13g2_decap_4 FILLER_69_2081 ();
 sg13g2_fill_1 FILLER_69_2090 ();
 sg13g2_decap_8 FILLER_69_2107 ();
 sg13g2_fill_2 FILLER_69_2114 ();
 sg13g2_decap_4 FILLER_69_2126 ();
 sg13g2_fill_2 FILLER_69_2130 ();
 sg13g2_fill_2 FILLER_69_2145 ();
 sg13g2_decap_8 FILLER_69_2164 ();
 sg13g2_decap_8 FILLER_69_2171 ();
 sg13g2_decap_4 FILLER_69_2187 ();
 sg13g2_fill_2 FILLER_69_2191 ();
 sg13g2_fill_2 FILLER_69_2197 ();
 sg13g2_decap_4 FILLER_69_2230 ();
 sg13g2_decap_4 FILLER_69_2238 ();
 sg13g2_fill_1 FILLER_69_2242 ();
 sg13g2_decap_8 FILLER_69_2249 ();
 sg13g2_decap_4 FILLER_69_2260 ();
 sg13g2_fill_2 FILLER_69_2272 ();
 sg13g2_fill_1 FILLER_69_2274 ();
 sg13g2_decap_8 FILLER_69_2285 ();
 sg13g2_fill_2 FILLER_69_2309 ();
 sg13g2_fill_1 FILLER_69_2311 ();
 sg13g2_fill_1 FILLER_69_2325 ();
 sg13g2_fill_2 FILLER_69_2397 ();
 sg13g2_decap_4 FILLER_69_2410 ();
 sg13g2_fill_2 FILLER_69_2414 ();
 sg13g2_fill_2 FILLER_69_2429 ();
 sg13g2_fill_1 FILLER_69_2444 ();
 sg13g2_decap_8 FILLER_69_2470 ();
 sg13g2_fill_1 FILLER_69_2477 ();
 sg13g2_fill_1 FILLER_69_2504 ();
 sg13g2_decap_8 FILLER_69_2537 ();
 sg13g2_fill_2 FILLER_69_2544 ();
 sg13g2_decap_8 FILLER_69_2550 ();
 sg13g2_fill_1 FILLER_69_2557 ();
 sg13g2_fill_1 FILLER_69_2567 ();
 sg13g2_fill_1 FILLER_69_2574 ();
 sg13g2_fill_1 FILLER_69_2584 ();
 sg13g2_decap_8 FILLER_69_2610 ();
 sg13g2_fill_2 FILLER_69_2617 ();
 sg13g2_fill_1 FILLER_69_2619 ();
 sg13g2_decap_8 FILLER_69_2633 ();
 sg13g2_fill_2 FILLER_69_2640 ();
 sg13g2_fill_1 FILLER_69_2642 ();
 sg13g2_fill_1 FILLER_69_2691 ();
 sg13g2_fill_1 FILLER_69_2700 ();
 sg13g2_fill_2 FILLER_69_2711 ();
 sg13g2_fill_1 FILLER_69_2744 ();
 sg13g2_fill_2 FILLER_69_2758 ();
 sg13g2_fill_1 FILLER_69_2760 ();
 sg13g2_fill_2 FILLER_69_2787 ();
 sg13g2_fill_2 FILLER_69_2811 ();
 sg13g2_fill_1 FILLER_69_2823 ();
 sg13g2_fill_2 FILLER_69_2843 ();
 sg13g2_decap_4 FILLER_69_2882 ();
 sg13g2_fill_2 FILLER_69_2910 ();
 sg13g2_fill_1 FILLER_69_2912 ();
 sg13g2_fill_1 FILLER_69_2928 ();
 sg13g2_decap_8 FILLER_69_2981 ();
 sg13g2_decap_8 FILLER_69_2988 ();
 sg13g2_decap_8 FILLER_69_2995 ();
 sg13g2_decap_8 FILLER_69_3002 ();
 sg13g2_decap_8 FILLER_69_3009 ();
 sg13g2_decap_8 FILLER_69_3016 ();
 sg13g2_decap_8 FILLER_69_3023 ();
 sg13g2_decap_8 FILLER_69_3030 ();
 sg13g2_decap_8 FILLER_69_3037 ();
 sg13g2_decap_8 FILLER_69_3044 ();
 sg13g2_decap_8 FILLER_69_3051 ();
 sg13g2_decap_8 FILLER_69_3058 ();
 sg13g2_decap_8 FILLER_69_3065 ();
 sg13g2_decap_8 FILLER_69_3072 ();
 sg13g2_decap_8 FILLER_69_3079 ();
 sg13g2_decap_8 FILLER_69_3086 ();
 sg13g2_decap_8 FILLER_69_3093 ();
 sg13g2_decap_8 FILLER_69_3100 ();
 sg13g2_decap_8 FILLER_69_3107 ();
 sg13g2_decap_8 FILLER_69_3114 ();
 sg13g2_decap_8 FILLER_69_3121 ();
 sg13g2_decap_8 FILLER_69_3128 ();
 sg13g2_decap_8 FILLER_69_3135 ();
 sg13g2_decap_8 FILLER_69_3142 ();
 sg13g2_decap_8 FILLER_69_3149 ();
 sg13g2_decap_8 FILLER_69_3156 ();
 sg13g2_decap_8 FILLER_69_3163 ();
 sg13g2_decap_8 FILLER_69_3170 ();
 sg13g2_decap_8 FILLER_69_3177 ();
 sg13g2_decap_8 FILLER_69_3184 ();
 sg13g2_decap_8 FILLER_69_3191 ();
 sg13g2_decap_8 FILLER_69_3198 ();
 sg13g2_decap_8 FILLER_69_3205 ();
 sg13g2_decap_8 FILLER_69_3212 ();
 sg13g2_decap_8 FILLER_69_3219 ();
 sg13g2_decap_8 FILLER_69_3226 ();
 sg13g2_decap_8 FILLER_69_3233 ();
 sg13g2_decap_8 FILLER_69_3240 ();
 sg13g2_decap_8 FILLER_69_3247 ();
 sg13g2_decap_8 FILLER_69_3254 ();
 sg13g2_decap_8 FILLER_69_3261 ();
 sg13g2_decap_8 FILLER_69_3268 ();
 sg13g2_decap_8 FILLER_69_3275 ();
 sg13g2_decap_8 FILLER_69_3282 ();
 sg13g2_decap_8 FILLER_69_3289 ();
 sg13g2_decap_8 FILLER_69_3296 ();
 sg13g2_decap_8 FILLER_69_3303 ();
 sg13g2_decap_8 FILLER_69_3310 ();
 sg13g2_decap_8 FILLER_69_3317 ();
 sg13g2_decap_8 FILLER_69_3324 ();
 sg13g2_decap_8 FILLER_69_3331 ();
 sg13g2_decap_8 FILLER_69_3338 ();
 sg13g2_decap_8 FILLER_69_3345 ();
 sg13g2_decap_8 FILLER_69_3352 ();
 sg13g2_decap_8 FILLER_69_3359 ();
 sg13g2_decap_8 FILLER_69_3366 ();
 sg13g2_decap_8 FILLER_69_3373 ();
 sg13g2_decap_8 FILLER_69_3380 ();
 sg13g2_decap_8 FILLER_69_3387 ();
 sg13g2_decap_8 FILLER_69_3394 ();
 sg13g2_decap_8 FILLER_69_3401 ();
 sg13g2_decap_8 FILLER_69_3408 ();
 sg13g2_decap_8 FILLER_69_3415 ();
 sg13g2_decap_8 FILLER_69_3422 ();
 sg13g2_decap_8 FILLER_69_3429 ();
 sg13g2_decap_8 FILLER_69_3436 ();
 sg13g2_decap_8 FILLER_69_3443 ();
 sg13g2_decap_8 FILLER_69_3450 ();
 sg13g2_decap_8 FILLER_69_3457 ();
 sg13g2_decap_8 FILLER_69_3464 ();
 sg13g2_decap_8 FILLER_69_3471 ();
 sg13g2_decap_8 FILLER_69_3478 ();
 sg13g2_decap_8 FILLER_69_3485 ();
 sg13g2_decap_8 FILLER_69_3492 ();
 sg13g2_decap_8 FILLER_69_3499 ();
 sg13g2_decap_8 FILLER_69_3506 ();
 sg13g2_decap_8 FILLER_69_3513 ();
 sg13g2_decap_8 FILLER_69_3520 ();
 sg13g2_decap_8 FILLER_69_3527 ();
 sg13g2_decap_8 FILLER_69_3534 ();
 sg13g2_decap_8 FILLER_69_3541 ();
 sg13g2_decap_8 FILLER_69_3548 ();
 sg13g2_decap_8 FILLER_69_3555 ();
 sg13g2_decap_8 FILLER_69_3562 ();
 sg13g2_decap_8 FILLER_69_3569 ();
 sg13g2_decap_4 FILLER_69_3576 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_fill_2 FILLER_70_28 ();
 sg13g2_fill_1 FILLER_70_30 ();
 sg13g2_decap_8 FILLER_70_40 ();
 sg13g2_decap_4 FILLER_70_47 ();
 sg13g2_fill_1 FILLER_70_51 ();
 sg13g2_decap_4 FILLER_70_56 ();
 sg13g2_fill_1 FILLER_70_60 ();
 sg13g2_fill_1 FILLER_70_87 ();
 sg13g2_fill_2 FILLER_70_114 ();
 sg13g2_fill_1 FILLER_70_116 ();
 sg13g2_fill_1 FILLER_70_122 ();
 sg13g2_decap_4 FILLER_70_135 ();
 sg13g2_fill_1 FILLER_70_143 ();
 sg13g2_decap_8 FILLER_70_179 ();
 sg13g2_decap_4 FILLER_70_186 ();
 sg13g2_fill_2 FILLER_70_190 ();
 sg13g2_decap_4 FILLER_70_196 ();
 sg13g2_fill_2 FILLER_70_257 ();
 sg13g2_decap_4 FILLER_70_275 ();
 sg13g2_fill_2 FILLER_70_279 ();
 sg13g2_fill_1 FILLER_70_291 ();
 sg13g2_decap_8 FILLER_70_344 ();
 sg13g2_fill_2 FILLER_70_351 ();
 sg13g2_fill_1 FILLER_70_358 ();
 sg13g2_fill_2 FILLER_70_388 ();
 sg13g2_fill_2 FILLER_70_400 ();
 sg13g2_fill_1 FILLER_70_406 ();
 sg13g2_fill_2 FILLER_70_429 ();
 sg13g2_decap_4 FILLER_70_457 ();
 sg13g2_fill_2 FILLER_70_504 ();
 sg13g2_fill_1 FILLER_70_541 ();
 sg13g2_fill_1 FILLER_70_551 ();
 sg13g2_decap_4 FILLER_70_582 ();
 sg13g2_fill_1 FILLER_70_586 ();
 sg13g2_fill_2 FILLER_70_631 ();
 sg13g2_fill_1 FILLER_70_633 ();
 sg13g2_fill_1 FILLER_70_664 ();
 sg13g2_fill_1 FILLER_70_670 ();
 sg13g2_decap_8 FILLER_70_698 ();
 sg13g2_decap_4 FILLER_70_705 ();
 sg13g2_decap_8 FILLER_70_718 ();
 sg13g2_decap_8 FILLER_70_725 ();
 sg13g2_fill_1 FILLER_70_732 ();
 sg13g2_decap_4 FILLER_70_738 ();
 sg13g2_fill_1 FILLER_70_742 ();
 sg13g2_decap_4 FILLER_70_746 ();
 sg13g2_fill_2 FILLER_70_750 ();
 sg13g2_decap_8 FILLER_70_769 ();
 sg13g2_fill_2 FILLER_70_776 ();
 sg13g2_fill_1 FILLER_70_778 ();
 sg13g2_fill_1 FILLER_70_793 ();
 sg13g2_decap_8 FILLER_70_815 ();
 sg13g2_decap_4 FILLER_70_822 ();
 sg13g2_fill_1 FILLER_70_826 ();
 sg13g2_decap_4 FILLER_70_853 ();
 sg13g2_fill_2 FILLER_70_857 ();
 sg13g2_fill_2 FILLER_70_924 ();
 sg13g2_fill_1 FILLER_70_926 ();
 sg13g2_fill_2 FILLER_70_953 ();
 sg13g2_fill_1 FILLER_70_955 ();
 sg13g2_decap_8 FILLER_70_971 ();
 sg13g2_decap_4 FILLER_70_978 ();
 sg13g2_decap_8 FILLER_70_1058 ();
 sg13g2_fill_2 FILLER_70_1071 ();
 sg13g2_decap_8 FILLER_70_1082 ();
 sg13g2_fill_1 FILLER_70_1112 ();
 sg13g2_fill_2 FILLER_70_1122 ();
 sg13g2_fill_2 FILLER_70_1133 ();
 sg13g2_fill_1 FILLER_70_1135 ();
 sg13g2_fill_2 FILLER_70_1145 ();
 sg13g2_fill_1 FILLER_70_1147 ();
 sg13g2_decap_8 FILLER_70_1170 ();
 sg13g2_decap_4 FILLER_70_1177 ();
 sg13g2_fill_1 FILLER_70_1181 ();
 sg13g2_fill_1 FILLER_70_1187 ();
 sg13g2_decap_8 FILLER_70_1198 ();
 sg13g2_fill_1 FILLER_70_1235 ();
 sg13g2_fill_2 FILLER_70_1241 ();
 sg13g2_fill_1 FILLER_70_1252 ();
 sg13g2_fill_1 FILLER_70_1279 ();
 sg13g2_decap_8 FILLER_70_1285 ();
 sg13g2_fill_2 FILLER_70_1292 ();
 sg13g2_decap_8 FILLER_70_1303 ();
 sg13g2_decap_4 FILLER_70_1310 ();
 sg13g2_fill_1 FILLER_70_1314 ();
 sg13g2_fill_2 FILLER_70_1341 ();
 sg13g2_fill_1 FILLER_70_1343 ();
 sg13g2_fill_2 FILLER_70_1383 ();
 sg13g2_fill_2 FILLER_70_1416 ();
 sg13g2_fill_1 FILLER_70_1467 ();
 sg13g2_fill_2 FILLER_70_1481 ();
 sg13g2_fill_1 FILLER_70_1483 ();
 sg13g2_decap_4 FILLER_70_1519 ();
 sg13g2_fill_2 FILLER_70_1592 ();
 sg13g2_fill_1 FILLER_70_1668 ();
 sg13g2_fill_1 FILLER_70_1678 ();
 sg13g2_decap_8 FILLER_70_1692 ();
 sg13g2_decap_8 FILLER_70_1699 ();
 sg13g2_decap_8 FILLER_70_1706 ();
 sg13g2_decap_4 FILLER_70_1721 ();
 sg13g2_decap_4 FILLER_70_1764 ();
 sg13g2_fill_1 FILLER_70_1768 ();
 sg13g2_fill_1 FILLER_70_1773 ();
 sg13g2_decap_8 FILLER_70_1778 ();
 sg13g2_fill_1 FILLER_70_1814 ();
 sg13g2_decap_4 FILLER_70_1847 ();
 sg13g2_fill_2 FILLER_70_1851 ();
 sg13g2_decap_8 FILLER_70_1879 ();
 sg13g2_decap_8 FILLER_70_1886 ();
 sg13g2_decap_4 FILLER_70_1902 ();
 sg13g2_decap_8 FILLER_70_1929 ();
 sg13g2_fill_1 FILLER_70_1936 ();
 sg13g2_fill_2 FILLER_70_1942 ();
 sg13g2_fill_1 FILLER_70_1944 ();
 sg13g2_fill_1 FILLER_70_1955 ();
 sg13g2_decap_4 FILLER_70_1985 ();
 sg13g2_fill_1 FILLER_70_2012 ();
 sg13g2_decap_8 FILLER_70_2018 ();
 sg13g2_decap_8 FILLER_70_2025 ();
 sg13g2_decap_4 FILLER_70_2032 ();
 sg13g2_fill_2 FILLER_70_2036 ();
 sg13g2_decap_8 FILLER_70_2042 ();
 sg13g2_fill_1 FILLER_70_2049 ();
 sg13g2_decap_8 FILLER_70_2055 ();
 sg13g2_decap_4 FILLER_70_2062 ();
 sg13g2_fill_2 FILLER_70_2070 ();
 sg13g2_fill_1 FILLER_70_2077 ();
 sg13g2_decap_8 FILLER_70_2082 ();
 sg13g2_fill_1 FILLER_70_2094 ();
 sg13g2_decap_8 FILLER_70_2108 ();
 sg13g2_fill_2 FILLER_70_2115 ();
 sg13g2_fill_1 FILLER_70_2117 ();
 sg13g2_fill_2 FILLER_70_2144 ();
 sg13g2_fill_1 FILLER_70_2146 ();
 sg13g2_fill_2 FILLER_70_2177 ();
 sg13g2_fill_1 FILLER_70_2179 ();
 sg13g2_decap_8 FILLER_70_2188 ();
 sg13g2_fill_1 FILLER_70_2195 ();
 sg13g2_fill_1 FILLER_70_2217 ();
 sg13g2_fill_1 FILLER_70_2232 ();
 sg13g2_fill_1 FILLER_70_2241 ();
 sg13g2_fill_2 FILLER_70_2259 ();
 sg13g2_decap_8 FILLER_70_2265 ();
 sg13g2_fill_1 FILLER_70_2272 ();
 sg13g2_decap_4 FILLER_70_2285 ();
 sg13g2_fill_1 FILLER_70_2289 ();
 sg13g2_fill_2 FILLER_70_2294 ();
 sg13g2_decap_8 FILLER_70_2319 ();
 sg13g2_fill_2 FILLER_70_2341 ();
 sg13g2_fill_1 FILLER_70_2352 ();
 sg13g2_decap_8 FILLER_70_2375 ();
 sg13g2_fill_2 FILLER_70_2390 ();
 sg13g2_fill_2 FILLER_70_2400 ();
 sg13g2_fill_1 FILLER_70_2402 ();
 sg13g2_fill_2 FILLER_70_2411 ();
 sg13g2_decap_4 FILLER_70_2439 ();
 sg13g2_fill_2 FILLER_70_2454 ();
 sg13g2_decap_8 FILLER_70_2470 ();
 sg13g2_decap_4 FILLER_70_2477 ();
 sg13g2_fill_1 FILLER_70_2481 ();
 sg13g2_fill_2 FILLER_70_2487 ();
 sg13g2_decap_8 FILLER_70_2493 ();
 sg13g2_decap_8 FILLER_70_2500 ();
 sg13g2_fill_1 FILLER_70_2512 ();
 sg13g2_decap_4 FILLER_70_2517 ();
 sg13g2_fill_1 FILLER_70_2521 ();
 sg13g2_decap_4 FILLER_70_2526 ();
 sg13g2_fill_2 FILLER_70_2530 ();
 sg13g2_fill_1 FILLER_70_2588 ();
 sg13g2_decap_4 FILLER_70_2598 ();
 sg13g2_fill_1 FILLER_70_2602 ();
 sg13g2_decap_4 FILLER_70_2629 ();
 sg13g2_fill_2 FILLER_70_2633 ();
 sg13g2_decap_4 FILLER_70_2639 ();
 sg13g2_fill_2 FILLER_70_2650 ();
 sg13g2_fill_1 FILLER_70_2652 ();
 sg13g2_fill_2 FILLER_70_2666 ();
 sg13g2_fill_1 FILLER_70_2668 ();
 sg13g2_decap_8 FILLER_70_2685 ();
 sg13g2_fill_1 FILLER_70_2692 ();
 sg13g2_decap_8 FILLER_70_2708 ();
 sg13g2_decap_8 FILLER_70_2715 ();
 sg13g2_fill_2 FILLER_70_2735 ();
 sg13g2_decap_8 FILLER_70_2752 ();
 sg13g2_decap_8 FILLER_70_2759 ();
 sg13g2_decap_8 FILLER_70_2766 ();
 sg13g2_fill_1 FILLER_70_2782 ();
 sg13g2_fill_2 FILLER_70_2788 ();
 sg13g2_decap_4 FILLER_70_2798 ();
 sg13g2_fill_1 FILLER_70_2820 ();
 sg13g2_decap_8 FILLER_70_2847 ();
 sg13g2_fill_2 FILLER_70_2854 ();
 sg13g2_fill_1 FILLER_70_2856 ();
 sg13g2_decap_4 FILLER_70_2861 ();
 sg13g2_fill_1 FILLER_70_2865 ();
 sg13g2_decap_4 FILLER_70_2879 ();
 sg13g2_decap_8 FILLER_70_2896 ();
 sg13g2_decap_4 FILLER_70_2903 ();
 sg13g2_fill_2 FILLER_70_2914 ();
 sg13g2_fill_1 FILLER_70_2938 ();
 sg13g2_decap_8 FILLER_70_2966 ();
 sg13g2_decap_8 FILLER_70_2973 ();
 sg13g2_decap_8 FILLER_70_2980 ();
 sg13g2_decap_8 FILLER_70_2987 ();
 sg13g2_decap_8 FILLER_70_2994 ();
 sg13g2_decap_8 FILLER_70_3001 ();
 sg13g2_decap_8 FILLER_70_3008 ();
 sg13g2_decap_8 FILLER_70_3015 ();
 sg13g2_decap_8 FILLER_70_3022 ();
 sg13g2_decap_8 FILLER_70_3029 ();
 sg13g2_decap_8 FILLER_70_3036 ();
 sg13g2_decap_8 FILLER_70_3043 ();
 sg13g2_decap_8 FILLER_70_3050 ();
 sg13g2_decap_8 FILLER_70_3057 ();
 sg13g2_decap_8 FILLER_70_3064 ();
 sg13g2_decap_8 FILLER_70_3071 ();
 sg13g2_decap_8 FILLER_70_3078 ();
 sg13g2_decap_8 FILLER_70_3085 ();
 sg13g2_decap_8 FILLER_70_3092 ();
 sg13g2_decap_8 FILLER_70_3099 ();
 sg13g2_decap_8 FILLER_70_3106 ();
 sg13g2_decap_8 FILLER_70_3113 ();
 sg13g2_decap_8 FILLER_70_3120 ();
 sg13g2_decap_8 FILLER_70_3127 ();
 sg13g2_decap_8 FILLER_70_3134 ();
 sg13g2_decap_8 FILLER_70_3141 ();
 sg13g2_decap_8 FILLER_70_3148 ();
 sg13g2_decap_8 FILLER_70_3155 ();
 sg13g2_decap_8 FILLER_70_3162 ();
 sg13g2_decap_8 FILLER_70_3169 ();
 sg13g2_decap_8 FILLER_70_3176 ();
 sg13g2_decap_8 FILLER_70_3183 ();
 sg13g2_decap_8 FILLER_70_3190 ();
 sg13g2_decap_8 FILLER_70_3197 ();
 sg13g2_decap_8 FILLER_70_3204 ();
 sg13g2_decap_8 FILLER_70_3211 ();
 sg13g2_decap_8 FILLER_70_3218 ();
 sg13g2_decap_8 FILLER_70_3225 ();
 sg13g2_decap_8 FILLER_70_3232 ();
 sg13g2_decap_8 FILLER_70_3239 ();
 sg13g2_decap_8 FILLER_70_3246 ();
 sg13g2_decap_8 FILLER_70_3253 ();
 sg13g2_decap_8 FILLER_70_3260 ();
 sg13g2_decap_8 FILLER_70_3267 ();
 sg13g2_decap_8 FILLER_70_3274 ();
 sg13g2_decap_8 FILLER_70_3281 ();
 sg13g2_decap_8 FILLER_70_3288 ();
 sg13g2_decap_8 FILLER_70_3295 ();
 sg13g2_decap_8 FILLER_70_3302 ();
 sg13g2_decap_8 FILLER_70_3309 ();
 sg13g2_decap_8 FILLER_70_3316 ();
 sg13g2_decap_8 FILLER_70_3323 ();
 sg13g2_decap_8 FILLER_70_3330 ();
 sg13g2_decap_8 FILLER_70_3337 ();
 sg13g2_decap_8 FILLER_70_3344 ();
 sg13g2_decap_8 FILLER_70_3351 ();
 sg13g2_decap_8 FILLER_70_3358 ();
 sg13g2_decap_8 FILLER_70_3365 ();
 sg13g2_decap_8 FILLER_70_3372 ();
 sg13g2_decap_8 FILLER_70_3379 ();
 sg13g2_decap_8 FILLER_70_3386 ();
 sg13g2_decap_8 FILLER_70_3393 ();
 sg13g2_decap_8 FILLER_70_3400 ();
 sg13g2_decap_8 FILLER_70_3407 ();
 sg13g2_decap_8 FILLER_70_3414 ();
 sg13g2_decap_8 FILLER_70_3421 ();
 sg13g2_decap_8 FILLER_70_3428 ();
 sg13g2_decap_8 FILLER_70_3435 ();
 sg13g2_decap_8 FILLER_70_3442 ();
 sg13g2_decap_8 FILLER_70_3449 ();
 sg13g2_decap_8 FILLER_70_3456 ();
 sg13g2_decap_8 FILLER_70_3463 ();
 sg13g2_decap_8 FILLER_70_3470 ();
 sg13g2_decap_8 FILLER_70_3477 ();
 sg13g2_decap_8 FILLER_70_3484 ();
 sg13g2_decap_8 FILLER_70_3491 ();
 sg13g2_decap_8 FILLER_70_3498 ();
 sg13g2_decap_8 FILLER_70_3505 ();
 sg13g2_decap_8 FILLER_70_3512 ();
 sg13g2_decap_8 FILLER_70_3519 ();
 sg13g2_decap_8 FILLER_70_3526 ();
 sg13g2_decap_8 FILLER_70_3533 ();
 sg13g2_decap_8 FILLER_70_3540 ();
 sg13g2_decap_8 FILLER_70_3547 ();
 sg13g2_decap_8 FILLER_70_3554 ();
 sg13g2_decap_8 FILLER_70_3561 ();
 sg13g2_decap_8 FILLER_70_3568 ();
 sg13g2_decap_4 FILLER_70_3575 ();
 sg13g2_fill_1 FILLER_70_3579 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_fill_2 FILLER_71_28 ();
 sg13g2_fill_2 FILLER_71_56 ();
 sg13g2_fill_1 FILLER_71_58 ();
 sg13g2_decap_8 FILLER_71_64 ();
 sg13g2_decap_8 FILLER_71_71 ();
 sg13g2_fill_2 FILLER_71_103 ();
 sg13g2_fill_1 FILLER_71_166 ();
 sg13g2_decap_4 FILLER_71_212 ();
 sg13g2_fill_1 FILLER_71_216 ();
 sg13g2_fill_2 FILLER_71_243 ();
 sg13g2_decap_8 FILLER_71_264 ();
 sg13g2_fill_2 FILLER_71_297 ();
 sg13g2_fill_1 FILLER_71_299 ();
 sg13g2_fill_2 FILLER_71_326 ();
 sg13g2_fill_1 FILLER_71_328 ();
 sg13g2_decap_4 FILLER_71_355 ();
 sg13g2_fill_2 FILLER_71_384 ();
 sg13g2_fill_1 FILLER_71_386 ();
 sg13g2_fill_2 FILLER_71_393 ();
 sg13g2_decap_8 FILLER_71_400 ();
 sg13g2_decap_4 FILLER_71_407 ();
 sg13g2_fill_2 FILLER_71_417 ();
 sg13g2_fill_1 FILLER_71_419 ();
 sg13g2_fill_1 FILLER_71_425 ();
 sg13g2_fill_2 FILLER_71_431 ();
 sg13g2_fill_1 FILLER_71_433 ();
 sg13g2_fill_2 FILLER_71_439 ();
 sg13g2_fill_1 FILLER_71_441 ();
 sg13g2_fill_2 FILLER_71_477 ();
 sg13g2_fill_2 FILLER_71_488 ();
 sg13g2_fill_1 FILLER_71_490 ();
 sg13g2_fill_2 FILLER_71_526 ();
 sg13g2_fill_2 FILLER_71_554 ();
 sg13g2_fill_2 FILLER_71_592 ();
 sg13g2_fill_1 FILLER_71_594 ();
 sg13g2_fill_2 FILLER_71_600 ();
 sg13g2_fill_1 FILLER_71_602 ();
 sg13g2_decap_8 FILLER_71_640 ();
 sg13g2_fill_1 FILLER_71_690 ();
 sg13g2_decap_8 FILLER_71_722 ();
 sg13g2_decap_8 FILLER_71_729 ();
 sg13g2_fill_2 FILLER_71_805 ();
 sg13g2_fill_1 FILLER_71_807 ();
 sg13g2_fill_1 FILLER_71_812 ();
 sg13g2_decap_4 FILLER_71_826 ();
 sg13g2_fill_1 FILLER_71_830 ();
 sg13g2_fill_2 FILLER_71_835 ();
 sg13g2_fill_1 FILLER_71_837 ();
 sg13g2_fill_1 FILLER_71_842 ();
 sg13g2_decap_8 FILLER_71_846 ();
 sg13g2_decap_8 FILLER_71_853 ();
 sg13g2_decap_8 FILLER_71_860 ();
 sg13g2_fill_2 FILLER_71_867 ();
 sg13g2_decap_4 FILLER_71_881 ();
 sg13g2_decap_4 FILLER_71_922 ();
 sg13g2_decap_4 FILLER_71_932 ();
 sg13g2_fill_1 FILLER_71_946 ();
 sg13g2_fill_1 FILLER_71_952 ();
 sg13g2_decap_8 FILLER_71_985 ();
 sg13g2_fill_1 FILLER_71_992 ();
 sg13g2_decap_4 FILLER_71_997 ();
 sg13g2_fill_2 FILLER_71_1001 ();
 sg13g2_decap_8 FILLER_71_1013 ();
 sg13g2_decap_4 FILLER_71_1020 ();
 sg13g2_fill_1 FILLER_71_1024 ();
 sg13g2_fill_2 FILLER_71_1049 ();
 sg13g2_fill_1 FILLER_71_1083 ();
 sg13g2_fill_1 FILLER_71_1119 ();
 sg13g2_decap_4 FILLER_71_1177 ();
 sg13g2_fill_2 FILLER_71_1216 ();
 sg13g2_fill_2 FILLER_71_1244 ();
 sg13g2_fill_1 FILLER_71_1246 ();
 sg13g2_fill_2 FILLER_71_1252 ();
 sg13g2_fill_1 FILLER_71_1259 ();
 sg13g2_fill_1 FILLER_71_1266 ();
 sg13g2_decap_4 FILLER_71_1276 ();
 sg13g2_decap_8 FILLER_71_1317 ();
 sg13g2_fill_1 FILLER_71_1324 ();
 sg13g2_decap_8 FILLER_71_1329 ();
 sg13g2_decap_4 FILLER_71_1336 ();
 sg13g2_fill_1 FILLER_71_1340 ();
 sg13g2_decap_4 FILLER_71_1345 ();
 sg13g2_fill_2 FILLER_71_1349 ();
 sg13g2_fill_1 FILLER_71_1356 ();
 sg13g2_decap_8 FILLER_71_1385 ();
 sg13g2_fill_1 FILLER_71_1392 ();
 sg13g2_fill_2 FILLER_71_1397 ();
 sg13g2_fill_1 FILLER_71_1399 ();
 sg13g2_fill_2 FILLER_71_1409 ();
 sg13g2_fill_1 FILLER_71_1416 ();
 sg13g2_fill_2 FILLER_71_1427 ();
 sg13g2_fill_1 FILLER_71_1433 ();
 sg13g2_decap_8 FILLER_71_1460 ();
 sg13g2_decap_4 FILLER_71_1467 ();
 sg13g2_fill_1 FILLER_71_1480 ();
 sg13g2_fill_2 FILLER_71_1485 ();
 sg13g2_fill_2 FILLER_71_1496 ();
 sg13g2_fill_1 FILLER_71_1518 ();
 sg13g2_fill_1 FILLER_71_1534 ();
 sg13g2_decap_4 FILLER_71_1554 ();
 sg13g2_fill_1 FILLER_71_1558 ();
 sg13g2_fill_1 FILLER_71_1566 ();
 sg13g2_fill_1 FILLER_71_1590 ();
 sg13g2_fill_1 FILLER_71_1617 ();
 sg13g2_fill_1 FILLER_71_1633 ();
 sg13g2_fill_2 FILLER_71_1690 ();
 sg13g2_fill_2 FILLER_71_1696 ();
 sg13g2_fill_1 FILLER_71_1698 ();
 sg13g2_decap_4 FILLER_71_1712 ();
 sg13g2_fill_1 FILLER_71_1716 ();
 sg13g2_fill_1 FILLER_71_1721 ();
 sg13g2_decap_8 FILLER_71_1728 ();
 sg13g2_decap_8 FILLER_71_1743 ();
 sg13g2_decap_8 FILLER_71_1754 ();
 sg13g2_fill_2 FILLER_71_1761 ();
 sg13g2_decap_8 FILLER_71_1824 ();
 sg13g2_fill_1 FILLER_71_1831 ();
 sg13g2_decap_8 FILLER_71_1836 ();
 sg13g2_fill_1 FILLER_71_1843 ();
 sg13g2_fill_1 FILLER_71_1853 ();
 sg13g2_fill_2 FILLER_71_1858 ();
 sg13g2_decap_8 FILLER_71_1873 ();
 sg13g2_decap_4 FILLER_71_1880 ();
 sg13g2_fill_1 FILLER_71_1884 ();
 sg13g2_fill_2 FILLER_71_1909 ();
 sg13g2_fill_1 FILLER_71_1911 ();
 sg13g2_fill_2 FILLER_71_1940 ();
 sg13g2_decap_4 FILLER_71_1952 ();
 sg13g2_fill_1 FILLER_71_1956 ();
 sg13g2_fill_2 FILLER_71_1993 ();
 sg13g2_decap_8 FILLER_71_2025 ();
 sg13g2_decap_8 FILLER_71_2032 ();
 sg13g2_fill_2 FILLER_71_2039 ();
 sg13g2_fill_2 FILLER_71_2045 ();
 sg13g2_fill_1 FILLER_71_2047 ();
 sg13g2_fill_1 FILLER_71_2056 ();
 sg13g2_fill_1 FILLER_71_2093 ();
 sg13g2_fill_1 FILLER_71_2099 ();
 sg13g2_fill_2 FILLER_71_2117 ();
 sg13g2_fill_2 FILLER_71_2124 ();
 sg13g2_fill_1 FILLER_71_2126 ();
 sg13g2_fill_2 FILLER_71_2141 ();
 sg13g2_fill_1 FILLER_71_2143 ();
 sg13g2_fill_1 FILLER_71_2149 ();
 sg13g2_decap_8 FILLER_71_2166 ();
 sg13g2_fill_1 FILLER_71_2188 ();
 sg13g2_fill_2 FILLER_71_2213 ();
 sg13g2_decap_4 FILLER_71_2219 ();
 sg13g2_fill_2 FILLER_71_2243 ();
 sg13g2_fill_1 FILLER_71_2245 ();
 sg13g2_fill_2 FILLER_71_2251 ();
 sg13g2_fill_1 FILLER_71_2277 ();
 sg13g2_decap_4 FILLER_71_2304 ();
 sg13g2_fill_2 FILLER_71_2317 ();
 sg13g2_fill_2 FILLER_71_2338 ();
 sg13g2_fill_1 FILLER_71_2340 ();
 sg13g2_fill_1 FILLER_71_2354 ();
 sg13g2_decap_4 FILLER_71_2381 ();
 sg13g2_fill_2 FILLER_71_2385 ();
 sg13g2_decap_4 FILLER_71_2395 ();
 sg13g2_fill_2 FILLER_71_2399 ();
 sg13g2_decap_4 FILLER_71_2419 ();
 sg13g2_fill_1 FILLER_71_2432 ();
 sg13g2_fill_2 FILLER_71_2445 ();
 sg13g2_fill_2 FILLER_71_2479 ();
 sg13g2_decap_8 FILLER_71_2526 ();
 sg13g2_decap_8 FILLER_71_2533 ();
 sg13g2_decap_8 FILLER_71_2540 ();
 sg13g2_decap_8 FILLER_71_2547 ();
 sg13g2_decap_8 FILLER_71_2554 ();
 sg13g2_fill_2 FILLER_71_2561 ();
 sg13g2_fill_1 FILLER_71_2578 ();
 sg13g2_fill_1 FILLER_71_2591 ();
 sg13g2_fill_2 FILLER_71_2606 ();
 sg13g2_fill_1 FILLER_71_2608 ();
 sg13g2_fill_2 FILLER_71_2637 ();
 sg13g2_fill_1 FILLER_71_2639 ();
 sg13g2_decap_4 FILLER_71_2650 ();
 sg13g2_fill_1 FILLER_71_2654 ();
 sg13g2_decap_4 FILLER_71_2658 ();
 sg13g2_fill_2 FILLER_71_2662 ();
 sg13g2_fill_2 FILLER_71_2669 ();
 sg13g2_decap_8 FILLER_71_2676 ();
 sg13g2_decap_8 FILLER_71_2683 ();
 sg13g2_decap_4 FILLER_71_2690 ();
 sg13g2_decap_4 FILLER_71_2710 ();
 sg13g2_fill_1 FILLER_71_2714 ();
 sg13g2_decap_8 FILLER_71_2728 ();
 sg13g2_fill_1 FILLER_71_2735 ();
 sg13g2_fill_2 FILLER_71_2749 ();
 sg13g2_fill_1 FILLER_71_2751 ();
 sg13g2_fill_2 FILLER_71_2757 ();
 sg13g2_decap_8 FILLER_71_2788 ();
 sg13g2_decap_4 FILLER_71_2795 ();
 sg13g2_fill_1 FILLER_71_2799 ();
 sg13g2_fill_1 FILLER_71_2812 ();
 sg13g2_decap_8 FILLER_71_2819 ();
 sg13g2_decap_8 FILLER_71_2839 ();
 sg13g2_fill_2 FILLER_71_2846 ();
 sg13g2_decap_8 FILLER_71_2864 ();
 sg13g2_fill_2 FILLER_71_2871 ();
 sg13g2_fill_1 FILLER_71_2873 ();
 sg13g2_fill_2 FILLER_71_2878 ();
 sg13g2_fill_1 FILLER_71_2880 ();
 sg13g2_decap_4 FILLER_71_2894 ();
 sg13g2_fill_1 FILLER_71_2898 ();
 sg13g2_decap_8 FILLER_71_2974 ();
 sg13g2_decap_8 FILLER_71_2981 ();
 sg13g2_decap_8 FILLER_71_2988 ();
 sg13g2_decap_8 FILLER_71_2995 ();
 sg13g2_decap_8 FILLER_71_3002 ();
 sg13g2_decap_8 FILLER_71_3009 ();
 sg13g2_decap_8 FILLER_71_3016 ();
 sg13g2_decap_8 FILLER_71_3023 ();
 sg13g2_decap_8 FILLER_71_3030 ();
 sg13g2_decap_8 FILLER_71_3037 ();
 sg13g2_decap_8 FILLER_71_3044 ();
 sg13g2_decap_8 FILLER_71_3051 ();
 sg13g2_decap_8 FILLER_71_3058 ();
 sg13g2_decap_8 FILLER_71_3065 ();
 sg13g2_decap_8 FILLER_71_3072 ();
 sg13g2_decap_8 FILLER_71_3079 ();
 sg13g2_decap_8 FILLER_71_3086 ();
 sg13g2_decap_8 FILLER_71_3093 ();
 sg13g2_decap_8 FILLER_71_3100 ();
 sg13g2_decap_8 FILLER_71_3107 ();
 sg13g2_decap_8 FILLER_71_3114 ();
 sg13g2_decap_8 FILLER_71_3121 ();
 sg13g2_decap_8 FILLER_71_3128 ();
 sg13g2_decap_8 FILLER_71_3135 ();
 sg13g2_decap_8 FILLER_71_3142 ();
 sg13g2_decap_8 FILLER_71_3149 ();
 sg13g2_decap_8 FILLER_71_3156 ();
 sg13g2_decap_8 FILLER_71_3163 ();
 sg13g2_decap_8 FILLER_71_3170 ();
 sg13g2_decap_8 FILLER_71_3177 ();
 sg13g2_decap_8 FILLER_71_3184 ();
 sg13g2_decap_8 FILLER_71_3191 ();
 sg13g2_decap_8 FILLER_71_3198 ();
 sg13g2_decap_8 FILLER_71_3205 ();
 sg13g2_decap_8 FILLER_71_3212 ();
 sg13g2_decap_8 FILLER_71_3219 ();
 sg13g2_decap_8 FILLER_71_3226 ();
 sg13g2_decap_8 FILLER_71_3233 ();
 sg13g2_decap_8 FILLER_71_3240 ();
 sg13g2_decap_8 FILLER_71_3247 ();
 sg13g2_decap_8 FILLER_71_3254 ();
 sg13g2_decap_8 FILLER_71_3261 ();
 sg13g2_decap_8 FILLER_71_3268 ();
 sg13g2_decap_8 FILLER_71_3275 ();
 sg13g2_decap_8 FILLER_71_3282 ();
 sg13g2_decap_8 FILLER_71_3289 ();
 sg13g2_decap_8 FILLER_71_3296 ();
 sg13g2_decap_8 FILLER_71_3303 ();
 sg13g2_decap_8 FILLER_71_3310 ();
 sg13g2_decap_8 FILLER_71_3317 ();
 sg13g2_decap_8 FILLER_71_3324 ();
 sg13g2_decap_8 FILLER_71_3331 ();
 sg13g2_decap_8 FILLER_71_3338 ();
 sg13g2_decap_8 FILLER_71_3345 ();
 sg13g2_decap_8 FILLER_71_3352 ();
 sg13g2_decap_8 FILLER_71_3359 ();
 sg13g2_decap_8 FILLER_71_3366 ();
 sg13g2_decap_8 FILLER_71_3373 ();
 sg13g2_decap_8 FILLER_71_3380 ();
 sg13g2_decap_8 FILLER_71_3387 ();
 sg13g2_decap_8 FILLER_71_3394 ();
 sg13g2_decap_8 FILLER_71_3401 ();
 sg13g2_decap_8 FILLER_71_3408 ();
 sg13g2_decap_8 FILLER_71_3415 ();
 sg13g2_decap_8 FILLER_71_3422 ();
 sg13g2_decap_8 FILLER_71_3429 ();
 sg13g2_decap_8 FILLER_71_3436 ();
 sg13g2_decap_8 FILLER_71_3443 ();
 sg13g2_decap_8 FILLER_71_3450 ();
 sg13g2_decap_8 FILLER_71_3457 ();
 sg13g2_decap_8 FILLER_71_3464 ();
 sg13g2_decap_8 FILLER_71_3471 ();
 sg13g2_decap_8 FILLER_71_3478 ();
 sg13g2_decap_8 FILLER_71_3485 ();
 sg13g2_decap_8 FILLER_71_3492 ();
 sg13g2_decap_8 FILLER_71_3499 ();
 sg13g2_decap_8 FILLER_71_3506 ();
 sg13g2_decap_8 FILLER_71_3513 ();
 sg13g2_decap_8 FILLER_71_3520 ();
 sg13g2_decap_8 FILLER_71_3527 ();
 sg13g2_decap_8 FILLER_71_3534 ();
 sg13g2_decap_8 FILLER_71_3541 ();
 sg13g2_decap_8 FILLER_71_3548 ();
 sg13g2_decap_8 FILLER_71_3555 ();
 sg13g2_decap_8 FILLER_71_3562 ();
 sg13g2_decap_8 FILLER_71_3569 ();
 sg13g2_decap_4 FILLER_71_3576 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_fill_2 FILLER_72_35 ();
 sg13g2_fill_2 FILLER_72_55 ();
 sg13g2_fill_2 FILLER_72_100 ();
 sg13g2_fill_1 FILLER_72_150 ();
 sg13g2_decap_8 FILLER_72_155 ();
 sg13g2_fill_2 FILLER_72_162 ();
 sg13g2_fill_1 FILLER_72_164 ();
 sg13g2_fill_1 FILLER_72_175 ();
 sg13g2_fill_2 FILLER_72_190 ();
 sg13g2_decap_8 FILLER_72_201 ();
 sg13g2_decap_8 FILLER_72_208 ();
 sg13g2_decap_4 FILLER_72_219 ();
 sg13g2_decap_8 FILLER_72_263 ();
 sg13g2_fill_2 FILLER_72_293 ();
 sg13g2_fill_1 FILLER_72_295 ();
 sg13g2_fill_2 FILLER_72_327 ();
 sg13g2_fill_1 FILLER_72_329 ();
 sg13g2_decap_4 FILLER_72_335 ();
 sg13g2_fill_1 FILLER_72_353 ();
 sg13g2_fill_2 FILLER_72_385 ();
 sg13g2_fill_1 FILLER_72_387 ();
 sg13g2_decap_8 FILLER_72_405 ();
 sg13g2_fill_2 FILLER_72_412 ();
 sg13g2_fill_1 FILLER_72_420 ();
 sg13g2_fill_2 FILLER_72_426 ();
 sg13g2_fill_1 FILLER_72_428 ();
 sg13g2_decap_8 FILLER_72_469 ();
 sg13g2_fill_1 FILLER_72_476 ();
 sg13g2_decap_8 FILLER_72_481 ();
 sg13g2_fill_2 FILLER_72_488 ();
 sg13g2_fill_1 FILLER_72_490 ();
 sg13g2_fill_1 FILLER_72_499 ();
 sg13g2_decap_8 FILLER_72_513 ();
 sg13g2_decap_8 FILLER_72_520 ();
 sg13g2_fill_2 FILLER_72_555 ();
 sg13g2_fill_1 FILLER_72_557 ();
 sg13g2_fill_1 FILLER_72_567 ();
 sg13g2_decap_8 FILLER_72_581 ();
 sg13g2_fill_2 FILLER_72_588 ();
 sg13g2_fill_1 FILLER_72_590 ();
 sg13g2_fill_1 FILLER_72_600 ();
 sg13g2_decap_8 FILLER_72_646 ();
 sg13g2_decap_4 FILLER_72_653 ();
 sg13g2_decap_4 FILLER_72_668 ();
 sg13g2_fill_2 FILLER_72_672 ();
 sg13g2_fill_2 FILLER_72_679 ();
 sg13g2_fill_1 FILLER_72_696 ();
 sg13g2_fill_1 FILLER_72_746 ();
 sg13g2_fill_2 FILLER_72_751 ();
 sg13g2_decap_4 FILLER_72_776 ();
 sg13g2_fill_1 FILLER_72_780 ();
 sg13g2_fill_1 FILLER_72_785 ();
 sg13g2_decap_4 FILLER_72_790 ();
 sg13g2_fill_2 FILLER_72_846 ();
 sg13g2_fill_1 FILLER_72_848 ();
 sg13g2_fill_2 FILLER_72_875 ();
 sg13g2_fill_2 FILLER_72_894 ();
 sg13g2_decap_4 FILLER_72_910 ();
 sg13g2_fill_2 FILLER_72_949 ();
 sg13g2_fill_1 FILLER_72_951 ();
 sg13g2_fill_1 FILLER_72_974 ();
 sg13g2_fill_2 FILLER_72_989 ();
 sg13g2_fill_1 FILLER_72_991 ();
 sg13g2_fill_2 FILLER_72_1023 ();
 sg13g2_decap_8 FILLER_72_1051 ();
 sg13g2_decap_4 FILLER_72_1058 ();
 sg13g2_decap_4 FILLER_72_1066 ();
 sg13g2_decap_8 FILLER_72_1076 ();
 sg13g2_decap_4 FILLER_72_1083 ();
 sg13g2_fill_2 FILLER_72_1087 ();
 sg13g2_fill_2 FILLER_72_1101 ();
 sg13g2_fill_1 FILLER_72_1103 ();
 sg13g2_decap_4 FILLER_72_1109 ();
 sg13g2_fill_1 FILLER_72_1113 ();
 sg13g2_decap_8 FILLER_72_1142 ();
 sg13g2_decap_8 FILLER_72_1149 ();
 sg13g2_decap_8 FILLER_72_1160 ();
 sg13g2_fill_2 FILLER_72_1167 ();
 sg13g2_fill_1 FILLER_72_1169 ();
 sg13g2_decap_4 FILLER_72_1196 ();
 sg13g2_fill_1 FILLER_72_1200 ();
 sg13g2_fill_2 FILLER_72_1250 ();
 sg13g2_fill_1 FILLER_72_1252 ();
 sg13g2_fill_1 FILLER_72_1291 ();
 sg13g2_fill_2 FILLER_72_1301 ();
 sg13g2_fill_1 FILLER_72_1303 ();
 sg13g2_fill_2 FILLER_72_1320 ();
 sg13g2_fill_1 FILLER_72_1322 ();
 sg13g2_fill_2 FILLER_72_1335 ();
 sg13g2_fill_1 FILLER_72_1381 ();
 sg13g2_fill_1 FILLER_72_1412 ();
 sg13g2_fill_2 FILLER_72_1422 ();
 sg13g2_fill_1 FILLER_72_1424 ();
 sg13g2_fill_1 FILLER_72_1441 ();
 sg13g2_fill_2 FILLER_72_1473 ();
 sg13g2_fill_2 FILLER_72_1531 ();
 sg13g2_fill_1 FILLER_72_1533 ();
 sg13g2_fill_1 FILLER_72_1539 ();
 sg13g2_fill_2 FILLER_72_1614 ();
 sg13g2_decap_8 FILLER_72_1659 ();
 sg13g2_decap_4 FILLER_72_1666 ();
 sg13g2_fill_1 FILLER_72_1670 ();
 sg13g2_decap_4 FILLER_72_1675 ();
 sg13g2_fill_1 FILLER_72_1679 ();
 sg13g2_fill_2 FILLER_72_1686 ();
 sg13g2_fill_2 FILLER_72_1732 ();
 sg13g2_fill_1 FILLER_72_1734 ();
 sg13g2_decap_8 FILLER_72_1765 ();
 sg13g2_decap_8 FILLER_72_1772 ();
 sg13g2_decap_8 FILLER_72_1779 ();
 sg13g2_decap_8 FILLER_72_1797 ();
 sg13g2_fill_2 FILLER_72_1804 ();
 sg13g2_fill_1 FILLER_72_1806 ();
 sg13g2_decap_8 FILLER_72_1824 ();
 sg13g2_fill_2 FILLER_72_1831 ();
 sg13g2_fill_2 FILLER_72_1869 ();
 sg13g2_fill_1 FILLER_72_1871 ();
 sg13g2_decap_8 FILLER_72_1921 ();
 sg13g2_decap_8 FILLER_72_1928 ();
 sg13g2_fill_2 FILLER_72_1935 ();
 sg13g2_fill_1 FILLER_72_1937 ();
 sg13g2_fill_2 FILLER_72_1948 ();
 sg13g2_fill_2 FILLER_72_1959 ();
 sg13g2_decap_4 FILLER_72_1979 ();
 sg13g2_fill_2 FILLER_72_2002 ();
 sg13g2_fill_2 FILLER_72_2030 ();
 sg13g2_fill_1 FILLER_72_2032 ();
 sg13g2_fill_1 FILLER_72_2095 ();
 sg13g2_decap_4 FILLER_72_2112 ();
 sg13g2_fill_1 FILLER_72_2121 ();
 sg13g2_fill_2 FILLER_72_2130 ();
 sg13g2_fill_1 FILLER_72_2132 ();
 sg13g2_decap_8 FILLER_72_2168 ();
 sg13g2_fill_1 FILLER_72_2175 ();
 sg13g2_fill_2 FILLER_72_2181 ();
 sg13g2_fill_1 FILLER_72_2183 ();
 sg13g2_decap_8 FILLER_72_2188 ();
 sg13g2_decap_8 FILLER_72_2195 ();
 sg13g2_decap_8 FILLER_72_2220 ();
 sg13g2_fill_2 FILLER_72_2227 ();
 sg13g2_fill_2 FILLER_72_2252 ();
 sg13g2_fill_2 FILLER_72_2272 ();
 sg13g2_fill_2 FILLER_72_2279 ();
 sg13g2_fill_1 FILLER_72_2281 ();
 sg13g2_fill_2 FILLER_72_2305 ();
 sg13g2_fill_1 FILLER_72_2307 ();
 sg13g2_decap_4 FILLER_72_2360 ();
 sg13g2_fill_2 FILLER_72_2364 ();
 sg13g2_decap_8 FILLER_72_2370 ();
 sg13g2_decap_8 FILLER_72_2377 ();
 sg13g2_fill_2 FILLER_72_2384 ();
 sg13g2_fill_1 FILLER_72_2386 ();
 sg13g2_fill_2 FILLER_72_2397 ();
 sg13g2_fill_1 FILLER_72_2404 ();
 sg13g2_fill_2 FILLER_72_2423 ();
 sg13g2_fill_1 FILLER_72_2425 ();
 sg13g2_decap_8 FILLER_72_2492 ();
 sg13g2_decap_4 FILLER_72_2499 ();
 sg13g2_decap_8 FILLER_72_2516 ();
 sg13g2_decap_4 FILLER_72_2523 ();
 sg13g2_fill_1 FILLER_72_2527 ();
 sg13g2_fill_1 FILLER_72_2562 ();
 sg13g2_fill_1 FILLER_72_2568 ();
 sg13g2_fill_1 FILLER_72_2580 ();
 sg13g2_fill_1 FILLER_72_2591 ();
 sg13g2_fill_1 FILLER_72_2597 ();
 sg13g2_decap_4 FILLER_72_2602 ();
 sg13g2_fill_2 FILLER_72_2611 ();
 sg13g2_fill_1 FILLER_72_2613 ();
 sg13g2_fill_1 FILLER_72_2618 ();
 sg13g2_fill_1 FILLER_72_2623 ();
 sg13g2_fill_2 FILLER_72_2629 ();
 sg13g2_fill_1 FILLER_72_2631 ();
 sg13g2_fill_2 FILLER_72_2687 ();
 sg13g2_fill_1 FILLER_72_2689 ();
 sg13g2_fill_1 FILLER_72_2700 ();
 sg13g2_fill_2 FILLER_72_2710 ();
 sg13g2_fill_1 FILLER_72_2712 ();
 sg13g2_fill_1 FILLER_72_2723 ();
 sg13g2_decap_4 FILLER_72_2729 ();
 sg13g2_fill_1 FILLER_72_2733 ();
 sg13g2_decap_4 FILLER_72_2743 ();
 sg13g2_fill_1 FILLER_72_2747 ();
 sg13g2_decap_4 FILLER_72_2778 ();
 sg13g2_fill_2 FILLER_72_2782 ();
 sg13g2_fill_2 FILLER_72_2791 ();
 sg13g2_fill_2 FILLER_72_2798 ();
 sg13g2_fill_1 FILLER_72_2800 ();
 sg13g2_fill_2 FILLER_72_2814 ();
 sg13g2_fill_2 FILLER_72_2884 ();
 sg13g2_decap_8 FILLER_72_2899 ();
 sg13g2_fill_2 FILLER_72_2906 ();
 sg13g2_fill_2 FILLER_72_2919 ();
 sg13g2_decap_8 FILLER_72_2926 ();
 sg13g2_fill_2 FILLER_72_2952 ();
 sg13g2_decap_8 FILLER_72_2967 ();
 sg13g2_decap_8 FILLER_72_2974 ();
 sg13g2_decap_8 FILLER_72_2981 ();
 sg13g2_decap_8 FILLER_72_2988 ();
 sg13g2_decap_8 FILLER_72_2995 ();
 sg13g2_decap_8 FILLER_72_3002 ();
 sg13g2_decap_8 FILLER_72_3009 ();
 sg13g2_decap_8 FILLER_72_3016 ();
 sg13g2_decap_8 FILLER_72_3023 ();
 sg13g2_decap_8 FILLER_72_3030 ();
 sg13g2_decap_8 FILLER_72_3037 ();
 sg13g2_decap_8 FILLER_72_3044 ();
 sg13g2_decap_8 FILLER_72_3051 ();
 sg13g2_decap_8 FILLER_72_3058 ();
 sg13g2_decap_8 FILLER_72_3065 ();
 sg13g2_decap_8 FILLER_72_3072 ();
 sg13g2_decap_8 FILLER_72_3079 ();
 sg13g2_decap_8 FILLER_72_3086 ();
 sg13g2_decap_8 FILLER_72_3093 ();
 sg13g2_decap_8 FILLER_72_3100 ();
 sg13g2_decap_8 FILLER_72_3107 ();
 sg13g2_decap_8 FILLER_72_3114 ();
 sg13g2_decap_8 FILLER_72_3121 ();
 sg13g2_decap_8 FILLER_72_3128 ();
 sg13g2_decap_8 FILLER_72_3135 ();
 sg13g2_decap_8 FILLER_72_3142 ();
 sg13g2_decap_8 FILLER_72_3149 ();
 sg13g2_decap_8 FILLER_72_3156 ();
 sg13g2_decap_8 FILLER_72_3163 ();
 sg13g2_decap_8 FILLER_72_3170 ();
 sg13g2_decap_8 FILLER_72_3177 ();
 sg13g2_decap_8 FILLER_72_3184 ();
 sg13g2_decap_8 FILLER_72_3191 ();
 sg13g2_decap_8 FILLER_72_3198 ();
 sg13g2_decap_8 FILLER_72_3205 ();
 sg13g2_decap_8 FILLER_72_3212 ();
 sg13g2_decap_8 FILLER_72_3219 ();
 sg13g2_decap_8 FILLER_72_3226 ();
 sg13g2_decap_8 FILLER_72_3233 ();
 sg13g2_decap_8 FILLER_72_3240 ();
 sg13g2_decap_8 FILLER_72_3247 ();
 sg13g2_decap_8 FILLER_72_3254 ();
 sg13g2_decap_8 FILLER_72_3261 ();
 sg13g2_decap_8 FILLER_72_3268 ();
 sg13g2_decap_8 FILLER_72_3275 ();
 sg13g2_decap_8 FILLER_72_3282 ();
 sg13g2_decap_8 FILLER_72_3289 ();
 sg13g2_decap_8 FILLER_72_3296 ();
 sg13g2_decap_8 FILLER_72_3303 ();
 sg13g2_decap_8 FILLER_72_3310 ();
 sg13g2_decap_8 FILLER_72_3317 ();
 sg13g2_decap_8 FILLER_72_3324 ();
 sg13g2_decap_8 FILLER_72_3331 ();
 sg13g2_decap_8 FILLER_72_3338 ();
 sg13g2_decap_8 FILLER_72_3345 ();
 sg13g2_decap_8 FILLER_72_3352 ();
 sg13g2_decap_8 FILLER_72_3359 ();
 sg13g2_decap_8 FILLER_72_3366 ();
 sg13g2_decap_8 FILLER_72_3373 ();
 sg13g2_decap_8 FILLER_72_3380 ();
 sg13g2_decap_8 FILLER_72_3387 ();
 sg13g2_decap_8 FILLER_72_3394 ();
 sg13g2_decap_8 FILLER_72_3401 ();
 sg13g2_decap_8 FILLER_72_3408 ();
 sg13g2_decap_8 FILLER_72_3415 ();
 sg13g2_decap_8 FILLER_72_3422 ();
 sg13g2_decap_8 FILLER_72_3429 ();
 sg13g2_decap_8 FILLER_72_3436 ();
 sg13g2_decap_8 FILLER_72_3443 ();
 sg13g2_decap_8 FILLER_72_3450 ();
 sg13g2_decap_8 FILLER_72_3457 ();
 sg13g2_decap_8 FILLER_72_3464 ();
 sg13g2_decap_8 FILLER_72_3471 ();
 sg13g2_decap_8 FILLER_72_3478 ();
 sg13g2_decap_8 FILLER_72_3485 ();
 sg13g2_decap_8 FILLER_72_3492 ();
 sg13g2_decap_8 FILLER_72_3499 ();
 sg13g2_decap_8 FILLER_72_3506 ();
 sg13g2_decap_8 FILLER_72_3513 ();
 sg13g2_decap_8 FILLER_72_3520 ();
 sg13g2_decap_8 FILLER_72_3527 ();
 sg13g2_decap_8 FILLER_72_3534 ();
 sg13g2_decap_8 FILLER_72_3541 ();
 sg13g2_decap_8 FILLER_72_3548 ();
 sg13g2_decap_8 FILLER_72_3555 ();
 sg13g2_decap_8 FILLER_72_3562 ();
 sg13g2_decap_8 FILLER_72_3569 ();
 sg13g2_decap_4 FILLER_72_3576 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_88 ();
 sg13g2_decap_4 FILLER_73_95 ();
 sg13g2_fill_1 FILLER_73_99 ();
 sg13g2_decap_4 FILLER_73_104 ();
 sg13g2_fill_2 FILLER_73_108 ();
 sg13g2_fill_2 FILLER_73_167 ();
 sg13g2_fill_1 FILLER_73_169 ();
 sg13g2_fill_2 FILLER_73_183 ();
 sg13g2_decap_8 FILLER_73_231 ();
 sg13g2_fill_2 FILLER_73_238 ();
 sg13g2_fill_1 FILLER_73_240 ();
 sg13g2_decap_4 FILLER_73_246 ();
 sg13g2_fill_2 FILLER_73_259 ();
 sg13g2_decap_8 FILLER_73_360 ();
 sg13g2_decap_8 FILLER_73_380 ();
 sg13g2_fill_2 FILLER_73_387 ();
 sg13g2_decap_8 FILLER_73_399 ();
 sg13g2_decap_8 FILLER_73_406 ();
 sg13g2_fill_2 FILLER_73_413 ();
 sg13g2_fill_1 FILLER_73_439 ();
 sg13g2_fill_2 FILLER_73_458 ();
 sg13g2_fill_2 FILLER_73_469 ();
 sg13g2_fill_1 FILLER_73_471 ();
 sg13g2_decap_4 FILLER_73_498 ();
 sg13g2_fill_1 FILLER_73_502 ();
 sg13g2_fill_2 FILLER_73_598 ();
 sg13g2_decap_8 FILLER_73_605 ();
 sg13g2_fill_2 FILLER_73_628 ();
 sg13g2_fill_1 FILLER_73_654 ();
 sg13g2_fill_1 FILLER_73_674 ();
 sg13g2_fill_1 FILLER_73_683 ();
 sg13g2_fill_1 FILLER_73_703 ();
 sg13g2_fill_2 FILLER_73_722 ();
 sg13g2_fill_1 FILLER_73_724 ();
 sg13g2_fill_1 FILLER_73_744 ();
 sg13g2_fill_2 FILLER_73_774 ();
 sg13g2_fill_1 FILLER_73_776 ();
 sg13g2_decap_8 FILLER_73_803 ();
 sg13g2_decap_8 FILLER_73_810 ();
 sg13g2_decap_4 FILLER_73_825 ();
 sg13g2_decap_8 FILLER_73_847 ();
 sg13g2_fill_2 FILLER_73_871 ();
 sg13g2_decap_8 FILLER_73_916 ();
 sg13g2_fill_2 FILLER_73_923 ();
 sg13g2_decap_4 FILLER_73_929 ();
 sg13g2_fill_2 FILLER_73_933 ();
 sg13g2_decap_8 FILLER_73_939 ();
 sg13g2_decap_8 FILLER_73_946 ();
 sg13g2_fill_2 FILLER_73_953 ();
 sg13g2_fill_1 FILLER_73_955 ();
 sg13g2_decap_8 FILLER_73_961 ();
 sg13g2_fill_1 FILLER_73_968 ();
 sg13g2_fill_2 FILLER_73_974 ();
 sg13g2_fill_1 FILLER_73_979 ();
 sg13g2_fill_2 FILLER_73_990 ();
 sg13g2_fill_2 FILLER_73_1000 ();
 sg13g2_fill_2 FILLER_73_1011 ();
 sg13g2_fill_1 FILLER_73_1013 ();
 sg13g2_fill_2 FILLER_73_1023 ();
 sg13g2_decap_4 FILLER_73_1030 ();
 sg13g2_fill_2 FILLER_73_1034 ();
 sg13g2_decap_8 FILLER_73_1040 ();
 sg13g2_decap_4 FILLER_73_1047 ();
 sg13g2_fill_1 FILLER_73_1051 ();
 sg13g2_fill_2 FILLER_73_1078 ();
 sg13g2_fill_1 FILLER_73_1080 ();
 sg13g2_fill_1 FILLER_73_1086 ();
 sg13g2_fill_2 FILLER_73_1097 ();
 sg13g2_decap_8 FILLER_73_1138 ();
 sg13g2_fill_2 FILLER_73_1145 ();
 sg13g2_fill_1 FILLER_73_1147 ();
 sg13g2_decap_4 FILLER_73_1153 ();
 sg13g2_fill_1 FILLER_73_1157 ();
 sg13g2_fill_1 FILLER_73_1189 ();
 sg13g2_decap_8 FILLER_73_1203 ();
 sg13g2_decap_8 FILLER_73_1210 ();
 sg13g2_fill_2 FILLER_73_1217 ();
 sg13g2_fill_2 FILLER_73_1245 ();
 sg13g2_fill_1 FILLER_73_1252 ();
 sg13g2_fill_2 FILLER_73_1268 ();
 sg13g2_fill_2 FILLER_73_1284 ();
 sg13g2_fill_1 FILLER_73_1313 ();
 sg13g2_decap_8 FILLER_73_1346 ();
 sg13g2_decap_8 FILLER_73_1353 ();
 sg13g2_fill_1 FILLER_73_1360 ();
 sg13g2_fill_2 FILLER_73_1365 ();
 sg13g2_decap_4 FILLER_73_1371 ();
 sg13g2_fill_1 FILLER_73_1375 ();
 sg13g2_fill_2 FILLER_73_1385 ();
 sg13g2_decap_8 FILLER_73_1392 ();
 sg13g2_fill_1 FILLER_73_1399 ();
 sg13g2_fill_2 FILLER_73_1406 ();
 sg13g2_fill_2 FILLER_73_1434 ();
 sg13g2_fill_1 FILLER_73_1453 ();
 sg13g2_fill_1 FILLER_73_1462 ();
 sg13g2_decap_8 FILLER_73_1472 ();
 sg13g2_decap_4 FILLER_73_1479 ();
 sg13g2_fill_2 FILLER_73_1483 ();
 sg13g2_fill_2 FILLER_73_1489 ();
 sg13g2_fill_1 FILLER_73_1491 ();
 sg13g2_fill_1 FILLER_73_1518 ();
 sg13g2_fill_2 FILLER_73_1540 ();
 sg13g2_fill_2 FILLER_73_1558 ();
 sg13g2_fill_1 FILLER_73_1560 ();
 sg13g2_decap_4 FILLER_73_1565 ();
 sg13g2_fill_1 FILLER_73_1569 ();
 sg13g2_fill_2 FILLER_73_1580 ();
 sg13g2_fill_2 FILLER_73_1617 ();
 sg13g2_fill_2 FILLER_73_1624 ();
 sg13g2_fill_1 FILLER_73_1626 ();
 sg13g2_fill_1 FILLER_73_1635 ();
 sg13g2_decap_8 FILLER_73_1667 ();
 sg13g2_decap_4 FILLER_73_1674 ();
 sg13g2_fill_1 FILLER_73_1678 ();
 sg13g2_decap_4 FILLER_73_1683 ();
 sg13g2_fill_2 FILLER_73_1687 ();
 sg13g2_fill_2 FILLER_73_1695 ();
 sg13g2_fill_1 FILLER_73_1697 ();
 sg13g2_decap_8 FILLER_73_1709 ();
 sg13g2_decap_4 FILLER_73_1716 ();
 sg13g2_fill_2 FILLER_73_1720 ();
 sg13g2_fill_2 FILLER_73_1757 ();
 sg13g2_fill_1 FILLER_73_1759 ();
 sg13g2_fill_1 FILLER_73_1786 ();
 sg13g2_decap_8 FILLER_73_1804 ();
 sg13g2_decap_4 FILLER_73_1811 ();
 sg13g2_decap_8 FILLER_73_1830 ();
 sg13g2_fill_2 FILLER_73_1837 ();
 sg13g2_fill_2 FILLER_73_1844 ();
 sg13g2_decap_8 FILLER_73_1850 ();
 sg13g2_fill_2 FILLER_73_1857 ();
 sg13g2_fill_1 FILLER_73_1859 ();
 sg13g2_decap_8 FILLER_73_1875 ();
 sg13g2_fill_2 FILLER_73_1882 ();
 sg13g2_fill_1 FILLER_73_1938 ();
 sg13g2_fill_2 FILLER_73_1991 ();
 sg13g2_fill_1 FILLER_73_1993 ();
 sg13g2_decap_4 FILLER_73_2039 ();
 sg13g2_fill_1 FILLER_73_2043 ();
 sg13g2_fill_1 FILLER_73_2060 ();
 sg13g2_fill_2 FILLER_73_2087 ();
 sg13g2_fill_1 FILLER_73_2089 ();
 sg13g2_fill_2 FILLER_73_2099 ();
 sg13g2_decap_8 FILLER_73_2111 ();
 sg13g2_fill_2 FILLER_73_2118 ();
 sg13g2_decap_4 FILLER_73_2127 ();
 sg13g2_decap_8 FILLER_73_2161 ();
 sg13g2_decap_4 FILLER_73_2168 ();
 sg13g2_fill_2 FILLER_73_2172 ();
 sg13g2_decap_4 FILLER_73_2200 ();
 sg13g2_fill_2 FILLER_73_2204 ();
 sg13g2_decap_4 FILLER_73_2224 ();
 sg13g2_fill_1 FILLER_73_2228 ();
 sg13g2_fill_2 FILLER_73_2317 ();
 sg13g2_decap_4 FILLER_73_2327 ();
 sg13g2_fill_1 FILLER_73_2331 ();
 sg13g2_decap_8 FILLER_73_2337 ();
 sg13g2_decap_8 FILLER_73_2344 ();
 sg13g2_fill_2 FILLER_73_2356 ();
 sg13g2_decap_8 FILLER_73_2363 ();
 sg13g2_decap_4 FILLER_73_2370 ();
 sg13g2_fill_1 FILLER_73_2374 ();
 sg13g2_fill_2 FILLER_73_2391 ();
 sg13g2_fill_1 FILLER_73_2393 ();
 sg13g2_decap_8 FILLER_73_2398 ();
 sg13g2_fill_2 FILLER_73_2405 ();
 sg13g2_decap_4 FILLER_73_2412 ();
 sg13g2_decap_4 FILLER_73_2420 ();
 sg13g2_fill_1 FILLER_73_2474 ();
 sg13g2_fill_2 FILLER_73_2497 ();
 sg13g2_fill_1 FILLER_73_2499 ();
 sg13g2_decap_8 FILLER_73_2531 ();
 sg13g2_decap_8 FILLER_73_2542 ();
 sg13g2_fill_2 FILLER_73_2562 ();
 sg13g2_fill_2 FILLER_73_2591 ();
 sg13g2_fill_2 FILLER_73_2603 ();
 sg13g2_decap_8 FILLER_73_2635 ();
 sg13g2_fill_1 FILLER_73_2642 ();
 sg13g2_decap_4 FILLER_73_2648 ();
 sg13g2_fill_1 FILLER_73_2652 ();
 sg13g2_fill_2 FILLER_73_2657 ();
 sg13g2_fill_1 FILLER_73_2659 ();
 sg13g2_fill_2 FILLER_73_2679 ();
 sg13g2_fill_1 FILLER_73_2681 ();
 sg13g2_fill_2 FILLER_73_2696 ();
 sg13g2_fill_1 FILLER_73_2698 ();
 sg13g2_fill_1 FILLER_73_2704 ();
 sg13g2_fill_2 FILLER_73_2725 ();
 sg13g2_fill_1 FILLER_73_2727 ();
 sg13g2_fill_2 FILLER_73_2741 ();
 sg13g2_fill_1 FILLER_73_2743 ();
 sg13g2_decap_8 FILLER_73_2752 ();
 sg13g2_fill_2 FILLER_73_2759 ();
 sg13g2_fill_1 FILLER_73_2761 ();
 sg13g2_fill_1 FILLER_73_2765 ();
 sg13g2_decap_8 FILLER_73_2770 ();
 sg13g2_fill_2 FILLER_73_2777 ();
 sg13g2_fill_1 FILLER_73_2779 ();
 sg13g2_fill_1 FILLER_73_2820 ();
 sg13g2_decap_8 FILLER_73_2829 ();
 sg13g2_decap_8 FILLER_73_2836 ();
 sg13g2_decap_8 FILLER_73_2843 ();
 sg13g2_fill_1 FILLER_73_2850 ();
 sg13g2_decap_8 FILLER_73_2859 ();
 sg13g2_fill_2 FILLER_73_2866 ();
 sg13g2_fill_1 FILLER_73_2868 ();
 sg13g2_decap_8 FILLER_73_2874 ();
 sg13g2_decap_8 FILLER_73_2881 ();
 sg13g2_decap_8 FILLER_73_2888 ();
 sg13g2_fill_2 FILLER_73_2895 ();
 sg13g2_fill_1 FILLER_73_2897 ();
 sg13g2_fill_1 FILLER_73_2902 ();
 sg13g2_fill_2 FILLER_73_2925 ();
 sg13g2_decap_8 FILLER_73_2953 ();
 sg13g2_decap_8 FILLER_73_2960 ();
 sg13g2_decap_8 FILLER_73_2967 ();
 sg13g2_decap_8 FILLER_73_2974 ();
 sg13g2_decap_8 FILLER_73_2981 ();
 sg13g2_decap_8 FILLER_73_2988 ();
 sg13g2_decap_8 FILLER_73_2995 ();
 sg13g2_decap_8 FILLER_73_3002 ();
 sg13g2_decap_8 FILLER_73_3009 ();
 sg13g2_decap_8 FILLER_73_3016 ();
 sg13g2_decap_8 FILLER_73_3023 ();
 sg13g2_decap_8 FILLER_73_3030 ();
 sg13g2_decap_8 FILLER_73_3037 ();
 sg13g2_decap_8 FILLER_73_3044 ();
 sg13g2_decap_8 FILLER_73_3051 ();
 sg13g2_decap_8 FILLER_73_3058 ();
 sg13g2_decap_8 FILLER_73_3065 ();
 sg13g2_decap_8 FILLER_73_3072 ();
 sg13g2_decap_8 FILLER_73_3079 ();
 sg13g2_decap_8 FILLER_73_3086 ();
 sg13g2_decap_8 FILLER_73_3093 ();
 sg13g2_decap_8 FILLER_73_3100 ();
 sg13g2_decap_8 FILLER_73_3107 ();
 sg13g2_decap_8 FILLER_73_3114 ();
 sg13g2_decap_8 FILLER_73_3121 ();
 sg13g2_decap_8 FILLER_73_3128 ();
 sg13g2_decap_8 FILLER_73_3135 ();
 sg13g2_decap_8 FILLER_73_3142 ();
 sg13g2_decap_8 FILLER_73_3149 ();
 sg13g2_decap_8 FILLER_73_3156 ();
 sg13g2_decap_8 FILLER_73_3163 ();
 sg13g2_decap_8 FILLER_73_3170 ();
 sg13g2_decap_8 FILLER_73_3177 ();
 sg13g2_decap_8 FILLER_73_3184 ();
 sg13g2_decap_8 FILLER_73_3191 ();
 sg13g2_decap_8 FILLER_73_3198 ();
 sg13g2_decap_8 FILLER_73_3205 ();
 sg13g2_decap_8 FILLER_73_3212 ();
 sg13g2_decap_8 FILLER_73_3219 ();
 sg13g2_decap_8 FILLER_73_3226 ();
 sg13g2_decap_8 FILLER_73_3233 ();
 sg13g2_decap_8 FILLER_73_3240 ();
 sg13g2_decap_8 FILLER_73_3247 ();
 sg13g2_decap_8 FILLER_73_3254 ();
 sg13g2_decap_8 FILLER_73_3261 ();
 sg13g2_decap_8 FILLER_73_3268 ();
 sg13g2_decap_8 FILLER_73_3275 ();
 sg13g2_decap_8 FILLER_73_3282 ();
 sg13g2_decap_8 FILLER_73_3289 ();
 sg13g2_decap_8 FILLER_73_3296 ();
 sg13g2_decap_8 FILLER_73_3303 ();
 sg13g2_decap_8 FILLER_73_3310 ();
 sg13g2_decap_8 FILLER_73_3317 ();
 sg13g2_decap_8 FILLER_73_3324 ();
 sg13g2_decap_8 FILLER_73_3331 ();
 sg13g2_decap_8 FILLER_73_3338 ();
 sg13g2_decap_8 FILLER_73_3345 ();
 sg13g2_decap_8 FILLER_73_3352 ();
 sg13g2_decap_8 FILLER_73_3359 ();
 sg13g2_decap_8 FILLER_73_3366 ();
 sg13g2_decap_8 FILLER_73_3373 ();
 sg13g2_decap_8 FILLER_73_3380 ();
 sg13g2_decap_8 FILLER_73_3387 ();
 sg13g2_decap_8 FILLER_73_3394 ();
 sg13g2_decap_8 FILLER_73_3401 ();
 sg13g2_decap_8 FILLER_73_3408 ();
 sg13g2_decap_8 FILLER_73_3415 ();
 sg13g2_decap_8 FILLER_73_3422 ();
 sg13g2_decap_8 FILLER_73_3429 ();
 sg13g2_decap_8 FILLER_73_3436 ();
 sg13g2_decap_8 FILLER_73_3443 ();
 sg13g2_decap_8 FILLER_73_3450 ();
 sg13g2_decap_8 FILLER_73_3457 ();
 sg13g2_decap_8 FILLER_73_3464 ();
 sg13g2_decap_8 FILLER_73_3471 ();
 sg13g2_decap_8 FILLER_73_3478 ();
 sg13g2_decap_8 FILLER_73_3485 ();
 sg13g2_decap_8 FILLER_73_3492 ();
 sg13g2_decap_8 FILLER_73_3499 ();
 sg13g2_decap_8 FILLER_73_3506 ();
 sg13g2_decap_8 FILLER_73_3513 ();
 sg13g2_decap_8 FILLER_73_3520 ();
 sg13g2_decap_8 FILLER_73_3527 ();
 sg13g2_decap_8 FILLER_73_3534 ();
 sg13g2_decap_8 FILLER_73_3541 ();
 sg13g2_decap_8 FILLER_73_3548 ();
 sg13g2_decap_8 FILLER_73_3555 ();
 sg13g2_decap_8 FILLER_73_3562 ();
 sg13g2_decap_8 FILLER_73_3569 ();
 sg13g2_decap_4 FILLER_73_3576 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_fill_2 FILLER_74_42 ();
 sg13g2_fill_1 FILLER_74_44 ();
 sg13g2_decap_8 FILLER_74_58 ();
 sg13g2_decap_8 FILLER_74_65 ();
 sg13g2_decap_8 FILLER_74_72 ();
 sg13g2_decap_8 FILLER_74_79 ();
 sg13g2_decap_4 FILLER_74_86 ();
 sg13g2_fill_2 FILLER_74_90 ();
 sg13g2_fill_1 FILLER_74_127 ();
 sg13g2_fill_1 FILLER_74_147 ();
 sg13g2_decap_8 FILLER_74_152 ();
 sg13g2_fill_2 FILLER_74_159 ();
 sg13g2_fill_2 FILLER_74_190 ();
 sg13g2_decap_4 FILLER_74_227 ();
 sg13g2_fill_2 FILLER_74_231 ();
 sg13g2_fill_2 FILLER_74_251 ();
 sg13g2_fill_2 FILLER_74_270 ();
 sg13g2_fill_2 FILLER_74_282 ();
 sg13g2_fill_1 FILLER_74_284 ();
 sg13g2_fill_2 FILLER_74_289 ();
 sg13g2_fill_2 FILLER_74_316 ();
 sg13g2_fill_1 FILLER_74_318 ();
 sg13g2_decap_4 FILLER_74_332 ();
 sg13g2_fill_2 FILLER_74_411 ();
 sg13g2_fill_1 FILLER_74_439 ();
 sg13g2_fill_2 FILLER_74_445 ();
 sg13g2_fill_1 FILLER_74_447 ();
 sg13g2_decap_8 FILLER_74_493 ();
 sg13g2_fill_1 FILLER_74_500 ();
 sg13g2_fill_1 FILLER_74_540 ();
 sg13g2_fill_1 FILLER_74_559 ();
 sg13g2_decap_8 FILLER_74_567 ();
 sg13g2_decap_4 FILLER_74_574 ();
 sg13g2_decap_8 FILLER_74_582 ();
 sg13g2_fill_2 FILLER_74_589 ();
 sg13g2_fill_1 FILLER_74_591 ();
 sg13g2_fill_2 FILLER_74_625 ();
 sg13g2_fill_1 FILLER_74_632 ();
 sg13g2_decap_8 FILLER_74_638 ();
 sg13g2_fill_1 FILLER_74_645 ();
 sg13g2_decap_8 FILLER_74_651 ();
 sg13g2_fill_2 FILLER_74_658 ();
 sg13g2_fill_1 FILLER_74_660 ();
 sg13g2_decap_4 FILLER_74_666 ();
 sg13g2_fill_2 FILLER_74_670 ();
 sg13g2_fill_1 FILLER_74_702 ();
 sg13g2_fill_2 FILLER_74_729 ();
 sg13g2_fill_1 FILLER_74_752 ();
 sg13g2_fill_2 FILLER_74_786 ();
 sg13g2_decap_4 FILLER_74_792 ();
 sg13g2_fill_2 FILLER_74_887 ();
 sg13g2_decap_4 FILLER_74_898 ();
 sg13g2_fill_2 FILLER_74_922 ();
 sg13g2_fill_1 FILLER_74_964 ();
 sg13g2_fill_2 FILLER_74_986 ();
 sg13g2_fill_1 FILLER_74_1014 ();
 sg13g2_fill_2 FILLER_74_1051 ();
 sg13g2_fill_1 FILLER_74_1053 ();
 sg13g2_fill_1 FILLER_74_1072 ();
 sg13g2_fill_2 FILLER_74_1078 ();
 sg13g2_decap_4 FILLER_74_1106 ();
 sg13g2_fill_2 FILLER_74_1155 ();
 sg13g2_fill_1 FILLER_74_1157 ();
 sg13g2_decap_8 FILLER_74_1217 ();
 sg13g2_fill_2 FILLER_74_1224 ();
 sg13g2_fill_1 FILLER_74_1226 ();
 sg13g2_fill_1 FILLER_74_1269 ();
 sg13g2_fill_1 FILLER_74_1280 ();
 sg13g2_decap_8 FILLER_74_1337 ();
 sg13g2_decap_4 FILLER_74_1344 ();
 sg13g2_fill_1 FILLER_74_1348 ();
 sg13g2_decap_8 FILLER_74_1353 ();
 sg13g2_fill_2 FILLER_74_1360 ();
 sg13g2_fill_1 FILLER_74_1362 ();
 sg13g2_fill_1 FILLER_74_1389 ();
 sg13g2_fill_1 FILLER_74_1395 ();
 sg13g2_fill_2 FILLER_74_1404 ();
 sg13g2_fill_2 FILLER_74_1412 ();
 sg13g2_fill_1 FILLER_74_1414 ();
 sg13g2_fill_2 FILLER_74_1441 ();
 sg13g2_fill_1 FILLER_74_1475 ();
 sg13g2_decap_4 FILLER_74_1516 ();
 sg13g2_fill_1 FILLER_74_1520 ();
 sg13g2_fill_1 FILLER_74_1540 ();
 sg13g2_fill_2 FILLER_74_1596 ();
 sg13g2_fill_2 FILLER_74_1606 ();
 sg13g2_fill_1 FILLER_74_1608 ();
 sg13g2_fill_2 FILLER_74_1694 ();
 sg13g2_fill_1 FILLER_74_1696 ();
 sg13g2_fill_2 FILLER_74_1706 ();
 sg13g2_fill_1 FILLER_74_1708 ();
 sg13g2_decap_8 FILLER_74_1761 ();
 sg13g2_fill_2 FILLER_74_1768 ();
 sg13g2_fill_1 FILLER_74_1770 ();
 sg13g2_decap_8 FILLER_74_1775 ();
 sg13g2_fill_2 FILLER_74_1782 ();
 sg13g2_fill_2 FILLER_74_1828 ();
 sg13g2_fill_1 FILLER_74_1830 ();
 sg13g2_decap_4 FILLER_74_1862 ();
 sg13g2_decap_8 FILLER_74_1877 ();
 sg13g2_fill_2 FILLER_74_1884 ();
 sg13g2_fill_1 FILLER_74_1886 ();
 sg13g2_fill_1 FILLER_74_1892 ();
 sg13g2_decap_4 FILLER_74_1903 ();
 sg13g2_fill_1 FILLER_74_1907 ();
 sg13g2_fill_2 FILLER_74_1937 ();
 sg13g2_fill_2 FILLER_74_1944 ();
 sg13g2_fill_1 FILLER_74_1946 ();
 sg13g2_decap_4 FILLER_74_1971 ();
 sg13g2_decap_8 FILLER_74_1979 ();
 sg13g2_fill_1 FILLER_74_1986 ();
 sg13g2_decap_8 FILLER_74_2017 ();
 sg13g2_decap_4 FILLER_74_2024 ();
 sg13g2_fill_2 FILLER_74_2028 ();
 sg13g2_fill_1 FILLER_74_2073 ();
 sg13g2_fill_2 FILLER_74_2095 ();
 sg13g2_decap_8 FILLER_74_2106 ();
 sg13g2_decap_4 FILLER_74_2113 ();
 sg13g2_fill_2 FILLER_74_2117 ();
 sg13g2_fill_2 FILLER_74_2142 ();
 sg13g2_fill_1 FILLER_74_2171 ();
 sg13g2_decap_8 FILLER_74_2176 ();
 sg13g2_decap_4 FILLER_74_2183 ();
 sg13g2_fill_2 FILLER_74_2187 ();
 sg13g2_fill_1 FILLER_74_2193 ();
 sg13g2_decap_4 FILLER_74_2199 ();
 sg13g2_fill_1 FILLER_74_2203 ();
 sg13g2_decap_8 FILLER_74_2208 ();
 sg13g2_fill_2 FILLER_74_2215 ();
 sg13g2_fill_1 FILLER_74_2225 ();
 sg13g2_decap_8 FILLER_74_2231 ();
 sg13g2_fill_2 FILLER_74_2238 ();
 sg13g2_decap_4 FILLER_74_2244 ();
 sg13g2_fill_2 FILLER_74_2248 ();
 sg13g2_decap_4 FILLER_74_2255 ();
 sg13g2_fill_1 FILLER_74_2259 ();
 sg13g2_decap_4 FILLER_74_2282 ();
 sg13g2_fill_2 FILLER_74_2286 ();
 sg13g2_fill_2 FILLER_74_2292 ();
 sg13g2_fill_1 FILLER_74_2320 ();
 sg13g2_fill_2 FILLER_74_2326 ();
 sg13g2_fill_2 FILLER_74_2338 ();
 sg13g2_fill_1 FILLER_74_2350 ();
 sg13g2_decap_8 FILLER_74_2377 ();
 sg13g2_fill_2 FILLER_74_2384 ();
 sg13g2_fill_1 FILLER_74_2386 ();
 sg13g2_fill_1 FILLER_74_2406 ();
 sg13g2_fill_1 FILLER_74_2412 ();
 sg13g2_fill_2 FILLER_74_2457 ();
 sg13g2_fill_1 FILLER_74_2465 ();
 sg13g2_decap_4 FILLER_74_2474 ();
 sg13g2_fill_1 FILLER_74_2504 ();
 sg13g2_decap_4 FILLER_74_2511 ();
 sg13g2_fill_1 FILLER_74_2515 ();
 sg13g2_decap_8 FILLER_74_2520 ();
 sg13g2_decap_4 FILLER_74_2527 ();
 sg13g2_fill_2 FILLER_74_2531 ();
 sg13g2_decap_8 FILLER_74_2537 ();
 sg13g2_fill_1 FILLER_74_2554 ();
 sg13g2_decap_8 FILLER_74_2594 ();
 sg13g2_decap_4 FILLER_74_2601 ();
 sg13g2_fill_1 FILLER_74_2605 ();
 sg13g2_decap_4 FILLER_74_2610 ();
 sg13g2_fill_1 FILLER_74_2614 ();
 sg13g2_decap_8 FILLER_74_2628 ();
 sg13g2_decap_4 FILLER_74_2635 ();
 sg13g2_fill_2 FILLER_74_2639 ();
 sg13g2_decap_8 FILLER_74_2648 ();
 sg13g2_decap_4 FILLER_74_2655 ();
 sg13g2_fill_1 FILLER_74_2664 ();
 sg13g2_decap_4 FILLER_74_2683 ();
 sg13g2_decap_8 FILLER_74_2692 ();
 sg13g2_decap_8 FILLER_74_2699 ();
 sg13g2_decap_4 FILLER_74_2706 ();
 sg13g2_fill_2 FILLER_74_2710 ();
 sg13g2_fill_2 FILLER_74_2726 ();
 sg13g2_decap_8 FILLER_74_2749 ();
 sg13g2_decap_4 FILLER_74_2756 ();
 sg13g2_decap_8 FILLER_74_2780 ();
 sg13g2_decap_4 FILLER_74_2787 ();
 sg13g2_decap_8 FILLER_74_2800 ();
 sg13g2_decap_4 FILLER_74_2807 ();
 sg13g2_fill_2 FILLER_74_2811 ();
 sg13g2_fill_2 FILLER_74_2821 ();
 sg13g2_fill_1 FILLER_74_2823 ();
 sg13g2_decap_8 FILLER_74_2839 ();
 sg13g2_fill_2 FILLER_74_2846 ();
 sg13g2_fill_1 FILLER_74_2848 ();
 sg13g2_decap_8 FILLER_74_2857 ();
 sg13g2_fill_2 FILLER_74_2864 ();
 sg13g2_fill_2 FILLER_74_2920 ();
 sg13g2_fill_2 FILLER_74_2935 ();
 sg13g2_fill_1 FILLER_74_2937 ();
 sg13g2_decap_8 FILLER_74_2942 ();
 sg13g2_decap_8 FILLER_74_2949 ();
 sg13g2_decap_8 FILLER_74_2956 ();
 sg13g2_decap_8 FILLER_74_2963 ();
 sg13g2_decap_8 FILLER_74_2970 ();
 sg13g2_decap_8 FILLER_74_2977 ();
 sg13g2_decap_8 FILLER_74_2984 ();
 sg13g2_decap_8 FILLER_74_2991 ();
 sg13g2_decap_8 FILLER_74_2998 ();
 sg13g2_decap_8 FILLER_74_3005 ();
 sg13g2_decap_8 FILLER_74_3012 ();
 sg13g2_decap_8 FILLER_74_3019 ();
 sg13g2_decap_8 FILLER_74_3026 ();
 sg13g2_decap_8 FILLER_74_3033 ();
 sg13g2_decap_8 FILLER_74_3040 ();
 sg13g2_decap_8 FILLER_74_3047 ();
 sg13g2_decap_8 FILLER_74_3054 ();
 sg13g2_decap_8 FILLER_74_3061 ();
 sg13g2_decap_8 FILLER_74_3068 ();
 sg13g2_decap_8 FILLER_74_3075 ();
 sg13g2_decap_8 FILLER_74_3082 ();
 sg13g2_decap_8 FILLER_74_3089 ();
 sg13g2_decap_8 FILLER_74_3096 ();
 sg13g2_decap_8 FILLER_74_3103 ();
 sg13g2_decap_8 FILLER_74_3110 ();
 sg13g2_decap_8 FILLER_74_3117 ();
 sg13g2_decap_8 FILLER_74_3124 ();
 sg13g2_decap_8 FILLER_74_3131 ();
 sg13g2_decap_8 FILLER_74_3138 ();
 sg13g2_decap_8 FILLER_74_3145 ();
 sg13g2_decap_8 FILLER_74_3152 ();
 sg13g2_decap_8 FILLER_74_3159 ();
 sg13g2_decap_8 FILLER_74_3166 ();
 sg13g2_decap_8 FILLER_74_3173 ();
 sg13g2_decap_8 FILLER_74_3180 ();
 sg13g2_decap_8 FILLER_74_3187 ();
 sg13g2_decap_8 FILLER_74_3194 ();
 sg13g2_decap_8 FILLER_74_3201 ();
 sg13g2_decap_8 FILLER_74_3208 ();
 sg13g2_decap_8 FILLER_74_3215 ();
 sg13g2_decap_8 FILLER_74_3222 ();
 sg13g2_decap_8 FILLER_74_3229 ();
 sg13g2_decap_8 FILLER_74_3236 ();
 sg13g2_decap_8 FILLER_74_3243 ();
 sg13g2_decap_8 FILLER_74_3250 ();
 sg13g2_decap_8 FILLER_74_3257 ();
 sg13g2_decap_8 FILLER_74_3264 ();
 sg13g2_decap_8 FILLER_74_3271 ();
 sg13g2_decap_8 FILLER_74_3278 ();
 sg13g2_decap_8 FILLER_74_3285 ();
 sg13g2_decap_8 FILLER_74_3292 ();
 sg13g2_decap_8 FILLER_74_3299 ();
 sg13g2_decap_8 FILLER_74_3306 ();
 sg13g2_decap_8 FILLER_74_3313 ();
 sg13g2_decap_8 FILLER_74_3320 ();
 sg13g2_decap_8 FILLER_74_3327 ();
 sg13g2_decap_8 FILLER_74_3334 ();
 sg13g2_decap_8 FILLER_74_3341 ();
 sg13g2_decap_8 FILLER_74_3348 ();
 sg13g2_decap_8 FILLER_74_3355 ();
 sg13g2_decap_8 FILLER_74_3362 ();
 sg13g2_decap_8 FILLER_74_3369 ();
 sg13g2_decap_8 FILLER_74_3376 ();
 sg13g2_decap_8 FILLER_74_3383 ();
 sg13g2_decap_8 FILLER_74_3390 ();
 sg13g2_decap_8 FILLER_74_3397 ();
 sg13g2_decap_8 FILLER_74_3404 ();
 sg13g2_decap_8 FILLER_74_3411 ();
 sg13g2_decap_8 FILLER_74_3418 ();
 sg13g2_decap_8 FILLER_74_3425 ();
 sg13g2_decap_8 FILLER_74_3432 ();
 sg13g2_decap_8 FILLER_74_3439 ();
 sg13g2_decap_8 FILLER_74_3446 ();
 sg13g2_decap_8 FILLER_74_3453 ();
 sg13g2_decap_8 FILLER_74_3460 ();
 sg13g2_decap_8 FILLER_74_3467 ();
 sg13g2_decap_8 FILLER_74_3474 ();
 sg13g2_decap_8 FILLER_74_3481 ();
 sg13g2_decap_8 FILLER_74_3488 ();
 sg13g2_decap_8 FILLER_74_3495 ();
 sg13g2_decap_8 FILLER_74_3502 ();
 sg13g2_decap_8 FILLER_74_3509 ();
 sg13g2_decap_8 FILLER_74_3516 ();
 sg13g2_decap_8 FILLER_74_3523 ();
 sg13g2_decap_8 FILLER_74_3530 ();
 sg13g2_decap_8 FILLER_74_3537 ();
 sg13g2_decap_8 FILLER_74_3544 ();
 sg13g2_decap_8 FILLER_74_3551 ();
 sg13g2_decap_8 FILLER_74_3558 ();
 sg13g2_decap_8 FILLER_74_3565 ();
 sg13g2_decap_8 FILLER_74_3572 ();
 sg13g2_fill_1 FILLER_74_3579 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_4 FILLER_75_98 ();
 sg13g2_fill_1 FILLER_75_102 ();
 sg13g2_fill_2 FILLER_75_107 ();
 sg13g2_fill_1 FILLER_75_109 ();
 sg13g2_fill_2 FILLER_75_171 ();
 sg13g2_fill_1 FILLER_75_173 ();
 sg13g2_fill_2 FILLER_75_188 ();
 sg13g2_fill_1 FILLER_75_195 ();
 sg13g2_fill_2 FILLER_75_206 ();
 sg13g2_fill_2 FILLER_75_231 ();
 sg13g2_fill_1 FILLER_75_233 ();
 sg13g2_fill_2 FILLER_75_280 ();
 sg13g2_fill_1 FILLER_75_282 ();
 sg13g2_fill_1 FILLER_75_318 ();
 sg13g2_fill_2 FILLER_75_343 ();
 sg13g2_fill_1 FILLER_75_345 ();
 sg13g2_fill_1 FILLER_75_356 ();
 sg13g2_fill_2 FILLER_75_362 ();
 sg13g2_decap_8 FILLER_75_377 ();
 sg13g2_decap_8 FILLER_75_384 ();
 sg13g2_fill_1 FILLER_75_395 ();
 sg13g2_fill_2 FILLER_75_413 ();
 sg13g2_fill_2 FILLER_75_453 ();
 sg13g2_fill_1 FILLER_75_464 ();
 sg13g2_fill_2 FILLER_75_491 ();
 sg13g2_fill_2 FILLER_75_499 ();
 sg13g2_fill_1 FILLER_75_522 ();
 sg13g2_fill_2 FILLER_75_538 ();
 sg13g2_fill_1 FILLER_75_540 ();
 sg13g2_fill_1 FILLER_75_561 ();
 sg13g2_fill_2 FILLER_75_614 ();
 sg13g2_fill_2 FILLER_75_636 ();
 sg13g2_fill_2 FILLER_75_643 ();
 sg13g2_fill_1 FILLER_75_645 ();
 sg13g2_fill_2 FILLER_75_653 ();
 sg13g2_fill_1 FILLER_75_655 ();
 sg13g2_fill_2 FILLER_75_673 ();
 sg13g2_fill_1 FILLER_75_675 ();
 sg13g2_fill_1 FILLER_75_690 ();
 sg13g2_fill_1 FILLER_75_696 ();
 sg13g2_fill_1 FILLER_75_766 ();
 sg13g2_decap_8 FILLER_75_793 ();
 sg13g2_fill_1 FILLER_75_800 ();
 sg13g2_fill_1 FILLER_75_815 ();
 sg13g2_decap_4 FILLER_75_834 ();
 sg13g2_fill_1 FILLER_75_838 ();
 sg13g2_fill_1 FILLER_75_869 ();
 sg13g2_decap_4 FILLER_75_899 ();
 sg13g2_decap_8 FILLER_75_930 ();
 sg13g2_fill_2 FILLER_75_937 ();
 sg13g2_fill_2 FILLER_75_967 ();
 sg13g2_fill_1 FILLER_75_969 ();
 sg13g2_fill_1 FILLER_75_984 ();
 sg13g2_fill_1 FILLER_75_1046 ();
 sg13g2_decap_8 FILLER_75_1073 ();
 sg13g2_decap_8 FILLER_75_1080 ();
 sg13g2_fill_2 FILLER_75_1099 ();
 sg13g2_fill_1 FILLER_75_1110 ();
 sg13g2_decap_8 FILLER_75_1119 ();
 sg13g2_fill_2 FILLER_75_1126 ();
 sg13g2_fill_1 FILLER_75_1128 ();
 sg13g2_fill_1 FILLER_75_1175 ();
 sg13g2_decap_4 FILLER_75_1214 ();
 sg13g2_fill_2 FILLER_75_1229 ();
 sg13g2_fill_1 FILLER_75_1253 ();
 sg13g2_fill_2 FILLER_75_1263 ();
 sg13g2_decap_8 FILLER_75_1269 ();
 sg13g2_decap_4 FILLER_75_1276 ();
 sg13g2_fill_1 FILLER_75_1280 ();
 sg13g2_fill_1 FILLER_75_1330 ();
 sg13g2_fill_1 FILLER_75_1337 ();
 sg13g2_fill_1 FILLER_75_1384 ();
 sg13g2_fill_2 FILLER_75_1400 ();
 sg13g2_decap_8 FILLER_75_1408 ();
 sg13g2_decap_8 FILLER_75_1415 ();
 sg13g2_decap_4 FILLER_75_1422 ();
 sg13g2_decap_8 FILLER_75_1434 ();
 sg13g2_fill_1 FILLER_75_1441 ();
 sg13g2_fill_1 FILLER_75_1448 ();
 sg13g2_decap_8 FILLER_75_1468 ();
 sg13g2_decap_8 FILLER_75_1480 ();
 sg13g2_decap_4 FILLER_75_1487 ();
 sg13g2_fill_1 FILLER_75_1495 ();
 sg13g2_decap_4 FILLER_75_1501 ();
 sg13g2_decap_8 FILLER_75_1529 ();
 sg13g2_fill_2 FILLER_75_1536 ();
 sg13g2_decap_8 FILLER_75_1542 ();
 sg13g2_decap_4 FILLER_75_1549 ();
 sg13g2_fill_1 FILLER_75_1553 ();
 sg13g2_decap_4 FILLER_75_1560 ();
 sg13g2_fill_2 FILLER_75_1564 ();
 sg13g2_decap_8 FILLER_75_1576 ();
 sg13g2_fill_1 FILLER_75_1583 ();
 sg13g2_fill_2 FILLER_75_1630 ();
 sg13g2_fill_1 FILLER_75_1632 ();
 sg13g2_decap_8 FILLER_75_1649 ();
 sg13g2_fill_1 FILLER_75_1656 ();
 sg13g2_decap_8 FILLER_75_1675 ();
 sg13g2_decap_4 FILLER_75_1682 ();
 sg13g2_fill_1 FILLER_75_1686 ();
 sg13g2_fill_1 FILLER_75_1692 ();
 sg13g2_decap_8 FILLER_75_1728 ();
 sg13g2_decap_8 FILLER_75_1735 ();
 sg13g2_decap_4 FILLER_75_1742 ();
 sg13g2_fill_2 FILLER_75_1750 ();
 sg13g2_fill_1 FILLER_75_1752 ();
 sg13g2_decap_8 FILLER_75_1779 ();
 sg13g2_fill_1 FILLER_75_1786 ();
 sg13g2_fill_2 FILLER_75_1791 ();
 sg13g2_decap_4 FILLER_75_1806 ();
 sg13g2_fill_2 FILLER_75_1906 ();
 sg13g2_decap_8 FILLER_75_1934 ();
 sg13g2_decap_4 FILLER_75_2006 ();
 sg13g2_fill_2 FILLER_75_2015 ();
 sg13g2_fill_1 FILLER_75_2017 ();
 sg13g2_fill_2 FILLER_75_2033 ();
 sg13g2_decap_4 FILLER_75_2087 ();
 sg13g2_fill_2 FILLER_75_2091 ();
 sg13g2_fill_2 FILLER_75_2161 ();
 sg13g2_fill_1 FILLER_75_2163 ();
 sg13g2_fill_2 FILLER_75_2174 ();
 sg13g2_fill_1 FILLER_75_2211 ();
 sg13g2_decap_4 FILLER_75_2217 ();
 sg13g2_decap_4 FILLER_75_2234 ();
 sg13g2_fill_1 FILLER_75_2238 ();
 sg13g2_decap_8 FILLER_75_2252 ();
 sg13g2_fill_1 FILLER_75_2277 ();
 sg13g2_decap_8 FILLER_75_2291 ();
 sg13g2_fill_2 FILLER_75_2306 ();
 sg13g2_decap_8 FILLER_75_2317 ();
 sg13g2_decap_4 FILLER_75_2324 ();
 sg13g2_fill_1 FILLER_75_2328 ();
 sg13g2_fill_1 FILLER_75_2334 ();
 sg13g2_decap_8 FILLER_75_2339 ();
 sg13g2_fill_1 FILLER_75_2346 ();
 sg13g2_fill_1 FILLER_75_2352 ();
 sg13g2_decap_4 FILLER_75_2366 ();
 sg13g2_fill_2 FILLER_75_2396 ();
 sg13g2_fill_1 FILLER_75_2398 ();
 sg13g2_decap_4 FILLER_75_2404 ();
 sg13g2_fill_1 FILLER_75_2408 ();
 sg13g2_decap_8 FILLER_75_2417 ();
 sg13g2_decap_4 FILLER_75_2428 ();
 sg13g2_fill_1 FILLER_75_2432 ();
 sg13g2_decap_4 FILLER_75_2439 ();
 sg13g2_fill_1 FILLER_75_2443 ();
 sg13g2_fill_2 FILLER_75_2453 ();
 sg13g2_decap_8 FILLER_75_2481 ();
 sg13g2_fill_1 FILLER_75_2488 ();
 sg13g2_decap_4 FILLER_75_2493 ();
 sg13g2_fill_2 FILLER_75_2501 ();
 sg13g2_fill_1 FILLER_75_2503 ();
 sg13g2_decap_8 FILLER_75_2515 ();
 sg13g2_fill_2 FILLER_75_2558 ();
 sg13g2_fill_1 FILLER_75_2560 ();
 sg13g2_fill_2 FILLER_75_2565 ();
 sg13g2_fill_1 FILLER_75_2567 ();
 sg13g2_decap_8 FILLER_75_2591 ();
 sg13g2_decap_4 FILLER_75_2598 ();
 sg13g2_fill_2 FILLER_75_2602 ();
 sg13g2_fill_1 FILLER_75_2613 ();
 sg13g2_fill_2 FILLER_75_2622 ();
 sg13g2_fill_1 FILLER_75_2672 ();
 sg13g2_decap_4 FILLER_75_2684 ();
 sg13g2_fill_2 FILLER_75_2688 ();
 sg13g2_fill_2 FILLER_75_2703 ();
 sg13g2_decap_4 FILLER_75_2746 ();
 sg13g2_fill_2 FILLER_75_2750 ();
 sg13g2_decap_4 FILLER_75_2757 ();
 sg13g2_fill_2 FILLER_75_2784 ();
 sg13g2_fill_1 FILLER_75_2786 ();
 sg13g2_decap_4 FILLER_75_2809 ();
 sg13g2_fill_1 FILLER_75_2813 ();
 sg13g2_fill_1 FILLER_75_2819 ();
 sg13g2_fill_2 FILLER_75_2838 ();
 sg13g2_fill_1 FILLER_75_2840 ();
 sg13g2_decap_8 FILLER_75_2858 ();
 sg13g2_fill_1 FILLER_75_2865 ();
 sg13g2_decap_8 FILLER_75_2893 ();
 sg13g2_fill_2 FILLER_75_2900 ();
 sg13g2_decap_8 FILLER_75_2932 ();
 sg13g2_decap_8 FILLER_75_2939 ();
 sg13g2_decap_8 FILLER_75_2946 ();
 sg13g2_decap_8 FILLER_75_2953 ();
 sg13g2_decap_8 FILLER_75_2960 ();
 sg13g2_decap_8 FILLER_75_2967 ();
 sg13g2_decap_8 FILLER_75_2974 ();
 sg13g2_decap_8 FILLER_75_2981 ();
 sg13g2_decap_8 FILLER_75_2988 ();
 sg13g2_decap_8 FILLER_75_2995 ();
 sg13g2_decap_8 FILLER_75_3002 ();
 sg13g2_decap_8 FILLER_75_3009 ();
 sg13g2_decap_8 FILLER_75_3016 ();
 sg13g2_decap_8 FILLER_75_3023 ();
 sg13g2_decap_8 FILLER_75_3030 ();
 sg13g2_decap_8 FILLER_75_3037 ();
 sg13g2_decap_8 FILLER_75_3044 ();
 sg13g2_decap_8 FILLER_75_3051 ();
 sg13g2_decap_8 FILLER_75_3058 ();
 sg13g2_decap_8 FILLER_75_3065 ();
 sg13g2_decap_8 FILLER_75_3072 ();
 sg13g2_decap_8 FILLER_75_3079 ();
 sg13g2_decap_8 FILLER_75_3086 ();
 sg13g2_decap_8 FILLER_75_3093 ();
 sg13g2_decap_8 FILLER_75_3100 ();
 sg13g2_decap_8 FILLER_75_3107 ();
 sg13g2_decap_8 FILLER_75_3114 ();
 sg13g2_decap_8 FILLER_75_3121 ();
 sg13g2_decap_8 FILLER_75_3128 ();
 sg13g2_decap_8 FILLER_75_3135 ();
 sg13g2_decap_8 FILLER_75_3142 ();
 sg13g2_decap_8 FILLER_75_3149 ();
 sg13g2_decap_8 FILLER_75_3156 ();
 sg13g2_decap_8 FILLER_75_3163 ();
 sg13g2_decap_8 FILLER_75_3170 ();
 sg13g2_decap_8 FILLER_75_3177 ();
 sg13g2_decap_8 FILLER_75_3184 ();
 sg13g2_decap_8 FILLER_75_3191 ();
 sg13g2_decap_8 FILLER_75_3198 ();
 sg13g2_decap_8 FILLER_75_3205 ();
 sg13g2_decap_8 FILLER_75_3212 ();
 sg13g2_decap_8 FILLER_75_3219 ();
 sg13g2_decap_8 FILLER_75_3226 ();
 sg13g2_decap_8 FILLER_75_3233 ();
 sg13g2_decap_8 FILLER_75_3240 ();
 sg13g2_decap_8 FILLER_75_3247 ();
 sg13g2_decap_8 FILLER_75_3254 ();
 sg13g2_decap_8 FILLER_75_3261 ();
 sg13g2_decap_8 FILLER_75_3268 ();
 sg13g2_decap_8 FILLER_75_3275 ();
 sg13g2_decap_8 FILLER_75_3282 ();
 sg13g2_decap_8 FILLER_75_3289 ();
 sg13g2_decap_8 FILLER_75_3296 ();
 sg13g2_decap_8 FILLER_75_3303 ();
 sg13g2_decap_8 FILLER_75_3310 ();
 sg13g2_decap_8 FILLER_75_3317 ();
 sg13g2_decap_8 FILLER_75_3324 ();
 sg13g2_decap_8 FILLER_75_3331 ();
 sg13g2_decap_8 FILLER_75_3338 ();
 sg13g2_decap_8 FILLER_75_3345 ();
 sg13g2_decap_8 FILLER_75_3352 ();
 sg13g2_decap_8 FILLER_75_3359 ();
 sg13g2_decap_8 FILLER_75_3366 ();
 sg13g2_decap_8 FILLER_75_3373 ();
 sg13g2_decap_8 FILLER_75_3380 ();
 sg13g2_decap_8 FILLER_75_3387 ();
 sg13g2_decap_8 FILLER_75_3394 ();
 sg13g2_decap_8 FILLER_75_3401 ();
 sg13g2_decap_8 FILLER_75_3408 ();
 sg13g2_decap_8 FILLER_75_3415 ();
 sg13g2_decap_8 FILLER_75_3422 ();
 sg13g2_decap_8 FILLER_75_3429 ();
 sg13g2_decap_8 FILLER_75_3436 ();
 sg13g2_decap_8 FILLER_75_3443 ();
 sg13g2_decap_8 FILLER_75_3450 ();
 sg13g2_decap_8 FILLER_75_3457 ();
 sg13g2_decap_8 FILLER_75_3464 ();
 sg13g2_decap_8 FILLER_75_3471 ();
 sg13g2_decap_8 FILLER_75_3478 ();
 sg13g2_decap_8 FILLER_75_3485 ();
 sg13g2_decap_8 FILLER_75_3492 ();
 sg13g2_decap_8 FILLER_75_3499 ();
 sg13g2_decap_8 FILLER_75_3506 ();
 sg13g2_decap_8 FILLER_75_3513 ();
 sg13g2_decap_8 FILLER_75_3520 ();
 sg13g2_decap_8 FILLER_75_3527 ();
 sg13g2_decap_8 FILLER_75_3534 ();
 sg13g2_decap_8 FILLER_75_3541 ();
 sg13g2_decap_8 FILLER_75_3548 ();
 sg13g2_decap_8 FILLER_75_3555 ();
 sg13g2_decap_8 FILLER_75_3562 ();
 sg13g2_decap_8 FILLER_75_3569 ();
 sg13g2_decap_4 FILLER_75_3576 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_fill_1 FILLER_76_119 ();
 sg13g2_fill_1 FILLER_76_133 ();
 sg13g2_decap_4 FILLER_76_143 ();
 sg13g2_fill_1 FILLER_76_147 ();
 sg13g2_decap_4 FILLER_76_198 ();
 sg13g2_fill_2 FILLER_76_246 ();
 sg13g2_fill_1 FILLER_76_248 ();
 sg13g2_fill_1 FILLER_76_310 ();
 sg13g2_fill_2 FILLER_76_316 ();
 sg13g2_fill_1 FILLER_76_323 ();
 sg13g2_fill_1 FILLER_76_332 ();
 sg13g2_decap_4 FILLER_76_377 ();
 sg13g2_fill_2 FILLER_76_381 ();
 sg13g2_decap_4 FILLER_76_401 ();
 sg13g2_fill_2 FILLER_76_418 ();
 sg13g2_fill_1 FILLER_76_420 ();
 sg13g2_fill_1 FILLER_76_426 ();
 sg13g2_fill_1 FILLER_76_436 ();
 sg13g2_fill_2 FILLER_76_446 ();
 sg13g2_fill_2 FILLER_76_489 ();
 sg13g2_fill_1 FILLER_76_491 ();
 sg13g2_fill_2 FILLER_76_535 ();
 sg13g2_fill_2 FILLER_76_542 ();
 sg13g2_fill_1 FILLER_76_550 ();
 sg13g2_fill_2 FILLER_76_569 ();
 sg13g2_fill_2 FILLER_76_597 ();
 sg13g2_decap_8 FILLER_76_603 ();
 sg13g2_fill_2 FILLER_76_610 ();
 sg13g2_fill_1 FILLER_76_612 ();
 sg13g2_decap_4 FILLER_76_639 ();
 sg13g2_fill_2 FILLER_76_643 ();
 sg13g2_fill_2 FILLER_76_656 ();
 sg13g2_fill_1 FILLER_76_658 ();
 sg13g2_fill_2 FILLER_76_692 ();
 sg13g2_decap_4 FILLER_76_703 ();
 sg13g2_fill_2 FILLER_76_707 ();
 sg13g2_fill_2 FILLER_76_745 ();
 sg13g2_fill_2 FILLER_76_753 ();
 sg13g2_fill_2 FILLER_76_764 ();
 sg13g2_fill_1 FILLER_76_766 ();
 sg13g2_fill_2 FILLER_76_784 ();
 sg13g2_fill_2 FILLER_76_803 ();
 sg13g2_fill_1 FILLER_76_805 ();
 sg13g2_fill_2 FILLER_76_815 ();
 sg13g2_fill_1 FILLER_76_817 ();
 sg13g2_fill_2 FILLER_76_834 ();
 sg13g2_fill_1 FILLER_76_843 ();
 sg13g2_fill_2 FILLER_76_870 ();
 sg13g2_fill_1 FILLER_76_872 ();
 sg13g2_fill_2 FILLER_76_917 ();
 sg13g2_fill_1 FILLER_76_919 ();
 sg13g2_decap_8 FILLER_76_966 ();
 sg13g2_fill_2 FILLER_76_973 ();
 sg13g2_fill_2 FILLER_76_1015 ();
 sg13g2_fill_1 FILLER_76_1026 ();
 sg13g2_fill_1 FILLER_76_1037 ();
 sg13g2_fill_1 FILLER_76_1048 ();
 sg13g2_fill_2 FILLER_76_1088 ();
 sg13g2_fill_1 FILLER_76_1090 ();
 sg13g2_decap_4 FILLER_76_1097 ();
 sg13g2_fill_2 FILLER_76_1101 ();
 sg13g2_fill_2 FILLER_76_1169 ();
 sg13g2_fill_2 FILLER_76_1183 ();
 sg13g2_fill_2 FILLER_76_1207 ();
 sg13g2_fill_2 FILLER_76_1222 ();
 sg13g2_fill_1 FILLER_76_1224 ();
 sg13g2_decap_4 FILLER_76_1270 ();
 sg13g2_decap_4 FILLER_76_1280 ();
 sg13g2_fill_2 FILLER_76_1321 ();
 sg13g2_fill_1 FILLER_76_1323 ();
 sg13g2_decap_8 FILLER_76_1337 ();
 sg13g2_fill_2 FILLER_76_1344 ();
 sg13g2_fill_2 FILLER_76_1355 ();
 sg13g2_fill_2 FILLER_76_1372 ();
 sg13g2_fill_2 FILLER_76_1379 ();
 sg13g2_fill_1 FILLER_76_1381 ();
 sg13g2_decap_8 FILLER_76_1390 ();
 sg13g2_fill_2 FILLER_76_1397 ();
 sg13g2_decap_8 FILLER_76_1430 ();
 sg13g2_fill_2 FILLER_76_1437 ();
 sg13g2_fill_1 FILLER_76_1439 ();
 sg13g2_fill_1 FILLER_76_1444 ();
 sg13g2_decap_8 FILLER_76_1451 ();
 sg13g2_decap_8 FILLER_76_1458 ();
 sg13g2_fill_2 FILLER_76_1465 ();
 sg13g2_decap_4 FILLER_76_1478 ();
 sg13g2_fill_1 FILLER_76_1482 ();
 sg13g2_decap_8 FILLER_76_1497 ();
 sg13g2_decap_8 FILLER_76_1504 ();
 sg13g2_decap_4 FILLER_76_1511 ();
 sg13g2_decap_8 FILLER_76_1536 ();
 sg13g2_fill_1 FILLER_76_1543 ();
 sg13g2_decap_4 FILLER_76_1548 ();
 sg13g2_fill_2 FILLER_76_1567 ();
 sg13g2_fill_2 FILLER_76_1609 ();
 sg13g2_fill_1 FILLER_76_1611 ();
 sg13g2_fill_1 FILLER_76_1634 ();
 sg13g2_decap_4 FILLER_76_1647 ();
 sg13g2_fill_2 FILLER_76_1682 ();
 sg13g2_fill_1 FILLER_76_1684 ();
 sg13g2_fill_1 FILLER_76_1693 ();
 sg13g2_decap_8 FILLER_76_1725 ();
 sg13g2_fill_1 FILLER_76_1732 ();
 sg13g2_decap_8 FILLER_76_1737 ();
 sg13g2_decap_8 FILLER_76_1744 ();
 sg13g2_decap_8 FILLER_76_1751 ();
 sg13g2_decap_4 FILLER_76_1758 ();
 sg13g2_fill_2 FILLER_76_1762 ();
 sg13g2_decap_8 FILLER_76_1768 ();
 sg13g2_fill_1 FILLER_76_1775 ();
 sg13g2_fill_2 FILLER_76_1802 ();
 sg13g2_decap_8 FILLER_76_1808 ();
 sg13g2_decap_4 FILLER_76_1815 ();
 sg13g2_fill_2 FILLER_76_1819 ();
 sg13g2_decap_8 FILLER_76_1860 ();
 sg13g2_decap_8 FILLER_76_1867 ();
 sg13g2_decap_4 FILLER_76_1874 ();
 sg13g2_fill_2 FILLER_76_1878 ();
 sg13g2_fill_2 FILLER_76_1884 ();
 sg13g2_decap_8 FILLER_76_1918 ();
 sg13g2_decap_4 FILLER_76_1925 ();
 sg13g2_fill_1 FILLER_76_1929 ();
 sg13g2_decap_8 FILLER_76_1963 ();
 sg13g2_decap_8 FILLER_76_1970 ();
 sg13g2_fill_2 FILLER_76_1977 ();
 sg13g2_fill_2 FILLER_76_2042 ();
 sg13g2_fill_2 FILLER_76_2049 ();
 sg13g2_fill_1 FILLER_76_2051 ();
 sg13g2_fill_2 FILLER_76_2059 ();
 sg13g2_decap_8 FILLER_76_2084 ();
 sg13g2_fill_2 FILLER_76_2091 ();
 sg13g2_fill_2 FILLER_76_2101 ();
 sg13g2_fill_1 FILLER_76_2103 ();
 sg13g2_decap_8 FILLER_76_2108 ();
 sg13g2_decap_4 FILLER_76_2115 ();
 sg13g2_fill_1 FILLER_76_2119 ();
 sg13g2_fill_2 FILLER_76_2156 ();
 sg13g2_fill_2 FILLER_76_2199 ();
 sg13g2_fill_1 FILLER_76_2201 ();
 sg13g2_decap_8 FILLER_76_2211 ();
 sg13g2_decap_8 FILLER_76_2226 ();
 sg13g2_decap_8 FILLER_76_2255 ();
 sg13g2_decap_8 FILLER_76_2267 ();
 sg13g2_fill_2 FILLER_76_2279 ();
 sg13g2_decap_4 FILLER_76_2301 ();
 sg13g2_decap_4 FILLER_76_2311 ();
 sg13g2_fill_2 FILLER_76_2338 ();
 sg13g2_fill_1 FILLER_76_2340 ();
 sg13g2_fill_2 FILLER_76_2346 ();
 sg13g2_fill_1 FILLER_76_2348 ();
 sg13g2_fill_2 FILLER_76_2371 ();
 sg13g2_fill_2 FILLER_76_2422 ();
 sg13g2_fill_1 FILLER_76_2424 ();
 sg13g2_fill_1 FILLER_76_2448 ();
 sg13g2_fill_1 FILLER_76_2452 ();
 sg13g2_fill_1 FILLER_76_2462 ();
 sg13g2_fill_1 FILLER_76_2467 ();
 sg13g2_fill_2 FILLER_76_2494 ();
 sg13g2_decap_8 FILLER_76_2517 ();
 sg13g2_decap_8 FILLER_76_2524 ();
 sg13g2_decap_4 FILLER_76_2531 ();
 sg13g2_fill_1 FILLER_76_2535 ();
 sg13g2_decap_4 FILLER_76_2540 ();
 sg13g2_fill_2 FILLER_76_2563 ();
 sg13g2_fill_1 FILLER_76_2565 ();
 sg13g2_decap_4 FILLER_76_2571 ();
 sg13g2_decap_8 FILLER_76_2580 ();
 sg13g2_decap_8 FILLER_76_2596 ();
 sg13g2_decap_4 FILLER_76_2603 ();
 sg13g2_decap_8 FILLER_76_2626 ();
 sg13g2_decap_4 FILLER_76_2633 ();
 sg13g2_fill_1 FILLER_76_2649 ();
 sg13g2_decap_4 FILLER_76_2659 ();
 sg13g2_fill_1 FILLER_76_2667 ();
 sg13g2_fill_1 FILLER_76_2672 ();
 sg13g2_decap_4 FILLER_76_2695 ();
 sg13g2_fill_1 FILLER_76_2699 ();
 sg13g2_decap_8 FILLER_76_2705 ();
 sg13g2_fill_1 FILLER_76_2712 ();
 sg13g2_fill_2 FILLER_76_2750 ();
 sg13g2_fill_1 FILLER_76_2752 ();
 sg13g2_fill_2 FILLER_76_2766 ();
 sg13g2_decap_4 FILLER_76_2776 ();
 sg13g2_fill_2 FILLER_76_2780 ();
 sg13g2_fill_2 FILLER_76_2799 ();
 sg13g2_decap_8 FILLER_76_2809 ();
 sg13g2_decap_8 FILLER_76_2816 ();
 sg13g2_fill_1 FILLER_76_2823 ();
 sg13g2_fill_1 FILLER_76_2842 ();
 sg13g2_decap_8 FILLER_76_2860 ();
 sg13g2_decap_4 FILLER_76_2872 ();
 sg13g2_fill_1 FILLER_76_2876 ();
 sg13g2_decap_8 FILLER_76_2885 ();
 sg13g2_fill_1 FILLER_76_2892 ();
 sg13g2_decap_4 FILLER_76_2904 ();
 sg13g2_fill_2 FILLER_76_2908 ();
 sg13g2_fill_1 FILLER_76_2923 ();
 sg13g2_fill_1 FILLER_76_2929 ();
 sg13g2_decap_8 FILLER_76_2946 ();
 sg13g2_decap_8 FILLER_76_2953 ();
 sg13g2_decap_8 FILLER_76_2960 ();
 sg13g2_decap_8 FILLER_76_2967 ();
 sg13g2_decap_8 FILLER_76_2974 ();
 sg13g2_decap_8 FILLER_76_2981 ();
 sg13g2_decap_8 FILLER_76_2988 ();
 sg13g2_decap_8 FILLER_76_2995 ();
 sg13g2_decap_8 FILLER_76_3002 ();
 sg13g2_decap_8 FILLER_76_3009 ();
 sg13g2_decap_8 FILLER_76_3016 ();
 sg13g2_decap_8 FILLER_76_3023 ();
 sg13g2_decap_8 FILLER_76_3030 ();
 sg13g2_decap_8 FILLER_76_3037 ();
 sg13g2_decap_8 FILLER_76_3044 ();
 sg13g2_decap_8 FILLER_76_3051 ();
 sg13g2_decap_8 FILLER_76_3058 ();
 sg13g2_decap_8 FILLER_76_3065 ();
 sg13g2_decap_8 FILLER_76_3072 ();
 sg13g2_decap_8 FILLER_76_3079 ();
 sg13g2_decap_8 FILLER_76_3086 ();
 sg13g2_decap_8 FILLER_76_3093 ();
 sg13g2_decap_8 FILLER_76_3100 ();
 sg13g2_decap_8 FILLER_76_3107 ();
 sg13g2_decap_8 FILLER_76_3114 ();
 sg13g2_decap_8 FILLER_76_3121 ();
 sg13g2_decap_8 FILLER_76_3128 ();
 sg13g2_decap_8 FILLER_76_3135 ();
 sg13g2_decap_8 FILLER_76_3142 ();
 sg13g2_decap_8 FILLER_76_3149 ();
 sg13g2_decap_8 FILLER_76_3156 ();
 sg13g2_decap_8 FILLER_76_3163 ();
 sg13g2_decap_8 FILLER_76_3170 ();
 sg13g2_decap_8 FILLER_76_3177 ();
 sg13g2_decap_8 FILLER_76_3184 ();
 sg13g2_decap_8 FILLER_76_3191 ();
 sg13g2_decap_8 FILLER_76_3198 ();
 sg13g2_decap_8 FILLER_76_3205 ();
 sg13g2_decap_8 FILLER_76_3212 ();
 sg13g2_decap_8 FILLER_76_3219 ();
 sg13g2_decap_8 FILLER_76_3226 ();
 sg13g2_decap_8 FILLER_76_3233 ();
 sg13g2_decap_8 FILLER_76_3240 ();
 sg13g2_decap_8 FILLER_76_3247 ();
 sg13g2_decap_8 FILLER_76_3254 ();
 sg13g2_decap_8 FILLER_76_3261 ();
 sg13g2_decap_8 FILLER_76_3268 ();
 sg13g2_decap_8 FILLER_76_3275 ();
 sg13g2_decap_8 FILLER_76_3282 ();
 sg13g2_decap_8 FILLER_76_3289 ();
 sg13g2_decap_8 FILLER_76_3296 ();
 sg13g2_decap_8 FILLER_76_3303 ();
 sg13g2_decap_8 FILLER_76_3310 ();
 sg13g2_decap_8 FILLER_76_3317 ();
 sg13g2_decap_8 FILLER_76_3324 ();
 sg13g2_decap_8 FILLER_76_3331 ();
 sg13g2_decap_8 FILLER_76_3338 ();
 sg13g2_decap_8 FILLER_76_3345 ();
 sg13g2_decap_8 FILLER_76_3352 ();
 sg13g2_decap_8 FILLER_76_3359 ();
 sg13g2_decap_8 FILLER_76_3366 ();
 sg13g2_decap_8 FILLER_76_3373 ();
 sg13g2_decap_8 FILLER_76_3380 ();
 sg13g2_decap_8 FILLER_76_3387 ();
 sg13g2_decap_8 FILLER_76_3394 ();
 sg13g2_decap_8 FILLER_76_3401 ();
 sg13g2_decap_8 FILLER_76_3408 ();
 sg13g2_decap_8 FILLER_76_3415 ();
 sg13g2_decap_8 FILLER_76_3422 ();
 sg13g2_decap_8 FILLER_76_3429 ();
 sg13g2_decap_8 FILLER_76_3436 ();
 sg13g2_decap_8 FILLER_76_3443 ();
 sg13g2_decap_8 FILLER_76_3450 ();
 sg13g2_decap_8 FILLER_76_3457 ();
 sg13g2_decap_8 FILLER_76_3464 ();
 sg13g2_decap_8 FILLER_76_3471 ();
 sg13g2_decap_8 FILLER_76_3478 ();
 sg13g2_decap_8 FILLER_76_3485 ();
 sg13g2_decap_8 FILLER_76_3492 ();
 sg13g2_decap_8 FILLER_76_3499 ();
 sg13g2_decap_8 FILLER_76_3506 ();
 sg13g2_decap_8 FILLER_76_3513 ();
 sg13g2_decap_8 FILLER_76_3520 ();
 sg13g2_decap_8 FILLER_76_3527 ();
 sg13g2_decap_8 FILLER_76_3534 ();
 sg13g2_decap_8 FILLER_76_3541 ();
 sg13g2_decap_8 FILLER_76_3548 ();
 sg13g2_decap_8 FILLER_76_3555 ();
 sg13g2_decap_8 FILLER_76_3562 ();
 sg13g2_decap_8 FILLER_76_3569 ();
 sg13g2_decap_4 FILLER_76_3576 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_4 FILLER_77_126 ();
 sg13g2_fill_1 FILLER_77_130 ();
 sg13g2_decap_8 FILLER_77_134 ();
 sg13g2_fill_1 FILLER_77_141 ();
 sg13g2_fill_2 FILLER_77_234 ();
 sg13g2_fill_2 FILLER_77_253 ();
 sg13g2_fill_2 FILLER_77_269 ();
 sg13g2_fill_2 FILLER_77_281 ();
 sg13g2_fill_1 FILLER_77_333 ();
 sg13g2_decap_4 FILLER_77_352 ();
 sg13g2_fill_1 FILLER_77_356 ();
 sg13g2_decap_4 FILLER_77_436 ();
 sg13g2_fill_2 FILLER_77_440 ();
 sg13g2_decap_8 FILLER_77_451 ();
 sg13g2_fill_2 FILLER_77_458 ();
 sg13g2_fill_2 FILLER_77_485 ();
 sg13g2_fill_1 FILLER_77_487 ();
 sg13g2_fill_2 FILLER_77_528 ();
 sg13g2_fill_1 FILLER_77_544 ();
 sg13g2_fill_2 FILLER_77_585 ();
 sg13g2_fill_1 FILLER_77_587 ();
 sg13g2_decap_8 FILLER_77_627 ();
 sg13g2_decap_8 FILLER_77_634 ();
 sg13g2_fill_2 FILLER_77_641 ();
 sg13g2_fill_1 FILLER_77_651 ();
 sg13g2_decap_4 FILLER_77_670 ();
 sg13g2_fill_1 FILLER_77_674 ();
 sg13g2_fill_1 FILLER_77_727 ();
 sg13g2_fill_1 FILLER_77_731 ();
 sg13g2_fill_1 FILLER_77_892 ();
 sg13g2_fill_1 FILLER_77_920 ();
 sg13g2_fill_2 FILLER_77_951 ();
 sg13g2_fill_1 FILLER_77_968 ();
 sg13g2_fill_1 FILLER_77_1027 ();
 sg13g2_fill_1 FILLER_77_1080 ();
 sg13g2_fill_1 FILLER_77_1165 ();
 sg13g2_fill_1 FILLER_77_1197 ();
 sg13g2_decap_4 FILLER_77_1276 ();
 sg13g2_decap_4 FILLER_77_1388 ();
 sg13g2_decap_4 FILLER_77_1459 ();
 sg13g2_fill_1 FILLER_77_1463 ();
 sg13g2_fill_2 FILLER_77_1504 ();
 sg13g2_fill_1 FILLER_77_1506 ();
 sg13g2_decap_4 FILLER_77_1591 ();
 sg13g2_fill_2 FILLER_77_1605 ();
 sg13g2_fill_1 FILLER_77_1607 ();
 sg13g2_fill_1 FILLER_77_1629 ();
 sg13g2_fill_2 FILLER_77_1638 ();
 sg13g2_fill_1 FILLER_77_1640 ();
 sg13g2_decap_4 FILLER_77_1646 ();
 sg13g2_decap_4 FILLER_77_1660 ();
 sg13g2_fill_1 FILLER_77_1668 ();
 sg13g2_decap_4 FILLER_77_1678 ();
 sg13g2_fill_2 FILLER_77_1687 ();
 sg13g2_fill_1 FILLER_77_1689 ();
 sg13g2_fill_2 FILLER_77_1719 ();
 sg13g2_fill_1 FILLER_77_1721 ();
 sg13g2_decap_8 FILLER_77_1748 ();
 sg13g2_decap_8 FILLER_77_1755 ();
 sg13g2_decap_8 FILLER_77_1762 ();
 sg13g2_decap_8 FILLER_77_1769 ();
 sg13g2_decap_8 FILLER_77_1776 ();
 sg13g2_decap_8 FILLER_77_1783 ();
 sg13g2_decap_4 FILLER_77_1790 ();
 sg13g2_decap_8 FILLER_77_1820 ();
 sg13g2_decap_8 FILLER_77_1827 ();
 sg13g2_fill_2 FILLER_77_1834 ();
 sg13g2_decap_8 FILLER_77_1844 ();
 sg13g2_decap_8 FILLER_77_1851 ();
 sg13g2_decap_8 FILLER_77_1858 ();
 sg13g2_decap_8 FILLER_77_1865 ();
 sg13g2_decap_8 FILLER_77_1872 ();
 sg13g2_decap_8 FILLER_77_1879 ();
 sg13g2_decap_8 FILLER_77_1886 ();
 sg13g2_decap_8 FILLER_77_1893 ();
 sg13g2_fill_2 FILLER_77_1900 ();
 sg13g2_fill_1 FILLER_77_1902 ();
 sg13g2_decap_8 FILLER_77_1907 ();
 sg13g2_decap_4 FILLER_77_1914 ();
 sg13g2_fill_1 FILLER_77_1918 ();
 sg13g2_decap_8 FILLER_77_1923 ();
 sg13g2_decap_8 FILLER_77_1930 ();
 sg13g2_decap_4 FILLER_77_1937 ();
 sg13g2_fill_2 FILLER_77_1941 ();
 sg13g2_decap_8 FILLER_77_1947 ();
 sg13g2_decap_8 FILLER_77_1954 ();
 sg13g2_decap_8 FILLER_77_1961 ();
 sg13g2_decap_8 FILLER_77_1968 ();
 sg13g2_decap_8 FILLER_77_1975 ();
 sg13g2_decap_8 FILLER_77_1986 ();
 sg13g2_fill_1 FILLER_77_1993 ();
 sg13g2_decap_8 FILLER_77_1998 ();
 sg13g2_fill_2 FILLER_77_2005 ();
 sg13g2_fill_1 FILLER_77_2007 ();
 sg13g2_decap_8 FILLER_77_2033 ();
 sg13g2_fill_2 FILLER_77_2066 ();
 sg13g2_fill_2 FILLER_77_2094 ();
 sg13g2_fill_2 FILLER_77_2122 ();
 sg13g2_fill_1 FILLER_77_2124 ();
 sg13g2_fill_1 FILLER_77_2147 ();
 sg13g2_decap_4 FILLER_77_2176 ();
 sg13g2_decap_8 FILLER_77_2223 ();
 sg13g2_fill_1 FILLER_77_2230 ();
 sg13g2_fill_1 FILLER_77_2246 ();
 sg13g2_decap_8 FILLER_77_2267 ();
 sg13g2_decap_8 FILLER_77_2274 ();
 sg13g2_decap_4 FILLER_77_2289 ();
 sg13g2_fill_1 FILLER_77_2293 ();
 sg13g2_fill_2 FILLER_77_2302 ();
 sg13g2_fill_1 FILLER_77_2304 ();
 sg13g2_decap_4 FILLER_77_2321 ();
 sg13g2_fill_2 FILLER_77_2335 ();
 sg13g2_fill_1 FILLER_77_2337 ();
 sg13g2_fill_1 FILLER_77_2347 ();
 sg13g2_decap_8 FILLER_77_2371 ();
 sg13g2_decap_8 FILLER_77_2378 ();
 sg13g2_fill_2 FILLER_77_2385 ();
 sg13g2_fill_1 FILLER_77_2398 ();
 sg13g2_decap_4 FILLER_77_2411 ();
 sg13g2_fill_1 FILLER_77_2424 ();
 sg13g2_fill_2 FILLER_77_2430 ();
 sg13g2_fill_1 FILLER_77_2432 ();
 sg13g2_decap_8 FILLER_77_2438 ();
 sg13g2_fill_1 FILLER_77_2445 ();
 sg13g2_decap_4 FILLER_77_2473 ();
 sg13g2_fill_2 FILLER_77_2477 ();
 sg13g2_decap_8 FILLER_77_2483 ();
 sg13g2_decap_8 FILLER_77_2490 ();
 sg13g2_decap_4 FILLER_77_2497 ();
 sg13g2_fill_2 FILLER_77_2573 ();
 sg13g2_fill_1 FILLER_77_2575 ();
 sg13g2_fill_1 FILLER_77_2594 ();
 sg13g2_fill_2 FILLER_77_2605 ();
 sg13g2_fill_1 FILLER_77_2607 ();
 sg13g2_fill_1 FILLER_77_2618 ();
 sg13g2_decap_8 FILLER_77_2630 ();
 sg13g2_decap_4 FILLER_77_2637 ();
 sg13g2_fill_1 FILLER_77_2650 ();
 sg13g2_decap_8 FILLER_77_2667 ();
 sg13g2_fill_1 FILLER_77_2674 ();
 sg13g2_fill_2 FILLER_77_2687 ();
 sg13g2_fill_1 FILLER_77_2694 ();
 sg13g2_decap_4 FILLER_77_2700 ();
 sg13g2_decap_8 FILLER_77_2716 ();
 sg13g2_fill_1 FILLER_77_2723 ();
 sg13g2_decap_8 FILLER_77_2728 ();
 sg13g2_decap_8 FILLER_77_2740 ();
 sg13g2_fill_1 FILLER_77_2747 ();
 sg13g2_fill_1 FILLER_77_2809 ();
 sg13g2_decap_8 FILLER_77_2824 ();
 sg13g2_fill_2 FILLER_77_2831 ();
 sg13g2_fill_1 FILLER_77_2843 ();
 sg13g2_fill_1 FILLER_77_2861 ();
 sg13g2_fill_1 FILLER_77_2867 ();
 sg13g2_decap_4 FILLER_77_2878 ();
 sg13g2_fill_2 FILLER_77_2882 ();
 sg13g2_fill_2 FILLER_77_2902 ();
 sg13g2_decap_8 FILLER_77_2930 ();
 sg13g2_decap_8 FILLER_77_2937 ();
 sg13g2_decap_8 FILLER_77_2944 ();
 sg13g2_decap_8 FILLER_77_2951 ();
 sg13g2_decap_8 FILLER_77_2958 ();
 sg13g2_decap_8 FILLER_77_2965 ();
 sg13g2_decap_8 FILLER_77_2972 ();
 sg13g2_decap_8 FILLER_77_2979 ();
 sg13g2_decap_8 FILLER_77_2986 ();
 sg13g2_decap_8 FILLER_77_2993 ();
 sg13g2_decap_8 FILLER_77_3000 ();
 sg13g2_decap_8 FILLER_77_3007 ();
 sg13g2_decap_8 FILLER_77_3014 ();
 sg13g2_decap_8 FILLER_77_3021 ();
 sg13g2_decap_8 FILLER_77_3028 ();
 sg13g2_decap_8 FILLER_77_3035 ();
 sg13g2_decap_8 FILLER_77_3042 ();
 sg13g2_decap_8 FILLER_77_3049 ();
 sg13g2_decap_8 FILLER_77_3056 ();
 sg13g2_decap_8 FILLER_77_3063 ();
 sg13g2_decap_8 FILLER_77_3070 ();
 sg13g2_decap_8 FILLER_77_3077 ();
 sg13g2_decap_8 FILLER_77_3084 ();
 sg13g2_decap_8 FILLER_77_3091 ();
 sg13g2_decap_8 FILLER_77_3098 ();
 sg13g2_decap_8 FILLER_77_3105 ();
 sg13g2_decap_8 FILLER_77_3112 ();
 sg13g2_decap_8 FILLER_77_3119 ();
 sg13g2_decap_8 FILLER_77_3126 ();
 sg13g2_decap_8 FILLER_77_3133 ();
 sg13g2_decap_8 FILLER_77_3140 ();
 sg13g2_decap_8 FILLER_77_3147 ();
 sg13g2_decap_8 FILLER_77_3154 ();
 sg13g2_decap_8 FILLER_77_3161 ();
 sg13g2_decap_8 FILLER_77_3168 ();
 sg13g2_decap_8 FILLER_77_3175 ();
 sg13g2_decap_8 FILLER_77_3182 ();
 sg13g2_decap_8 FILLER_77_3189 ();
 sg13g2_decap_8 FILLER_77_3196 ();
 sg13g2_decap_8 FILLER_77_3203 ();
 sg13g2_decap_8 FILLER_77_3210 ();
 sg13g2_decap_8 FILLER_77_3217 ();
 sg13g2_decap_8 FILLER_77_3224 ();
 sg13g2_decap_8 FILLER_77_3231 ();
 sg13g2_decap_8 FILLER_77_3238 ();
 sg13g2_decap_8 FILLER_77_3245 ();
 sg13g2_decap_8 FILLER_77_3252 ();
 sg13g2_decap_8 FILLER_77_3259 ();
 sg13g2_decap_8 FILLER_77_3266 ();
 sg13g2_decap_8 FILLER_77_3273 ();
 sg13g2_decap_8 FILLER_77_3280 ();
 sg13g2_decap_8 FILLER_77_3287 ();
 sg13g2_decap_8 FILLER_77_3294 ();
 sg13g2_decap_8 FILLER_77_3301 ();
 sg13g2_decap_8 FILLER_77_3308 ();
 sg13g2_decap_8 FILLER_77_3315 ();
 sg13g2_decap_8 FILLER_77_3322 ();
 sg13g2_decap_8 FILLER_77_3329 ();
 sg13g2_decap_8 FILLER_77_3336 ();
 sg13g2_decap_8 FILLER_77_3343 ();
 sg13g2_decap_8 FILLER_77_3350 ();
 sg13g2_decap_8 FILLER_77_3357 ();
 sg13g2_decap_8 FILLER_77_3364 ();
 sg13g2_decap_8 FILLER_77_3371 ();
 sg13g2_decap_8 FILLER_77_3378 ();
 sg13g2_decap_8 FILLER_77_3385 ();
 sg13g2_decap_8 FILLER_77_3392 ();
 sg13g2_decap_8 FILLER_77_3399 ();
 sg13g2_decap_8 FILLER_77_3406 ();
 sg13g2_decap_8 FILLER_77_3413 ();
 sg13g2_decap_8 FILLER_77_3420 ();
 sg13g2_decap_8 FILLER_77_3427 ();
 sg13g2_decap_8 FILLER_77_3434 ();
 sg13g2_decap_8 FILLER_77_3441 ();
 sg13g2_decap_8 FILLER_77_3448 ();
 sg13g2_decap_8 FILLER_77_3455 ();
 sg13g2_decap_8 FILLER_77_3462 ();
 sg13g2_decap_8 FILLER_77_3469 ();
 sg13g2_decap_8 FILLER_77_3476 ();
 sg13g2_decap_8 FILLER_77_3483 ();
 sg13g2_decap_8 FILLER_77_3490 ();
 sg13g2_decap_8 FILLER_77_3497 ();
 sg13g2_decap_8 FILLER_77_3504 ();
 sg13g2_decap_8 FILLER_77_3511 ();
 sg13g2_decap_8 FILLER_77_3518 ();
 sg13g2_decap_8 FILLER_77_3525 ();
 sg13g2_decap_8 FILLER_77_3532 ();
 sg13g2_decap_8 FILLER_77_3539 ();
 sg13g2_decap_8 FILLER_77_3546 ();
 sg13g2_decap_8 FILLER_77_3553 ();
 sg13g2_decap_8 FILLER_77_3560 ();
 sg13g2_decap_8 FILLER_77_3567 ();
 sg13g2_decap_4 FILLER_77_3574 ();
 sg13g2_fill_2 FILLER_77_3578 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_8 FILLER_78_140 ();
 sg13g2_decap_8 FILLER_78_147 ();
 sg13g2_fill_2 FILLER_78_154 ();
 sg13g2_fill_1 FILLER_78_156 ();
 sg13g2_decap_8 FILLER_78_161 ();
 sg13g2_fill_1 FILLER_78_168 ();
 sg13g2_decap_8 FILLER_78_186 ();
 sg13g2_fill_1 FILLER_78_193 ();
 sg13g2_decap_4 FILLER_78_199 ();
 sg13g2_fill_2 FILLER_78_208 ();
 sg13g2_decap_8 FILLER_78_214 ();
 sg13g2_decap_8 FILLER_78_221 ();
 sg13g2_fill_1 FILLER_78_228 ();
 sg13g2_fill_1 FILLER_78_271 ();
 sg13g2_fill_1 FILLER_78_315 ();
 sg13g2_fill_2 FILLER_78_347 ();
 sg13g2_fill_1 FILLER_78_395 ();
 sg13g2_decap_8 FILLER_78_425 ();
 sg13g2_fill_2 FILLER_78_432 ();
 sg13g2_fill_1 FILLER_78_460 ();
 sg13g2_fill_1 FILLER_78_482 ();
 sg13g2_fill_2 FILLER_78_509 ();
 sg13g2_fill_1 FILLER_78_580 ();
 sg13g2_fill_2 FILLER_78_607 ();
 sg13g2_fill_2 FILLER_78_623 ();
 sg13g2_decap_4 FILLER_78_634 ();
 sg13g2_fill_2 FILLER_78_673 ();
 sg13g2_fill_1 FILLER_78_675 ();
 sg13g2_fill_2 FILLER_78_711 ();
 sg13g2_fill_1 FILLER_78_737 ();
 sg13g2_fill_2 FILLER_78_763 ();
 sg13g2_fill_1 FILLER_78_774 ();
 sg13g2_decap_4 FILLER_78_820 ();
 sg13g2_decap_4 FILLER_78_850 ();
 sg13g2_fill_1 FILLER_78_854 ();
 sg13g2_fill_1 FILLER_78_864 ();
 sg13g2_fill_1 FILLER_78_878 ();
 sg13g2_fill_2 FILLER_78_902 ();
 sg13g2_fill_1 FILLER_78_904 ();
 sg13g2_fill_1 FILLER_78_928 ();
 sg13g2_fill_2 FILLER_78_944 ();
 sg13g2_fill_1 FILLER_78_946 ();
 sg13g2_fill_2 FILLER_78_964 ();
 sg13g2_fill_2 FILLER_78_987 ();
 sg13g2_fill_1 FILLER_78_989 ();
 sg13g2_decap_4 FILLER_78_1004 ();
 sg13g2_fill_1 FILLER_78_1008 ();
 sg13g2_fill_2 FILLER_78_1054 ();
 sg13g2_decap_4 FILLER_78_1068 ();
 sg13g2_fill_1 FILLER_78_1072 ();
 sg13g2_fill_1 FILLER_78_1105 ();
 sg13g2_fill_2 FILLER_78_1119 ();
 sg13g2_fill_1 FILLER_78_1121 ();
 sg13g2_decap_4 FILLER_78_1178 ();
 sg13g2_fill_2 FILLER_78_1189 ();
 sg13g2_fill_2 FILLER_78_1200 ();
 sg13g2_fill_1 FILLER_78_1202 ();
 sg13g2_fill_2 FILLER_78_1244 ();
 sg13g2_fill_2 FILLER_78_1255 ();
 sg13g2_fill_1 FILLER_78_1257 ();
 sg13g2_fill_1 FILLER_78_1290 ();
 sg13g2_fill_2 FILLER_78_1300 ();
 sg13g2_decap_8 FILLER_78_1322 ();
 sg13g2_decap_8 FILLER_78_1329 ();
 sg13g2_decap_8 FILLER_78_1336 ();
 sg13g2_decap_4 FILLER_78_1347 ();
 sg13g2_fill_2 FILLER_78_1351 ();
 sg13g2_fill_2 FILLER_78_1363 ();
 sg13g2_fill_1 FILLER_78_1389 ();
 sg13g2_fill_2 FILLER_78_1395 ();
 sg13g2_decap_8 FILLER_78_1420 ();
 sg13g2_decap_8 FILLER_78_1427 ();
 sg13g2_fill_1 FILLER_78_1448 ();
 sg13g2_fill_2 FILLER_78_1463 ();
 sg13g2_decap_8 FILLER_78_1475 ();
 sg13g2_fill_2 FILLER_78_1482 ();
 sg13g2_decap_4 FILLER_78_1488 ();
 sg13g2_fill_2 FILLER_78_1492 ();
 sg13g2_fill_2 FILLER_78_1533 ();
 sg13g2_decap_8 FILLER_78_1549 ();
 sg13g2_fill_2 FILLER_78_1556 ();
 sg13g2_fill_1 FILLER_78_1558 ();
 sg13g2_fill_2 FILLER_78_1582 ();
 sg13g2_fill_1 FILLER_78_1584 ();
 sg13g2_fill_2 FILLER_78_1644 ();
 sg13g2_fill_1 FILLER_78_1646 ();
 sg13g2_fill_1 FILLER_78_1652 ();
 sg13g2_fill_2 FILLER_78_1679 ();
 sg13g2_decap_8 FILLER_78_1735 ();
 sg13g2_decap_8 FILLER_78_1742 ();
 sg13g2_decap_8 FILLER_78_1749 ();
 sg13g2_decap_8 FILLER_78_1756 ();
 sg13g2_decap_8 FILLER_78_1763 ();
 sg13g2_decap_8 FILLER_78_1770 ();
 sg13g2_decap_8 FILLER_78_1777 ();
 sg13g2_decap_8 FILLER_78_1784 ();
 sg13g2_decap_8 FILLER_78_1791 ();
 sg13g2_decap_8 FILLER_78_1798 ();
 sg13g2_decap_8 FILLER_78_1805 ();
 sg13g2_decap_8 FILLER_78_1812 ();
 sg13g2_decap_8 FILLER_78_1819 ();
 sg13g2_decap_8 FILLER_78_1826 ();
 sg13g2_decap_8 FILLER_78_1833 ();
 sg13g2_decap_8 FILLER_78_1840 ();
 sg13g2_decap_8 FILLER_78_1847 ();
 sg13g2_decap_8 FILLER_78_1854 ();
 sg13g2_decap_8 FILLER_78_1861 ();
 sg13g2_decap_8 FILLER_78_1868 ();
 sg13g2_decap_8 FILLER_78_1875 ();
 sg13g2_fill_2 FILLER_78_1882 ();
 sg13g2_decap_8 FILLER_78_1892 ();
 sg13g2_decap_8 FILLER_78_1899 ();
 sg13g2_decap_8 FILLER_78_1906 ();
 sg13g2_decap_8 FILLER_78_1913 ();
 sg13g2_decap_8 FILLER_78_1920 ();
 sg13g2_decap_8 FILLER_78_1927 ();
 sg13g2_decap_8 FILLER_78_1934 ();
 sg13g2_decap_8 FILLER_78_1941 ();
 sg13g2_decap_8 FILLER_78_1948 ();
 sg13g2_decap_8 FILLER_78_1955 ();
 sg13g2_decap_4 FILLER_78_1962 ();
 sg13g2_fill_2 FILLER_78_1966 ();
 sg13g2_decap_4 FILLER_78_1998 ();
 sg13g2_fill_2 FILLER_78_2002 ();
 sg13g2_decap_4 FILLER_78_2038 ();
 sg13g2_fill_1 FILLER_78_2042 ();
 sg13g2_decap_4 FILLER_78_2075 ();
 sg13g2_decap_4 FILLER_78_2083 ();
 sg13g2_fill_2 FILLER_78_2087 ();
 sg13g2_decap_8 FILLER_78_2094 ();
 sg13g2_decap_4 FILLER_78_2101 ();
 sg13g2_fill_2 FILLER_78_2105 ();
 sg13g2_fill_1 FILLER_78_2111 ();
 sg13g2_fill_1 FILLER_78_2121 ();
 sg13g2_fill_2 FILLER_78_2152 ();
 sg13g2_fill_2 FILLER_78_2189 ();
 sg13g2_fill_1 FILLER_78_2225 ();
 sg13g2_decap_4 FILLER_78_2242 ();
 sg13g2_decap_4 FILLER_78_2316 ();
 sg13g2_fill_2 FILLER_78_2334 ();
 sg13g2_fill_1 FILLER_78_2336 ();
 sg13g2_decap_8 FILLER_78_2363 ();
 sg13g2_decap_4 FILLER_78_2370 ();
 sg13g2_fill_2 FILLER_78_2381 ();
 sg13g2_fill_1 FILLER_78_2383 ();
 sg13g2_decap_4 FILLER_78_2399 ();
 sg13g2_decap_4 FILLER_78_2419 ();
 sg13g2_fill_2 FILLER_78_2423 ();
 sg13g2_fill_2 FILLER_78_2457 ();
 sg13g2_fill_2 FILLER_78_2478 ();
 sg13g2_decap_8 FILLER_78_2484 ();
 sg13g2_decap_8 FILLER_78_2491 ();
 sg13g2_decap_8 FILLER_78_2498 ();
 sg13g2_decap_8 FILLER_78_2505 ();
 sg13g2_decap_8 FILLER_78_2516 ();
 sg13g2_decap_8 FILLER_78_2523 ();
 sg13g2_decap_8 FILLER_78_2530 ();
 sg13g2_decap_8 FILLER_78_2537 ();
 sg13g2_decap_8 FILLER_78_2544 ();
 sg13g2_decap_8 FILLER_78_2551 ();
 sg13g2_fill_1 FILLER_78_2558 ();
 sg13g2_decap_8 FILLER_78_2573 ();
 sg13g2_fill_2 FILLER_78_2580 ();
 sg13g2_fill_2 FILLER_78_2608 ();
 sg13g2_fill_1 FILLER_78_2644 ();
 sg13g2_decap_8 FILLER_78_2666 ();
 sg13g2_decap_4 FILLER_78_2673 ();
 sg13g2_fill_1 FILLER_78_2677 ();
 sg13g2_fill_1 FILLER_78_2699 ();
 sg13g2_decap_8 FILLER_78_2726 ();
 sg13g2_decap_4 FILLER_78_2736 ();
 sg13g2_fill_2 FILLER_78_2745 ();
 sg13g2_fill_1 FILLER_78_2747 ();
 sg13g2_fill_1 FILLER_78_2787 ();
 sg13g2_decap_8 FILLER_78_2799 ();
 sg13g2_decap_8 FILLER_78_2806 ();
 sg13g2_fill_1 FILLER_78_2830 ();
 sg13g2_decap_4 FILLER_78_2844 ();
 sg13g2_decap_4 FILLER_78_2862 ();
 sg13g2_decap_8 FILLER_78_2870 ();
 sg13g2_fill_2 FILLER_78_2877 ();
 sg13g2_fill_2 FILLER_78_2892 ();
 sg13g2_fill_1 FILLER_78_2894 ();
 sg13g2_fill_2 FILLER_78_2910 ();
 sg13g2_fill_1 FILLER_78_2912 ();
 sg13g2_decap_8 FILLER_78_2926 ();
 sg13g2_decap_8 FILLER_78_2933 ();
 sg13g2_decap_8 FILLER_78_2940 ();
 sg13g2_decap_8 FILLER_78_2947 ();
 sg13g2_decap_8 FILLER_78_2954 ();
 sg13g2_decap_8 FILLER_78_2961 ();
 sg13g2_decap_8 FILLER_78_2968 ();
 sg13g2_decap_8 FILLER_78_2975 ();
 sg13g2_decap_8 FILLER_78_2982 ();
 sg13g2_decap_8 FILLER_78_2989 ();
 sg13g2_decap_8 FILLER_78_2996 ();
 sg13g2_decap_8 FILLER_78_3003 ();
 sg13g2_decap_8 FILLER_78_3010 ();
 sg13g2_decap_8 FILLER_78_3017 ();
 sg13g2_decap_8 FILLER_78_3024 ();
 sg13g2_decap_8 FILLER_78_3031 ();
 sg13g2_decap_8 FILLER_78_3038 ();
 sg13g2_decap_8 FILLER_78_3045 ();
 sg13g2_decap_8 FILLER_78_3052 ();
 sg13g2_decap_8 FILLER_78_3059 ();
 sg13g2_decap_8 FILLER_78_3066 ();
 sg13g2_decap_8 FILLER_78_3073 ();
 sg13g2_decap_8 FILLER_78_3080 ();
 sg13g2_decap_8 FILLER_78_3087 ();
 sg13g2_decap_8 FILLER_78_3094 ();
 sg13g2_decap_8 FILLER_78_3101 ();
 sg13g2_decap_8 FILLER_78_3108 ();
 sg13g2_decap_8 FILLER_78_3115 ();
 sg13g2_decap_8 FILLER_78_3122 ();
 sg13g2_decap_8 FILLER_78_3129 ();
 sg13g2_decap_8 FILLER_78_3136 ();
 sg13g2_decap_8 FILLER_78_3143 ();
 sg13g2_decap_8 FILLER_78_3150 ();
 sg13g2_decap_8 FILLER_78_3157 ();
 sg13g2_decap_8 FILLER_78_3164 ();
 sg13g2_decap_8 FILLER_78_3171 ();
 sg13g2_decap_8 FILLER_78_3178 ();
 sg13g2_decap_8 FILLER_78_3185 ();
 sg13g2_decap_8 FILLER_78_3192 ();
 sg13g2_decap_8 FILLER_78_3199 ();
 sg13g2_decap_8 FILLER_78_3206 ();
 sg13g2_decap_8 FILLER_78_3213 ();
 sg13g2_decap_8 FILLER_78_3220 ();
 sg13g2_decap_8 FILLER_78_3227 ();
 sg13g2_decap_8 FILLER_78_3234 ();
 sg13g2_decap_8 FILLER_78_3241 ();
 sg13g2_decap_8 FILLER_78_3248 ();
 sg13g2_decap_8 FILLER_78_3255 ();
 sg13g2_decap_8 FILLER_78_3262 ();
 sg13g2_decap_8 FILLER_78_3269 ();
 sg13g2_decap_8 FILLER_78_3276 ();
 sg13g2_decap_8 FILLER_78_3283 ();
 sg13g2_decap_8 FILLER_78_3290 ();
 sg13g2_decap_8 FILLER_78_3297 ();
 sg13g2_decap_8 FILLER_78_3304 ();
 sg13g2_decap_8 FILLER_78_3311 ();
 sg13g2_decap_8 FILLER_78_3318 ();
 sg13g2_decap_8 FILLER_78_3325 ();
 sg13g2_decap_8 FILLER_78_3332 ();
 sg13g2_decap_8 FILLER_78_3339 ();
 sg13g2_decap_8 FILLER_78_3346 ();
 sg13g2_decap_8 FILLER_78_3353 ();
 sg13g2_decap_8 FILLER_78_3360 ();
 sg13g2_decap_8 FILLER_78_3367 ();
 sg13g2_decap_8 FILLER_78_3374 ();
 sg13g2_decap_8 FILLER_78_3381 ();
 sg13g2_decap_8 FILLER_78_3388 ();
 sg13g2_decap_8 FILLER_78_3395 ();
 sg13g2_decap_8 FILLER_78_3402 ();
 sg13g2_decap_8 FILLER_78_3409 ();
 sg13g2_decap_8 FILLER_78_3416 ();
 sg13g2_decap_8 FILLER_78_3423 ();
 sg13g2_decap_8 FILLER_78_3430 ();
 sg13g2_decap_8 FILLER_78_3437 ();
 sg13g2_decap_8 FILLER_78_3444 ();
 sg13g2_decap_8 FILLER_78_3451 ();
 sg13g2_decap_8 FILLER_78_3458 ();
 sg13g2_decap_8 FILLER_78_3465 ();
 sg13g2_decap_8 FILLER_78_3472 ();
 sg13g2_decap_8 FILLER_78_3479 ();
 sg13g2_decap_8 FILLER_78_3486 ();
 sg13g2_decap_8 FILLER_78_3493 ();
 sg13g2_decap_8 FILLER_78_3500 ();
 sg13g2_decap_8 FILLER_78_3507 ();
 sg13g2_decap_8 FILLER_78_3514 ();
 sg13g2_decap_8 FILLER_78_3521 ();
 sg13g2_decap_8 FILLER_78_3528 ();
 sg13g2_decap_8 FILLER_78_3535 ();
 sg13g2_decap_8 FILLER_78_3542 ();
 sg13g2_decap_8 FILLER_78_3549 ();
 sg13g2_decap_8 FILLER_78_3556 ();
 sg13g2_decap_8 FILLER_78_3563 ();
 sg13g2_decap_8 FILLER_78_3570 ();
 sg13g2_fill_2 FILLER_78_3577 ();
 sg13g2_fill_1 FILLER_78_3579 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_decap_8 FILLER_79_154 ();
 sg13g2_decap_8 FILLER_79_161 ();
 sg13g2_decap_8 FILLER_79_168 ();
 sg13g2_decap_8 FILLER_79_175 ();
 sg13g2_decap_8 FILLER_79_182 ();
 sg13g2_decap_8 FILLER_79_189 ();
 sg13g2_decap_8 FILLER_79_196 ();
 sg13g2_decap_8 FILLER_79_203 ();
 sg13g2_decap_8 FILLER_79_210 ();
 sg13g2_decap_8 FILLER_79_217 ();
 sg13g2_decap_8 FILLER_79_224 ();
 sg13g2_fill_2 FILLER_79_231 ();
 sg13g2_fill_2 FILLER_79_267 ();
 sg13g2_fill_1 FILLER_79_269 ();
 sg13g2_fill_1 FILLER_79_287 ();
 sg13g2_fill_2 FILLER_79_296 ();
 sg13g2_fill_1 FILLER_79_323 ();
 sg13g2_fill_1 FILLER_79_383 ();
 sg13g2_fill_2 FILLER_79_410 ();
 sg13g2_fill_2 FILLER_79_445 ();
 sg13g2_fill_1 FILLER_79_473 ();
 sg13g2_fill_2 FILLER_79_483 ();
 sg13g2_fill_2 FILLER_79_494 ();
 sg13g2_fill_2 FILLER_79_505 ();
 sg13g2_fill_1 FILLER_79_507 ();
 sg13g2_fill_2 FILLER_79_513 ();
 sg13g2_fill_1 FILLER_79_515 ();
 sg13g2_fill_2 FILLER_79_525 ();
 sg13g2_fill_1 FILLER_79_527 ();
 sg13g2_fill_1 FILLER_79_567 ();
 sg13g2_fill_2 FILLER_79_582 ();
 sg13g2_fill_2 FILLER_79_647 ();
 sg13g2_decap_8 FILLER_79_688 ();
 sg13g2_fill_1 FILLER_79_695 ();
 sg13g2_decap_8 FILLER_79_700 ();
 sg13g2_decap_8 FILLER_79_707 ();
 sg13g2_fill_1 FILLER_79_714 ();
 sg13g2_fill_1 FILLER_79_767 ();
 sg13g2_fill_2 FILLER_79_794 ();
 sg13g2_fill_1 FILLER_79_830 ();
 sg13g2_fill_2 FILLER_79_918 ();
 sg13g2_fill_1 FILLER_79_920 ();
 sg13g2_fill_1 FILLER_79_947 ();
 sg13g2_fill_2 FILLER_79_964 ();
 sg13g2_decap_8 FILLER_79_1013 ();
 sg13g2_fill_2 FILLER_79_1020 ();
 sg13g2_decap_4 FILLER_79_1029 ();
 sg13g2_decap_8 FILLER_79_1067 ();
 sg13g2_fill_2 FILLER_79_1118 ();
 sg13g2_fill_1 FILLER_79_1120 ();
 sg13g2_decap_4 FILLER_79_1134 ();
 sg13g2_fill_1 FILLER_79_1138 ();
 sg13g2_fill_2 FILLER_79_1149 ();
 sg13g2_fill_1 FILLER_79_1160 ();
 sg13g2_fill_2 FILLER_79_1179 ();
 sg13g2_fill_1 FILLER_79_1181 ();
 sg13g2_fill_2 FILLER_79_1239 ();
 sg13g2_fill_2 FILLER_79_1271 ();
 sg13g2_decap_4 FILLER_79_1299 ();
 sg13g2_fill_2 FILLER_79_1329 ();
 sg13g2_fill_1 FILLER_79_1331 ();
 sg13g2_fill_1 FILLER_79_1372 ();
 sg13g2_decap_8 FILLER_79_1425 ();
 sg13g2_fill_2 FILLER_79_1432 ();
 sg13g2_fill_1 FILLER_79_1434 ();
 sg13g2_decap_4 FILLER_79_1461 ();
 sg13g2_fill_1 FILLER_79_1465 ();
 sg13g2_fill_1 FILLER_79_1506 ();
 sg13g2_fill_2 FILLER_79_1590 ();
 sg13g2_fill_1 FILLER_79_1592 ();
 sg13g2_fill_2 FILLER_79_1660 ();
 sg13g2_fill_1 FILLER_79_1662 ();
 sg13g2_fill_2 FILLER_79_1672 ();
 sg13g2_fill_1 FILLER_79_1674 ();
 sg13g2_fill_1 FILLER_79_1710 ();
 sg13g2_decap_8 FILLER_79_1715 ();
 sg13g2_decap_8 FILLER_79_1722 ();
 sg13g2_decap_8 FILLER_79_1729 ();
 sg13g2_decap_8 FILLER_79_1736 ();
 sg13g2_decap_8 FILLER_79_1743 ();
 sg13g2_decap_8 FILLER_79_1750 ();
 sg13g2_decap_8 FILLER_79_1757 ();
 sg13g2_decap_8 FILLER_79_1764 ();
 sg13g2_decap_8 FILLER_79_1771 ();
 sg13g2_decap_8 FILLER_79_1778 ();
 sg13g2_decap_8 FILLER_79_1785 ();
 sg13g2_decap_8 FILLER_79_1792 ();
 sg13g2_decap_8 FILLER_79_1799 ();
 sg13g2_decap_8 FILLER_79_1806 ();
 sg13g2_decap_8 FILLER_79_1813 ();
 sg13g2_decap_8 FILLER_79_1820 ();
 sg13g2_decap_8 FILLER_79_1827 ();
 sg13g2_decap_8 FILLER_79_1834 ();
 sg13g2_decap_8 FILLER_79_1841 ();
 sg13g2_decap_8 FILLER_79_1848 ();
 sg13g2_decap_8 FILLER_79_1855 ();
 sg13g2_decap_8 FILLER_79_1862 ();
 sg13g2_decap_8 FILLER_79_1869 ();
 sg13g2_decap_8 FILLER_79_1876 ();
 sg13g2_decap_8 FILLER_79_1883 ();
 sg13g2_decap_8 FILLER_79_1890 ();
 sg13g2_decap_8 FILLER_79_1897 ();
 sg13g2_decap_8 FILLER_79_1904 ();
 sg13g2_decap_8 FILLER_79_1911 ();
 sg13g2_decap_8 FILLER_79_1918 ();
 sg13g2_decap_8 FILLER_79_1925 ();
 sg13g2_decap_8 FILLER_79_1932 ();
 sg13g2_decap_8 FILLER_79_1939 ();
 sg13g2_decap_8 FILLER_79_1946 ();
 sg13g2_decap_8 FILLER_79_1953 ();
 sg13g2_decap_8 FILLER_79_1960 ();
 sg13g2_decap_8 FILLER_79_1967 ();
 sg13g2_decap_8 FILLER_79_1974 ();
 sg13g2_decap_8 FILLER_79_1981 ();
 sg13g2_decap_4 FILLER_79_1988 ();
 sg13g2_fill_2 FILLER_79_1992 ();
 sg13g2_fill_2 FILLER_79_1998 ();
 sg13g2_fill_2 FILLER_79_2045 ();
 sg13g2_decap_8 FILLER_79_2065 ();
 sg13g2_decap_8 FILLER_79_2072 ();
 sg13g2_decap_8 FILLER_79_2079 ();
 sg13g2_decap_8 FILLER_79_2086 ();
 sg13g2_decap_8 FILLER_79_2093 ();
 sg13g2_decap_8 FILLER_79_2100 ();
 sg13g2_decap_8 FILLER_79_2107 ();
 sg13g2_decap_8 FILLER_79_2114 ();
 sg13g2_decap_8 FILLER_79_2121 ();
 sg13g2_decap_8 FILLER_79_2128 ();
 sg13g2_fill_2 FILLER_79_2135 ();
 sg13g2_decap_8 FILLER_79_2141 ();
 sg13g2_decap_8 FILLER_79_2148 ();
 sg13g2_fill_1 FILLER_79_2155 ();
 sg13g2_fill_1 FILLER_79_2160 ();
 sg13g2_decap_4 FILLER_79_2169 ();
 sg13g2_fill_2 FILLER_79_2173 ();
 sg13g2_decap_8 FILLER_79_2179 ();
 sg13g2_decap_4 FILLER_79_2186 ();
 sg13g2_fill_1 FILLER_79_2205 ();
 sg13g2_fill_2 FILLER_79_2234 ();
 sg13g2_fill_1 FILLER_79_2236 ();
 sg13g2_decap_8 FILLER_79_2256 ();
 sg13g2_decap_8 FILLER_79_2263 ();
 sg13g2_decap_8 FILLER_79_2270 ();
 sg13g2_fill_1 FILLER_79_2295 ();
 sg13g2_fill_2 FILLER_79_2345 ();
 sg13g2_fill_1 FILLER_79_2347 ();
 sg13g2_decap_8 FILLER_79_2352 ();
 sg13g2_decap_4 FILLER_79_2363 ();
 sg13g2_decap_4 FILLER_79_2371 ();
 sg13g2_fill_2 FILLER_79_2375 ();
 sg13g2_fill_2 FILLER_79_2390 ();
 sg13g2_fill_1 FILLER_79_2392 ();
 sg13g2_fill_2 FILLER_79_2399 ();
 sg13g2_fill_1 FILLER_79_2401 ();
 sg13g2_fill_2 FILLER_79_2430 ();
 sg13g2_fill_1 FILLER_79_2432 ();
 sg13g2_fill_2 FILLER_79_2439 ();
 sg13g2_fill_1 FILLER_79_2441 ();
 sg13g2_fill_1 FILLER_79_2468 ();
 sg13g2_decap_8 FILLER_79_2495 ();
 sg13g2_decap_8 FILLER_79_2502 ();
 sg13g2_decap_8 FILLER_79_2509 ();
 sg13g2_decap_8 FILLER_79_2516 ();
 sg13g2_decap_8 FILLER_79_2523 ();
 sg13g2_decap_8 FILLER_79_2530 ();
 sg13g2_decap_8 FILLER_79_2537 ();
 sg13g2_decap_8 FILLER_79_2544 ();
 sg13g2_decap_8 FILLER_79_2551 ();
 sg13g2_decap_4 FILLER_79_2558 ();
 sg13g2_fill_2 FILLER_79_2610 ();
 sg13g2_decap_8 FILLER_79_2643 ();
 sg13g2_fill_2 FILLER_79_2650 ();
 sg13g2_fill_1 FILLER_79_2661 ();
 sg13g2_decap_4 FILLER_79_2671 ();
 sg13g2_fill_1 FILLER_79_2675 ();
 sg13g2_fill_1 FILLER_79_2694 ();
 sg13g2_decap_8 FILLER_79_2704 ();
 sg13g2_decap_8 FILLER_79_2715 ();
 sg13g2_decap_8 FILLER_79_2722 ();
 sg13g2_decap_4 FILLER_79_2755 ();
 sg13g2_fill_2 FILLER_79_2763 ();
 sg13g2_decap_8 FILLER_79_2769 ();
 sg13g2_decap_8 FILLER_79_2776 ();
 sg13g2_fill_1 FILLER_79_2799 ();
 sg13g2_decap_8 FILLER_79_2805 ();
 sg13g2_fill_2 FILLER_79_2812 ();
 sg13g2_decap_4 FILLER_79_2823 ();
 sg13g2_fill_1 FILLER_79_2827 ();
 sg13g2_fill_2 FILLER_79_2846 ();
 sg13g2_fill_1 FILLER_79_2860 ();
 sg13g2_decap_4 FILLER_79_2865 ();
 sg13g2_fill_2 FILLER_79_2869 ();
 sg13g2_decap_8 FILLER_79_2897 ();
 sg13g2_decap_8 FILLER_79_2904 ();
 sg13g2_decap_8 FILLER_79_2911 ();
 sg13g2_decap_8 FILLER_79_2918 ();
 sg13g2_decap_8 FILLER_79_2925 ();
 sg13g2_decap_8 FILLER_79_2932 ();
 sg13g2_decap_8 FILLER_79_2939 ();
 sg13g2_decap_8 FILLER_79_2946 ();
 sg13g2_decap_8 FILLER_79_2953 ();
 sg13g2_decap_8 FILLER_79_2960 ();
 sg13g2_decap_8 FILLER_79_2967 ();
 sg13g2_decap_8 FILLER_79_2974 ();
 sg13g2_decap_8 FILLER_79_2981 ();
 sg13g2_decap_8 FILLER_79_2988 ();
 sg13g2_decap_8 FILLER_79_2995 ();
 sg13g2_decap_8 FILLER_79_3002 ();
 sg13g2_decap_8 FILLER_79_3009 ();
 sg13g2_decap_8 FILLER_79_3016 ();
 sg13g2_decap_8 FILLER_79_3023 ();
 sg13g2_decap_8 FILLER_79_3030 ();
 sg13g2_decap_8 FILLER_79_3037 ();
 sg13g2_decap_8 FILLER_79_3044 ();
 sg13g2_decap_8 FILLER_79_3051 ();
 sg13g2_decap_8 FILLER_79_3058 ();
 sg13g2_decap_8 FILLER_79_3065 ();
 sg13g2_decap_8 FILLER_79_3072 ();
 sg13g2_decap_8 FILLER_79_3079 ();
 sg13g2_decap_8 FILLER_79_3086 ();
 sg13g2_decap_8 FILLER_79_3093 ();
 sg13g2_decap_8 FILLER_79_3100 ();
 sg13g2_decap_8 FILLER_79_3107 ();
 sg13g2_decap_8 FILLER_79_3114 ();
 sg13g2_decap_8 FILLER_79_3121 ();
 sg13g2_decap_8 FILLER_79_3128 ();
 sg13g2_decap_8 FILLER_79_3135 ();
 sg13g2_decap_8 FILLER_79_3142 ();
 sg13g2_decap_8 FILLER_79_3149 ();
 sg13g2_decap_8 FILLER_79_3156 ();
 sg13g2_decap_8 FILLER_79_3163 ();
 sg13g2_decap_8 FILLER_79_3170 ();
 sg13g2_decap_8 FILLER_79_3177 ();
 sg13g2_decap_8 FILLER_79_3184 ();
 sg13g2_decap_8 FILLER_79_3191 ();
 sg13g2_decap_8 FILLER_79_3198 ();
 sg13g2_decap_8 FILLER_79_3205 ();
 sg13g2_decap_8 FILLER_79_3212 ();
 sg13g2_decap_8 FILLER_79_3219 ();
 sg13g2_decap_8 FILLER_79_3226 ();
 sg13g2_decap_8 FILLER_79_3233 ();
 sg13g2_decap_8 FILLER_79_3240 ();
 sg13g2_decap_8 FILLER_79_3247 ();
 sg13g2_decap_8 FILLER_79_3254 ();
 sg13g2_decap_8 FILLER_79_3261 ();
 sg13g2_decap_8 FILLER_79_3268 ();
 sg13g2_decap_8 FILLER_79_3275 ();
 sg13g2_decap_8 FILLER_79_3282 ();
 sg13g2_decap_8 FILLER_79_3289 ();
 sg13g2_decap_8 FILLER_79_3296 ();
 sg13g2_decap_8 FILLER_79_3303 ();
 sg13g2_decap_8 FILLER_79_3310 ();
 sg13g2_decap_8 FILLER_79_3317 ();
 sg13g2_decap_8 FILLER_79_3324 ();
 sg13g2_decap_8 FILLER_79_3331 ();
 sg13g2_decap_8 FILLER_79_3338 ();
 sg13g2_decap_8 FILLER_79_3345 ();
 sg13g2_decap_8 FILLER_79_3352 ();
 sg13g2_decap_8 FILLER_79_3359 ();
 sg13g2_decap_8 FILLER_79_3366 ();
 sg13g2_decap_8 FILLER_79_3373 ();
 sg13g2_decap_8 FILLER_79_3380 ();
 sg13g2_decap_8 FILLER_79_3387 ();
 sg13g2_decap_8 FILLER_79_3394 ();
 sg13g2_decap_8 FILLER_79_3401 ();
 sg13g2_decap_8 FILLER_79_3408 ();
 sg13g2_decap_8 FILLER_79_3415 ();
 sg13g2_decap_8 FILLER_79_3422 ();
 sg13g2_decap_8 FILLER_79_3429 ();
 sg13g2_decap_8 FILLER_79_3436 ();
 sg13g2_decap_8 FILLER_79_3443 ();
 sg13g2_decap_8 FILLER_79_3450 ();
 sg13g2_decap_8 FILLER_79_3457 ();
 sg13g2_decap_8 FILLER_79_3464 ();
 sg13g2_decap_8 FILLER_79_3471 ();
 sg13g2_decap_8 FILLER_79_3478 ();
 sg13g2_decap_8 FILLER_79_3485 ();
 sg13g2_decap_8 FILLER_79_3492 ();
 sg13g2_decap_8 FILLER_79_3499 ();
 sg13g2_decap_8 FILLER_79_3506 ();
 sg13g2_decap_8 FILLER_79_3513 ();
 sg13g2_decap_8 FILLER_79_3520 ();
 sg13g2_decap_8 FILLER_79_3527 ();
 sg13g2_decap_8 FILLER_79_3534 ();
 sg13g2_decap_8 FILLER_79_3541 ();
 sg13g2_decap_8 FILLER_79_3548 ();
 sg13g2_decap_8 FILLER_79_3555 ();
 sg13g2_decap_8 FILLER_79_3562 ();
 sg13g2_decap_8 FILLER_79_3569 ();
 sg13g2_decap_4 FILLER_79_3576 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_8 FILLER_80_68 ();
 sg13g2_decap_8 FILLER_80_75 ();
 sg13g2_decap_4 FILLER_80_82 ();
 sg13g2_fill_2 FILLER_80_86 ();
 sg13g2_decap_8 FILLER_80_92 ();
 sg13g2_decap_8 FILLER_80_99 ();
 sg13g2_decap_4 FILLER_80_106 ();
 sg13g2_fill_2 FILLER_80_110 ();
 sg13g2_decap_8 FILLER_80_116 ();
 sg13g2_decap_8 FILLER_80_123 ();
 sg13g2_decap_8 FILLER_80_130 ();
 sg13g2_decap_8 FILLER_80_137 ();
 sg13g2_decap_8 FILLER_80_144 ();
 sg13g2_decap_8 FILLER_80_151 ();
 sg13g2_decap_8 FILLER_80_158 ();
 sg13g2_decap_8 FILLER_80_165 ();
 sg13g2_decap_8 FILLER_80_172 ();
 sg13g2_decap_8 FILLER_80_179 ();
 sg13g2_decap_8 FILLER_80_186 ();
 sg13g2_decap_8 FILLER_80_193 ();
 sg13g2_decap_8 FILLER_80_200 ();
 sg13g2_decap_8 FILLER_80_207 ();
 sg13g2_decap_8 FILLER_80_214 ();
 sg13g2_decap_8 FILLER_80_221 ();
 sg13g2_decap_8 FILLER_80_228 ();
 sg13g2_fill_2 FILLER_80_235 ();
 sg13g2_fill_1 FILLER_80_237 ();
 sg13g2_fill_2 FILLER_80_302 ();
 sg13g2_fill_1 FILLER_80_304 ();
 sg13g2_fill_2 FILLER_80_357 ();
 sg13g2_fill_1 FILLER_80_359 ();
 sg13g2_decap_8 FILLER_80_399 ();
 sg13g2_decap_4 FILLER_80_406 ();
 sg13g2_fill_2 FILLER_80_410 ();
 sg13g2_decap_4 FILLER_80_417 ();
 sg13g2_decap_8 FILLER_80_447 ();
 sg13g2_decap_4 FILLER_80_454 ();
 sg13g2_fill_1 FILLER_80_462 ();
 sg13g2_fill_2 FILLER_80_472 ();
 sg13g2_fill_1 FILLER_80_505 ();
 sg13g2_fill_2 FILLER_80_550 ();
 sg13g2_decap_8 FILLER_80_582 ();
 sg13g2_fill_2 FILLER_80_589 ();
 sg13g2_fill_1 FILLER_80_591 ();
 sg13g2_fill_2 FILLER_80_599 ();
 sg13g2_decap_8 FILLER_80_614 ();
 sg13g2_decap_8 FILLER_80_621 ();
 sg13g2_decap_8 FILLER_80_628 ();
 sg13g2_fill_2 FILLER_80_635 ();
 sg13g2_decap_8 FILLER_80_676 ();
 sg13g2_decap_8 FILLER_80_683 ();
 sg13g2_decap_8 FILLER_80_690 ();
 sg13g2_decap_8 FILLER_80_697 ();
 sg13g2_decap_8 FILLER_80_704 ();
 sg13g2_decap_8 FILLER_80_711 ();
 sg13g2_decap_8 FILLER_80_718 ();
 sg13g2_fill_2 FILLER_80_732 ();
 sg13g2_fill_2 FILLER_80_741 ();
 sg13g2_fill_1 FILLER_80_751 ();
 sg13g2_decap_8 FILLER_80_756 ();
 sg13g2_decap_8 FILLER_80_763 ();
 sg13g2_fill_1 FILLER_80_770 ();
 sg13g2_fill_2 FILLER_80_775 ();
 sg13g2_fill_1 FILLER_80_777 ();
 sg13g2_fill_1 FILLER_80_782 ();
 sg13g2_fill_1 FILLER_80_811 ();
 sg13g2_decap_4 FILLER_80_826 ();
 sg13g2_decap_8 FILLER_80_847 ();
 sg13g2_fill_1 FILLER_80_854 ();
 sg13g2_decap_4 FILLER_80_859 ();
 sg13g2_fill_2 FILLER_80_867 ();
 sg13g2_decap_8 FILLER_80_885 ();
 sg13g2_decap_4 FILLER_80_892 ();
 sg13g2_fill_1 FILLER_80_896 ();
 sg13g2_fill_2 FILLER_80_901 ();
 sg13g2_decap_8 FILLER_80_907 ();
 sg13g2_decap_8 FILLER_80_914 ();
 sg13g2_decap_4 FILLER_80_982 ();
 sg13g2_decap_8 FILLER_80_1008 ();
 sg13g2_decap_8 FILLER_80_1015 ();
 sg13g2_decap_8 FILLER_80_1022 ();
 sg13g2_decap_4 FILLER_80_1029 ();
 sg13g2_fill_1 FILLER_80_1033 ();
 sg13g2_fill_2 FILLER_80_1038 ();
 sg13g2_fill_1 FILLER_80_1040 ();
 sg13g2_decap_8 FILLER_80_1063 ();
 sg13g2_decap_8 FILLER_80_1070 ();
 sg13g2_fill_2 FILLER_80_1077 ();
 sg13g2_fill_1 FILLER_80_1088 ();
 sg13g2_decap_4 FILLER_80_1093 ();
 sg13g2_fill_1 FILLER_80_1136 ();
 sg13g2_fill_2 FILLER_80_1142 ();
 sg13g2_decap_8 FILLER_80_1174 ();
 sg13g2_decap_4 FILLER_80_1181 ();
 sg13g2_fill_2 FILLER_80_1220 ();
 sg13g2_fill_1 FILLER_80_1222 ();
 sg13g2_fill_2 FILLER_80_1237 ();
 sg13g2_fill_1 FILLER_80_1253 ();
 sg13g2_fill_2 FILLER_80_1275 ();
 sg13g2_fill_2 FILLER_80_1281 ();
 sg13g2_fill_1 FILLER_80_1315 ();
 sg13g2_decap_8 FILLER_80_1329 ();
 sg13g2_decap_8 FILLER_80_1336 ();
 sg13g2_fill_1 FILLER_80_1343 ();
 sg13g2_decap_8 FILLER_80_1398 ();
 sg13g2_decap_4 FILLER_80_1405 ();
 sg13g2_fill_1 FILLER_80_1409 ();
 sg13g2_decap_8 FILLER_80_1414 ();
 sg13g2_decap_8 FILLER_80_1421 ();
 sg13g2_decap_8 FILLER_80_1428 ();
 sg13g2_decap_8 FILLER_80_1435 ();
 sg13g2_fill_2 FILLER_80_1442 ();
 sg13g2_fill_1 FILLER_80_1444 ();
 sg13g2_decap_8 FILLER_80_1449 ();
 sg13g2_fill_1 FILLER_80_1456 ();
 sg13g2_decap_8 FILLER_80_1466 ();
 sg13g2_decap_4 FILLER_80_1473 ();
 sg13g2_decap_8 FILLER_80_1481 ();
 sg13g2_decap_4 FILLER_80_1488 ();
 sg13g2_fill_2 FILLER_80_1492 ();
 sg13g2_decap_4 FILLER_80_1499 ();
 sg13g2_fill_1 FILLER_80_1503 ();
 sg13g2_decap_8 FILLER_80_1508 ();
 sg13g2_fill_1 FILLER_80_1529 ();
 sg13g2_fill_2 FILLER_80_1534 ();
 sg13g2_fill_1 FILLER_80_1536 ();
 sg13g2_decap_8 FILLER_80_1542 ();
 sg13g2_fill_1 FILLER_80_1549 ();
 sg13g2_fill_2 FILLER_80_1563 ();
 sg13g2_decap_4 FILLER_80_1570 ();
 sg13g2_decap_8 FILLER_80_1578 ();
 sg13g2_decap_8 FILLER_80_1585 ();
 sg13g2_decap_4 FILLER_80_1592 ();
 sg13g2_decap_4 FILLER_80_1600 ();
 sg13g2_fill_2 FILLER_80_1604 ();
 sg13g2_decap_4 FILLER_80_1615 ();
 sg13g2_decap_8 FILLER_80_1628 ();
 sg13g2_decap_4 FILLER_80_1635 ();
 sg13g2_decap_8 FILLER_80_1643 ();
 sg13g2_fill_2 FILLER_80_1650 ();
 sg13g2_fill_1 FILLER_80_1652 ();
 sg13g2_decap_8 FILLER_80_1696 ();
 sg13g2_decap_8 FILLER_80_1703 ();
 sg13g2_decap_8 FILLER_80_1710 ();
 sg13g2_decap_8 FILLER_80_1717 ();
 sg13g2_decap_8 FILLER_80_1724 ();
 sg13g2_decap_8 FILLER_80_1731 ();
 sg13g2_decap_8 FILLER_80_1738 ();
 sg13g2_decap_8 FILLER_80_1745 ();
 sg13g2_decap_8 FILLER_80_1752 ();
 sg13g2_decap_8 FILLER_80_1759 ();
 sg13g2_decap_8 FILLER_80_1766 ();
 sg13g2_decap_8 FILLER_80_1773 ();
 sg13g2_decap_8 FILLER_80_1780 ();
 sg13g2_decap_8 FILLER_80_1787 ();
 sg13g2_decap_8 FILLER_80_1794 ();
 sg13g2_decap_8 FILLER_80_1801 ();
 sg13g2_decap_8 FILLER_80_1808 ();
 sg13g2_decap_8 FILLER_80_1815 ();
 sg13g2_decap_8 FILLER_80_1822 ();
 sg13g2_decap_8 FILLER_80_1829 ();
 sg13g2_decap_8 FILLER_80_1836 ();
 sg13g2_decap_8 FILLER_80_1843 ();
 sg13g2_decap_8 FILLER_80_1850 ();
 sg13g2_decap_8 FILLER_80_1857 ();
 sg13g2_decap_8 FILLER_80_1864 ();
 sg13g2_decap_8 FILLER_80_1871 ();
 sg13g2_decap_8 FILLER_80_1878 ();
 sg13g2_decap_8 FILLER_80_1885 ();
 sg13g2_decap_8 FILLER_80_1892 ();
 sg13g2_decap_8 FILLER_80_1899 ();
 sg13g2_decap_8 FILLER_80_1906 ();
 sg13g2_decap_8 FILLER_80_1913 ();
 sg13g2_decap_8 FILLER_80_1920 ();
 sg13g2_decap_8 FILLER_80_1927 ();
 sg13g2_decap_8 FILLER_80_1934 ();
 sg13g2_decap_8 FILLER_80_1941 ();
 sg13g2_decap_8 FILLER_80_1948 ();
 sg13g2_decap_8 FILLER_80_1955 ();
 sg13g2_decap_8 FILLER_80_1962 ();
 sg13g2_decap_8 FILLER_80_1969 ();
 sg13g2_decap_8 FILLER_80_1976 ();
 sg13g2_fill_1 FILLER_80_1983 ();
 sg13g2_fill_2 FILLER_80_2010 ();
 sg13g2_decap_8 FILLER_80_2038 ();
 sg13g2_decap_8 FILLER_80_2045 ();
 sg13g2_decap_8 FILLER_80_2052 ();
 sg13g2_decap_8 FILLER_80_2059 ();
 sg13g2_decap_8 FILLER_80_2066 ();
 sg13g2_decap_8 FILLER_80_2073 ();
 sg13g2_decap_8 FILLER_80_2080 ();
 sg13g2_decap_8 FILLER_80_2087 ();
 sg13g2_decap_8 FILLER_80_2094 ();
 sg13g2_decap_8 FILLER_80_2101 ();
 sg13g2_decap_8 FILLER_80_2108 ();
 sg13g2_decap_8 FILLER_80_2115 ();
 sg13g2_decap_8 FILLER_80_2122 ();
 sg13g2_decap_8 FILLER_80_2129 ();
 sg13g2_decap_8 FILLER_80_2136 ();
 sg13g2_decap_8 FILLER_80_2143 ();
 sg13g2_decap_8 FILLER_80_2150 ();
 sg13g2_decap_8 FILLER_80_2157 ();
 sg13g2_decap_4 FILLER_80_2230 ();
 sg13g2_decap_4 FILLER_80_2260 ();
 sg13g2_fill_2 FILLER_80_2264 ();
 sg13g2_fill_2 FILLER_80_2296 ();
 sg13g2_decap_8 FILLER_80_2346 ();
 sg13g2_fill_2 FILLER_80_2353 ();
 sg13g2_fill_1 FILLER_80_2355 ();
 sg13g2_fill_1 FILLER_80_2410 ();
 sg13g2_decap_8 FILLER_80_2416 ();
 sg13g2_decap_8 FILLER_80_2427 ();
 sg13g2_decap_4 FILLER_80_2460 ();
 sg13g2_fill_2 FILLER_80_2464 ();
 sg13g2_decap_8 FILLER_80_2475 ();
 sg13g2_decap_8 FILLER_80_2482 ();
 sg13g2_decap_8 FILLER_80_2489 ();
 sg13g2_decap_8 FILLER_80_2496 ();
 sg13g2_decap_8 FILLER_80_2503 ();
 sg13g2_decap_8 FILLER_80_2510 ();
 sg13g2_decap_8 FILLER_80_2517 ();
 sg13g2_decap_8 FILLER_80_2524 ();
 sg13g2_decap_8 FILLER_80_2531 ();
 sg13g2_decap_8 FILLER_80_2538 ();
 sg13g2_decap_8 FILLER_80_2545 ();
 sg13g2_decap_8 FILLER_80_2552 ();
 sg13g2_decap_8 FILLER_80_2559 ();
 sg13g2_decap_8 FILLER_80_2566 ();
 sg13g2_decap_8 FILLER_80_2577 ();
 sg13g2_decap_8 FILLER_80_2584 ();
 sg13g2_decap_4 FILLER_80_2591 ();
 sg13g2_decap_4 FILLER_80_2634 ();
 sg13g2_fill_2 FILLER_80_2638 ();
 sg13g2_decap_4 FILLER_80_2670 ();
 sg13g2_decap_8 FILLER_80_2709 ();
 sg13g2_decap_8 FILLER_80_2716 ();
 sg13g2_decap_8 FILLER_80_2723 ();
 sg13g2_decap_8 FILLER_80_2730 ();
 sg13g2_fill_2 FILLER_80_2737 ();
 sg13g2_fill_1 FILLER_80_2739 ();
 sg13g2_decap_8 FILLER_80_2744 ();
 sg13g2_decap_8 FILLER_80_2751 ();
 sg13g2_decap_8 FILLER_80_2758 ();
 sg13g2_decap_8 FILLER_80_2765 ();
 sg13g2_decap_8 FILLER_80_2772 ();
 sg13g2_fill_2 FILLER_80_2779 ();
 sg13g2_fill_1 FILLER_80_2781 ();
 sg13g2_fill_1 FILLER_80_2817 ();
 sg13g2_decap_4 FILLER_80_2844 ();
 sg13g2_fill_2 FILLER_80_2848 ();
 sg13g2_decap_8 FILLER_80_2876 ();
 sg13g2_decap_8 FILLER_80_2883 ();
 sg13g2_decap_8 FILLER_80_2890 ();
 sg13g2_decap_8 FILLER_80_2897 ();
 sg13g2_decap_8 FILLER_80_2904 ();
 sg13g2_decap_8 FILLER_80_2911 ();
 sg13g2_decap_8 FILLER_80_2918 ();
 sg13g2_decap_8 FILLER_80_2925 ();
 sg13g2_decap_8 FILLER_80_2932 ();
 sg13g2_decap_8 FILLER_80_2939 ();
 sg13g2_decap_8 FILLER_80_2946 ();
 sg13g2_decap_8 FILLER_80_2953 ();
 sg13g2_decap_8 FILLER_80_2960 ();
 sg13g2_decap_8 FILLER_80_2967 ();
 sg13g2_decap_8 FILLER_80_2974 ();
 sg13g2_decap_8 FILLER_80_2981 ();
 sg13g2_decap_8 FILLER_80_2988 ();
 sg13g2_decap_8 FILLER_80_2995 ();
 sg13g2_decap_8 FILLER_80_3002 ();
 sg13g2_decap_8 FILLER_80_3009 ();
 sg13g2_decap_8 FILLER_80_3016 ();
 sg13g2_decap_8 FILLER_80_3023 ();
 sg13g2_decap_8 FILLER_80_3030 ();
 sg13g2_decap_8 FILLER_80_3037 ();
 sg13g2_decap_8 FILLER_80_3044 ();
 sg13g2_decap_8 FILLER_80_3051 ();
 sg13g2_decap_8 FILLER_80_3058 ();
 sg13g2_decap_8 FILLER_80_3065 ();
 sg13g2_decap_8 FILLER_80_3072 ();
 sg13g2_decap_8 FILLER_80_3079 ();
 sg13g2_decap_8 FILLER_80_3086 ();
 sg13g2_decap_8 FILLER_80_3093 ();
 sg13g2_decap_8 FILLER_80_3100 ();
 sg13g2_decap_8 FILLER_80_3107 ();
 sg13g2_decap_8 FILLER_80_3114 ();
 sg13g2_decap_8 FILLER_80_3121 ();
 sg13g2_decap_8 FILLER_80_3128 ();
 sg13g2_decap_8 FILLER_80_3135 ();
 sg13g2_decap_8 FILLER_80_3142 ();
 sg13g2_decap_8 FILLER_80_3149 ();
 sg13g2_decap_8 FILLER_80_3156 ();
 sg13g2_decap_8 FILLER_80_3163 ();
 sg13g2_decap_8 FILLER_80_3170 ();
 sg13g2_decap_8 FILLER_80_3177 ();
 sg13g2_decap_8 FILLER_80_3184 ();
 sg13g2_decap_8 FILLER_80_3191 ();
 sg13g2_decap_8 FILLER_80_3198 ();
 sg13g2_decap_8 FILLER_80_3205 ();
 sg13g2_decap_8 FILLER_80_3212 ();
 sg13g2_decap_8 FILLER_80_3219 ();
 sg13g2_decap_8 FILLER_80_3226 ();
 sg13g2_decap_8 FILLER_80_3233 ();
 sg13g2_decap_8 FILLER_80_3240 ();
 sg13g2_decap_8 FILLER_80_3247 ();
 sg13g2_decap_8 FILLER_80_3254 ();
 sg13g2_decap_8 FILLER_80_3261 ();
 sg13g2_decap_8 FILLER_80_3268 ();
 sg13g2_decap_8 FILLER_80_3275 ();
 sg13g2_decap_8 FILLER_80_3282 ();
 sg13g2_decap_8 FILLER_80_3289 ();
 sg13g2_decap_8 FILLER_80_3296 ();
 sg13g2_decap_8 FILLER_80_3303 ();
 sg13g2_decap_8 FILLER_80_3310 ();
 sg13g2_decap_8 FILLER_80_3317 ();
 sg13g2_decap_8 FILLER_80_3324 ();
 sg13g2_decap_8 FILLER_80_3331 ();
 sg13g2_decap_8 FILLER_80_3338 ();
 sg13g2_decap_8 FILLER_80_3345 ();
 sg13g2_decap_8 FILLER_80_3352 ();
 sg13g2_decap_8 FILLER_80_3359 ();
 sg13g2_decap_8 FILLER_80_3366 ();
 sg13g2_decap_8 FILLER_80_3373 ();
 sg13g2_decap_8 FILLER_80_3380 ();
 sg13g2_decap_8 FILLER_80_3387 ();
 sg13g2_decap_8 FILLER_80_3394 ();
 sg13g2_decap_8 FILLER_80_3401 ();
 sg13g2_decap_8 FILLER_80_3408 ();
 sg13g2_decap_8 FILLER_80_3415 ();
 sg13g2_decap_8 FILLER_80_3422 ();
 sg13g2_decap_8 FILLER_80_3429 ();
 sg13g2_decap_8 FILLER_80_3436 ();
 sg13g2_decap_8 FILLER_80_3443 ();
 sg13g2_decap_8 FILLER_80_3450 ();
 sg13g2_decap_8 FILLER_80_3457 ();
 sg13g2_decap_8 FILLER_80_3464 ();
 sg13g2_decap_8 FILLER_80_3471 ();
 sg13g2_decap_8 FILLER_80_3478 ();
 sg13g2_decap_8 FILLER_80_3485 ();
 sg13g2_decap_8 FILLER_80_3492 ();
 sg13g2_decap_8 FILLER_80_3499 ();
 sg13g2_decap_8 FILLER_80_3506 ();
 sg13g2_decap_8 FILLER_80_3513 ();
 sg13g2_decap_8 FILLER_80_3520 ();
 sg13g2_decap_8 FILLER_80_3527 ();
 sg13g2_decap_8 FILLER_80_3534 ();
 sg13g2_decap_8 FILLER_80_3541 ();
 sg13g2_decap_8 FILLER_80_3548 ();
 sg13g2_decap_8 FILLER_80_3555 ();
 sg13g2_decap_8 FILLER_80_3562 ();
 sg13g2_decap_8 FILLER_80_3569 ();
 sg13g2_decap_4 FILLER_80_3576 ();
 assign uio_oe[0] = net2594;
 assign uio_oe[3] = net2595;
 assign uio_oe[6] = net2596;
 assign uio_oe[7] = net2597;
endmodule
