module tt_um_rte_eink_driver (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire clk_regs;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire \counter[0] ;
 wire \counter[10] ;
 wire \counter[11] ;
 wire \counter[12] ;
 wire \counter[13] ;
 wire \counter[14] ;
 wire \counter[15] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire \counter[9] ;
 wire csb;
 wire \data_out[0] ;
 wire \data_out[1] ;
 wire \data_out[2] ;
 wire \data_out[3] ;
 wire \data_out[4] ;
 wire \data_out[5] ;
 wire \data_out[6] ;
 wire \data_out[7] ;
 wire dcb;
 wire \inbuf[0] ;
 wire \inbuf[1] ;
 wire \inbuf[2] ;
 wire \inbuf[3] ;
 wire \inbuf[4] ;
 wire \inbuf[5] ;
 wire \inbuf[6] ;
 wire \inbuf[7] ;
 wire \inval[0] ;
 wire \inval[1] ;
 wire \inval[2] ;
 wire \inval[3] ;
 wire \inval[4] ;
 wire \inval[5] ;
 wire \inval[6] ;
 wire \inval[7] ;
 wire mosi;
 wire resetb;
 wire sck;
 wire \spi.count[0] ;
 wire \spi.count[1] ;
 wire \spi.count[2] ;
 wire \spi.count[3] ;
 wire \spi.count[4] ;
 wire \spi.count[5] ;
 wire \spi.count[6] ;
 wire \spi.count[7] ;
 wire \spi.d_latched[0] ;
 wire \spi.d_latched[1] ;
 wire \spi.d_latched[2] ;
 wire \spi.d_latched[3] ;
 wire \spi.d_latched[4] ;
 wire \spi.d_latched[5] ;
 wire \spi.d_latched[6] ;
 wire \spi.d_latched[7] ;
 wire \spi.done ;
 wire \spi.hsck ;
 wire \spi.nbit[0] ;
 wire \spi.nbit[1] ;
 wire \spi.nbit[2] ;
 wire \spi.reg_dat_we ;
 wire \spi.state[0] ;
 wire \spi.state[1] ;
 wire \spi.state[2] ;
 wire \spi.state[3] ;
 wire \spi.stream ;
 wire \spi.treg[0] ;
 wire \spi.treg[1] ;
 wire \spi.treg[2] ;
 wire \spi.treg[3] ;
 wire \spi.treg[4] ;
 wire \spi.treg[5] ;
 wire \spi.treg[6] ;
 wire \spi.treg[7] ;
 wire \spi.w_latched ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire \state[4] ;
 wire stream;
 wire \timer[0] ;
 wire \timer[1] ;
 wire \timer[2] ;
 wire \timer[3] ;
 wire net23;
 wire net11;
 wire net24;
 wire net25;
 wire net26;
 wire net12;
 wire net27;
 wire net13;
 wire net28;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_4_0_0_clk_regs;
 wire clknet_4_1_0_clk_regs;
 wire clknet_4_2_0_clk_regs;
 wire clknet_4_3_0_clk_regs;
 wire clknet_4_4_0_clk_regs;
 wire clknet_4_5_0_clk_regs;
 wire clknet_4_6_0_clk_regs;
 wire clknet_4_7_0_clk_regs;
 wire clknet_4_8_0_clk_regs;
 wire clknet_4_9_0_clk_regs;
 wire clknet_4_10_0_clk_regs;
 wire clknet_4_11_0_clk_regs;
 wire clknet_4_12_0_clk_regs;
 wire clknet_4_13_0_clk_regs;
 wire clknet_4_14_0_clk_regs;
 wire clknet_4_15_0_clk_regs;
 wire delaynet_0_clk;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;

 sg13g2_inv_1 _0606_ (.Y(_0105_),
    .A(net66));
 sg13g2_inv_1 _0607_ (.Y(_0106_),
    .A(net67));
 sg13g2_inv_1 _0608_ (.Y(_0107_),
    .A(_0031_));
 sg13g2_inv_1 _0609_ (.Y(_0108_),
    .A(net144));
 sg13g2_inv_1 _0610_ (.Y(_0109_),
    .A(\spi.state[0] ));
 sg13g2_inv_1 _0611_ (.Y(_0110_),
    .A(\spi.state[1] ));
 sg13g2_inv_2 _0612_ (.Y(_0111_),
    .A(net165));
 sg13g2_inv_1 _0613_ (.Y(_0112_),
    .A(net162));
 sg13g2_inv_2 _0614_ (.Y(_0113_),
    .A(net117));
 sg13g2_inv_1 _0615_ (.Y(_0114_),
    .A(\counter[13] ));
 sg13g2_inv_1 _0616_ (.Y(_0115_),
    .A(net119));
 sg13g2_inv_1 _0617_ (.Y(_0116_),
    .A(\spi.done ));
 sg13g2_inv_1 _0618_ (.Y(_0117_),
    .A(net70));
 sg13g2_inv_1 _0619_ (.Y(_0118_),
    .A(\inval[0] ));
 sg13g2_inv_1 _0620_ (.Y(_0119_),
    .A(\inval[2] ));
 sg13g2_inv_1 _0621_ (.Y(_0120_),
    .A(\inbuf[2] ));
 sg13g2_inv_1 _0622_ (.Y(_0121_),
    .A(\inval[3] ));
 sg13g2_inv_1 _0623_ (.Y(_0122_),
    .A(\inval[4] ));
 sg13g2_inv_1 _0624_ (.Y(_0123_),
    .A(\inbuf[4] ));
 sg13g2_inv_1 _0625_ (.Y(_0124_),
    .A(net84));
 sg13g2_inv_1 _0626_ (.Y(_0125_),
    .A(\spi.treg[7] ));
 sg13g2_inv_1 _0627_ (.Y(_0126_),
    .A(_0019_));
 sg13g2_inv_1 _0628_ (.Y(uio_oe[1]),
    .A(csb));
 sg13g2_inv_1 _1114__2 (.Y(net29),
    .A(clknet_1_0__leaf_clk));
 sg13g2_nor2_2 _0630_ (.A(\spi.state[1] ),
    .B(\spi.state[2] ),
    .Y(_0127_));
 sg13g2_a21oi_1 _0631_ (.A1(\spi.w_latched ),
    .A2(_0116_),
    .Y(_0128_),
    .B1(_0015_));
 sg13g2_nand2_2 _0632_ (.Y(_0129_),
    .A(_0127_),
    .B(_0128_));
 sg13g2_mux2_1 _0633_ (.A0(\data_out[7] ),
    .A1(net74),
    .S(net142),
    .X(_0104_));
 sg13g2_mux2_1 _0634_ (.A0(\data_out[6] ),
    .A1(net80),
    .S(_0129_),
    .X(_0103_));
 sg13g2_mux2_1 _0635_ (.A0(\data_out[5] ),
    .A1(net88),
    .S(net142),
    .X(_0102_));
 sg13g2_nand2_1 _0636_ (.Y(_0130_),
    .A(net65),
    .B(net142));
 sg13g2_o21ai_1 _0637_ (.B1(_0130_),
    .Y(_0101_),
    .A1(_0105_),
    .A2(net142));
 sg13g2_mux2_1 _0638_ (.A0(\data_out[3] ),
    .A1(net91),
    .S(net142),
    .X(_0100_));
 sg13g2_mux2_1 _0639_ (.A0(\data_out[2] ),
    .A1(net94),
    .S(net142),
    .X(_0099_));
 sg13g2_nand2_1 _0640_ (.Y(_0131_),
    .A(net64),
    .B(net142));
 sg13g2_o21ai_1 _0641_ (.B1(_0131_),
    .Y(_0098_),
    .A1(_0106_),
    .A2(net142));
 sg13g2_mux2_1 _0642_ (.A0(\data_out[0] ),
    .A1(net99),
    .S(_0129_),
    .X(_0097_));
 sg13g2_o21ai_1 _0643_ (.B1(_0127_),
    .Y(_0132_),
    .A1(net144),
    .A2(\spi.reg_dat_we ));
 sg13g2_o21ai_1 _0644_ (.B1(_0132_),
    .Y(_0044_),
    .A1(_0108_),
    .A2(_0015_));
 sg13g2_a21oi_1 _0645_ (.A1(_0108_),
    .A2(\spi.state[0] ),
    .Y(_0033_),
    .B1(\spi.state[3] ));
 sg13g2_nand2_1 _0646_ (.Y(_0133_),
    .A(\spi.nbit[0] ),
    .B(\spi.nbit[1] ));
 sg13g2_o21ai_1 _0647_ (.B1(\spi.state[1] ),
    .Y(_0134_),
    .A1(_0013_),
    .A2(_0133_));
 sg13g2_nand2_1 _0648_ (.Y(_0135_),
    .A(net144),
    .B(\spi.state[0] ));
 sg13g2_nand2_1 _0649_ (.Y(_0001_),
    .A(_0134_),
    .B(_0135_));
 sg13g2_or4_1 _0650_ (.A(\spi.count[5] ),
    .B(\spi.count[4] ),
    .C(net59),
    .D(net68),
    .X(_0136_));
 sg13g2_nand2b_1 _0651_ (.Y(_0137_),
    .B(net95),
    .A_N(net62));
 sg13g2_nor4_2 _0652_ (.A(net84),
    .B(\spi.count[2] ),
    .C(_0136_),
    .Y(_0138_),
    .D(_0137_));
 sg13g2_nor2_1 _0653_ (.A(net62),
    .B(_0138_),
    .Y(_0002_));
 sg13g2_xnor2_1 _0654_ (.Y(_0139_),
    .A(net62),
    .B(net95));
 sg13g2_nor2_1 _0655_ (.A(_0138_),
    .B(_0139_),
    .Y(_0003_));
 sg13g2_nand3_1 _0656_ (.B(net95),
    .C(net111),
    .A(net62),
    .Y(_0140_));
 sg13g2_a21o_1 _0657_ (.A2(net95),
    .A1(net62),
    .B1(net111),
    .X(_0141_));
 sg13g2_and2_1 _0658_ (.A(_0140_),
    .B(_0141_),
    .X(_0004_));
 sg13g2_nor2_2 _0659_ (.A(_0124_),
    .B(_0140_),
    .Y(_0142_));
 sg13g2_xnor2_1 _0660_ (.Y(_0005_),
    .A(net84),
    .B(_0140_));
 sg13g2_xor2_1 _0661_ (.B(_0142_),
    .A(net86),
    .X(_0006_));
 sg13g2_nand3_1 _0662_ (.B(net86),
    .C(_0142_),
    .A(net112),
    .Y(_0143_));
 sg13g2_a21o_1 _0663_ (.A2(_0142_),
    .A1(net86),
    .B1(net112),
    .X(_0144_));
 sg13g2_and2_1 _0664_ (.A(_0143_),
    .B(_0144_),
    .X(_0007_));
 sg13g2_nand4_1 _0665_ (.B(\spi.count[4] ),
    .C(\spi.count[6] ),
    .A(\spi.count[5] ),
    .Y(_0145_),
    .D(_0142_));
 sg13g2_xnor2_1 _0666_ (.Y(_0008_),
    .A(net68),
    .B(_0143_));
 sg13g2_xnor2_1 _0667_ (.Y(_0009_),
    .A(net59),
    .B(_0145_));
 sg13g2_nor3_1 _0668_ (.A(\spi.state[0] ),
    .B(sck),
    .C(\spi.state[3] ),
    .Y(_0010_));
 sg13g2_nor3_1 _0669_ (.A(_0110_),
    .B(_0013_),
    .C(_0133_),
    .Y(_0000_));
 sg13g2_nor2_1 _0670_ (.A(net143),
    .B(_0021_),
    .Y(_0146_));
 sg13g2_a21oi_1 _0671_ (.A1(\spi.d_latched[0] ),
    .A2(net143),
    .Y(_0043_),
    .B1(_0146_));
 sg13g2_nor2_1 _0672_ (.A(\counter[4] ),
    .B(\counter[5] ),
    .Y(_0147_));
 sg13g2_nand2b_2 _0673_ (.Y(_0148_),
    .B(net163),
    .A_N(net165));
 sg13g2_nand2_2 _0674_ (.Y(_0149_),
    .A(net159),
    .B(net160));
 sg13g2_nor2_1 _0675_ (.A(_0148_),
    .B(_0149_),
    .Y(_0150_));
 sg13g2_nand2_1 _0676_ (.Y(_0151_),
    .A(_0147_),
    .B(_0150_));
 sg13g2_nor2b_2 _0677_ (.A(net106),
    .B_N(\counter[4] ),
    .Y(_0152_));
 sg13g2_nor2_2 _0678_ (.A(net164),
    .B(net162),
    .Y(_0153_));
 sg13g2_nand2b_2 _0679_ (.Y(_0154_),
    .B(net160),
    .A_N(net159));
 sg13g2_and2_1 _0680_ (.A(net160),
    .B(_0153_),
    .X(_0155_));
 sg13g2_nor3_2 _0681_ (.A(net164),
    .B(net162),
    .C(_0154_),
    .Y(_0156_));
 sg13g2_nor2_2 _0682_ (.A(net158),
    .B(net161),
    .Y(_0157_));
 sg13g2_nand2b_2 _0683_ (.Y(_0158_),
    .B(net165),
    .A_N(net162));
 sg13g2_nor3_2 _0684_ (.A(net158),
    .B(net161),
    .C(_0158_),
    .Y(_0159_));
 sg13g2_nand2_1 _0685_ (.Y(_0160_),
    .A(net145),
    .B(_0156_));
 sg13g2_o21ai_1 _0686_ (.B1(net145),
    .Y(_0161_),
    .A1(_0156_),
    .A2(_0159_));
 sg13g2_nand2_2 _0687_ (.Y(_0162_),
    .A(net146),
    .B(_0156_));
 sg13g2_nor2_1 _0688_ (.A(net158),
    .B(_0148_),
    .Y(_0163_));
 sg13g2_nor2b_2 _0689_ (.A(_0148_),
    .B_N(_0157_),
    .Y(_0164_));
 sg13g2_nand2_1 _0690_ (.Y(_0165_),
    .A(net146),
    .B(_0164_));
 sg13g2_o21ai_1 _0691_ (.B1(net146),
    .Y(_0166_),
    .A1(_0156_),
    .A2(_0164_));
 sg13g2_nand2b_2 _0692_ (.Y(_0167_),
    .B(net158),
    .A_N(net160));
 sg13g2_nor2_2 _0693_ (.A(_0158_),
    .B(_0167_),
    .Y(_0168_));
 sg13g2_nor2_2 _0694_ (.A(_0149_),
    .B(_0158_),
    .Y(_0169_));
 sg13g2_and2_1 _0695_ (.A(_0152_),
    .B(_0169_),
    .X(_0170_));
 sg13g2_and2_1 _0696_ (.A(_0153_),
    .B(_0157_),
    .X(_0171_));
 sg13g2_nand2_1 _0697_ (.Y(_0172_),
    .A(net146),
    .B(_0171_));
 sg13g2_a221oi_1 _0698_ (.B2(net147),
    .C1(_0170_),
    .B1(_0171_),
    .A1(net145),
    .Y(_0173_),
    .A2(_0168_));
 sg13g2_nand4_1 _0699_ (.B(_0161_),
    .C(_0166_),
    .A(_0151_),
    .Y(_0174_),
    .D(_0173_));
 sg13g2_and3_1 _0700_ (.X(_0175_),
    .A(net158),
    .B(net147),
    .C(_0153_));
 sg13g2_nor4_2 _0701_ (.A(\counter[4] ),
    .B(\counter[5] ),
    .C(_0148_),
    .Y(_0176_),
    .D(_0154_));
 sg13g2_nor3_1 _0702_ (.A(_0174_),
    .B(_0175_),
    .C(_0176_),
    .Y(_0177_));
 sg13g2_nand2_1 _0703_ (.Y(_0178_),
    .A(net169),
    .B(net168));
 sg13g2_nand3b_1 _0704_ (.B(_0012_),
    .C(\state[3] ),
    .Y(_0179_),
    .A_N(\state[2] ));
 sg13g2_inv_1 _0705_ (.Y(_0180_),
    .A(_0179_));
 sg13g2_nand3_1 _0706_ (.B(\state[1] ),
    .C(net166),
    .A(net169),
    .Y(_0181_));
 sg13g2_nor2_2 _0707_ (.A(_0178_),
    .B(_0179_),
    .Y(_0182_));
 sg13g2_nand2_2 _0708_ (.Y(_0183_),
    .A(net164),
    .B(net162));
 sg13g2_nor2_2 _0709_ (.A(_0167_),
    .B(_0183_),
    .Y(_0184_));
 sg13g2_nand2_2 _0710_ (.Y(_0185_),
    .A(net147),
    .B(_0184_));
 sg13g2_nor4_2 _0711_ (.A(_0111_),
    .B(\counter[4] ),
    .C(\counter[5] ),
    .Y(_0186_),
    .D(_0154_));
 sg13g2_inv_1 _0712_ (.Y(_0187_),
    .A(_0186_));
 sg13g2_nand3_1 _0713_ (.B(net145),
    .C(_0153_),
    .A(net158),
    .Y(_0188_));
 sg13g2_and4_1 _0714_ (.A(_0182_),
    .B(_0185_),
    .C(_0187_),
    .D(_0188_),
    .X(_0189_));
 sg13g2_a22oi_1 _0715_ (.Y(_0190_),
    .B1(_0171_),
    .B2(net145),
    .A2(_0169_),
    .A1(net147));
 sg13g2_and2_1 _0716_ (.A(net146),
    .B(_0159_),
    .X(_0191_));
 sg13g2_nand2_1 _0717_ (.Y(_0192_),
    .A(net146),
    .B(_0159_));
 sg13g2_nor3_1 _0718_ (.A(net158),
    .B(net160),
    .C(_0183_),
    .Y(_0193_));
 sg13g2_nand3_1 _0719_ (.B(net162),
    .C(_0157_),
    .A(net164),
    .Y(_0194_));
 sg13g2_nand2_1 _0720_ (.Y(_0195_),
    .A(net146),
    .B(_0193_));
 sg13g2_nand3_1 _0721_ (.B(net147),
    .C(_0157_),
    .A(net164),
    .Y(_0196_));
 sg13g2_nand2_1 _0722_ (.Y(_0197_),
    .A(net145),
    .B(_0193_));
 sg13g2_nand4_1 _0723_ (.B(_0190_),
    .C(_0196_),
    .A(_0189_),
    .Y(_0198_),
    .D(_0197_));
 sg13g2_nor4_1 _0724_ (.A(_0174_),
    .B(_0175_),
    .C(_0176_),
    .D(_0198_),
    .Y(_0199_));
 sg13g2_nor2_2 _0725_ (.A(\state[3] ),
    .B(\state[2] ),
    .Y(_0200_));
 sg13g2_and2_1 _0726_ (.A(net166),
    .B(_0200_),
    .X(_0201_));
 sg13g2_nor2b_1 _0727_ (.A(_0181_),
    .B_N(_0200_),
    .Y(_0202_));
 sg13g2_nor2_2 _0728_ (.A(\state[0] ),
    .B(net168),
    .Y(_0203_));
 sg13g2_a21oi_1 _0729_ (.A1(_0180_),
    .A2(_0203_),
    .Y(_0204_),
    .B1(_0202_));
 sg13g2_nor2b_2 _0730_ (.A(\state[0] ),
    .B_N(\state[1] ),
    .Y(_0205_));
 sg13g2_nand2b_1 _0731_ (.Y(_0206_),
    .B(net168),
    .A_N(net169));
 sg13g2_nand2_2 _0732_ (.Y(_0207_),
    .A(net167),
    .B(_0200_));
 sg13g2_o21ai_1 _0733_ (.B1(_0204_),
    .Y(_0208_),
    .A1(_0206_),
    .A2(_0207_));
 sg13g2_nor2b_2 _0734_ (.A(net168),
    .B_N(net169),
    .Y(_0209_));
 sg13g2_nand2b_1 _0735_ (.Y(_0210_),
    .B(net169),
    .A_N(net168));
 sg13g2_nor2b_2 _0736_ (.A(\state[3] ),
    .B_N(\state[2] ),
    .Y(_0211_));
 sg13g2_and3_1 _0737_ (.X(_0212_),
    .A(net167),
    .B(_0209_),
    .C(_0211_));
 sg13g2_nand3_1 _0738_ (.B(_0209_),
    .C(_0211_),
    .A(net167),
    .Y(_0213_));
 sg13g2_nor2_1 _0739_ (.A(_0182_),
    .B(_0212_),
    .Y(_0214_));
 sg13g2_nand2b_1 _0740_ (.Y(_0215_),
    .B(_0213_),
    .A_N(_0182_));
 sg13g2_nand2_2 _0741_ (.Y(_0216_),
    .A(\state[3] ),
    .B(\state[2] ));
 sg13g2_nor3_1 _0742_ (.A(net167),
    .B(_0210_),
    .C(_0216_),
    .Y(_0217_));
 sg13g2_nor3_1 _0743_ (.A(_0208_),
    .B(_0215_),
    .C(_0217_),
    .Y(_0218_));
 sg13g2_nor2_1 _0744_ (.A(\spi.done ),
    .B(_0214_),
    .Y(_0219_));
 sg13g2_a21oi_1 _0745_ (.A1(_0111_),
    .A2(_0014_),
    .Y(_0220_),
    .B1(_0155_));
 sg13g2_nor4_1 _0746_ (.A(_0116_),
    .B(_0014_),
    .C(_0155_),
    .D(_0213_),
    .Y(_0221_));
 sg13g2_nor4_2 _0747_ (.A(_0199_),
    .B(_0218_),
    .C(_0219_),
    .Y(_0222_),
    .D(_0221_));
 sg13g2_nor3_1 _0748_ (.A(_0177_),
    .B(_0208_),
    .C(_0212_),
    .Y(_0223_));
 sg13g2_nand4_1 _0749_ (.B(\state[2] ),
    .C(_0012_),
    .A(\state[3] ),
    .Y(_0224_),
    .D(_0209_));
 sg13g2_o21ai_1 _0750_ (.B1(_0224_),
    .Y(_0225_),
    .A1(_0213_),
    .A2(_0220_));
 sg13g2_nor2_1 _0751_ (.A(_0223_),
    .B(_0225_),
    .Y(_0226_));
 sg13g2_mux2_1 _0752_ (.A0(net61),
    .A1(_0226_),
    .S(_0222_),
    .X(_0045_));
 sg13g2_nand2_2 _0753_ (.Y(_0227_),
    .A(_0201_),
    .B(_0209_));
 sg13g2_nand2_2 _0754_ (.Y(_0228_),
    .A(net166),
    .B(_0205_));
 sg13g2_nand2_1 _0755_ (.Y(_0229_),
    .A(_0201_),
    .B(_0205_));
 sg13g2_and2_1 _0756_ (.A(\timer[1] ),
    .B(\timer[0] ),
    .X(_0230_));
 sg13g2_nor2_2 _0757_ (.A(_0149_),
    .B(_0183_),
    .Y(_0231_));
 sg13g2_and2_1 _0758_ (.A(\counter[4] ),
    .B(_0231_),
    .X(_0232_));
 sg13g2_nand3_1 _0759_ (.B(\counter[6] ),
    .C(_0232_),
    .A(\counter[5] ),
    .Y(_0233_));
 sg13g2_nand3_1 _0760_ (.B(net97),
    .C(\counter[14] ),
    .A(\counter[13] ),
    .Y(_0234_));
 sg13g2_and2_2 _0761_ (.A(net157),
    .B(net156),
    .X(_0235_));
 sg13g2_nand4_1 _0762_ (.B(net156),
    .C(net155),
    .A(\counter[7] ),
    .Y(_0236_),
    .D(net153));
 sg13g2_nand4_1 _0763_ (.B(net153),
    .C(net151),
    .A(net154),
    .Y(_0237_),
    .D(_0235_));
 sg13g2_nor4_2 _0764_ (.A(\counter[15] ),
    .B(_0233_),
    .C(_0234_),
    .Y(_0238_),
    .D(_0237_));
 sg13g2_nor4_2 _0765_ (.A(net101),
    .B(_0233_),
    .C(_0234_),
    .Y(_0239_),
    .D(_0237_));
 sg13g2_nand4_1 _0766_ (.B(\timer[3] ),
    .C(_0230_),
    .A(\timer[2] ),
    .Y(_0240_),
    .D(_0239_));
 sg13g2_nor2_1 _0767_ (.A(_0233_),
    .B(_0236_),
    .Y(_0241_));
 sg13g2_o21ai_1 _0768_ (.B1(net57),
    .Y(_0242_),
    .A1(_0229_),
    .A2(_0240_));
 sg13g2_nand2_1 _0769_ (.Y(_0046_),
    .A(_0227_),
    .B(net58));
 sg13g2_and2_1 _0770_ (.A(_0203_),
    .B(_0211_),
    .X(_0243_));
 sg13g2_a22oi_1 _0771_ (.Y(_0244_),
    .B1(_0243_),
    .B2(net166),
    .A2(_0205_),
    .A1(_0180_));
 sg13g2_nand2_1 _0772_ (.Y(_0245_),
    .A(net167),
    .B(_0243_));
 sg13g2_and2_1 _0773_ (.A(_0244_),
    .B(_0245_),
    .X(_0246_));
 sg13g2_o21ai_1 _0774_ (.B1(_0246_),
    .Y(_0247_),
    .A1(_0181_),
    .A2(_0216_));
 sg13g2_mux2_1 _0775_ (.A0(net108),
    .A1(\spi.done ),
    .S(_0247_),
    .X(_0248_));
 sg13g2_nand3_1 _0776_ (.B(_0209_),
    .C(_0211_),
    .A(net166),
    .Y(_0249_));
 sg13g2_nor3_2 _0777_ (.A(net169),
    .B(net168),
    .C(_0207_),
    .Y(_0250_));
 sg13g2_nor2_2 _0778_ (.A(_0215_),
    .B(_0250_),
    .Y(_0251_));
 sg13g2_and3_1 _0779_ (.X(_0047_),
    .A(_0248_),
    .B(_0249_),
    .C(_0251_));
 sg13g2_a221oi_1 _0780_ (.B2(net160),
    .C1(_0213_),
    .B1(_0153_),
    .A1(net164),
    .Y(_0252_),
    .A2(_0014_));
 sg13g2_nor2_1 _0781_ (.A(\spi.done ),
    .B(_0249_),
    .Y(_0253_));
 sg13g2_nor3_1 _0782_ (.A(_0219_),
    .B(_0252_),
    .C(_0253_),
    .Y(_0254_));
 sg13g2_nand3_1 _0783_ (.B(_0200_),
    .C(_0209_),
    .A(net167),
    .Y(_0255_));
 sg13g2_nand3b_1 _0784_ (.B(_0205_),
    .C(net167),
    .Y(_0256_),
    .A_N(\state[3] ));
 sg13g2_nand3_1 _0785_ (.B(_0205_),
    .C(_0211_),
    .A(\state[4] ),
    .Y(_0257_));
 sg13g2_nand4_1 _0786_ (.B(_0249_),
    .C(_0255_),
    .A(_0214_),
    .Y(_0258_),
    .D(_0257_));
 sg13g2_nand3_1 _0787_ (.B(_0254_),
    .C(_0258_),
    .A(_0198_),
    .Y(_0259_));
 sg13g2_nand2_1 _0788_ (.Y(_0260_),
    .A(net54),
    .B(_0259_));
 sg13g2_nor2_1 _0789_ (.A(_0178_),
    .B(_0207_),
    .Y(_0261_));
 sg13g2_or2_2 _0790_ (.X(_0262_),
    .B(_0207_),
    .A(_0178_));
 sg13g2_nand3_1 _0791_ (.B(_0260_),
    .C(_0262_),
    .A(net83),
    .Y(_0048_));
 sg13g2_nor2_1 _0792_ (.A(_0154_),
    .B(_0183_),
    .Y(_0263_));
 sg13g2_nor2_2 _0793_ (.A(net165),
    .B(_0167_),
    .Y(_0264_));
 sg13g2_a21oi_1 _0794_ (.A1(net162),
    .A2(_0264_),
    .Y(_0265_),
    .B1(_0263_));
 sg13g2_nand2b_2 _0795_ (.Y(_0266_),
    .B(net145),
    .A_N(_0265_));
 sg13g2_nor2_1 _0796_ (.A(_0112_),
    .B(_0187_),
    .Y(_0267_));
 sg13g2_a21oi_1 _0797_ (.A1(net145),
    .A2(_0168_),
    .Y(_0268_),
    .B1(_0267_));
 sg13g2_nand2_1 _0798_ (.Y(_0269_),
    .A(_0266_),
    .B(_0268_));
 sg13g2_nor3_2 _0799_ (.A(_0176_),
    .B(_0191_),
    .C(_0269_),
    .Y(_0270_));
 sg13g2_and2_1 _0800_ (.A(_0151_),
    .B(_0197_),
    .X(_0271_));
 sg13g2_and2_1 _0801_ (.A(_0195_),
    .B(_0271_),
    .X(_0272_));
 sg13g2_nand3_1 _0802_ (.B(_0165_),
    .C(_0272_),
    .A(_0161_),
    .Y(_0273_));
 sg13g2_nor2_2 _0803_ (.A(net162),
    .B(_0154_),
    .Y(_0274_));
 sg13g2_a21oi_2 _0804_ (.B1(_0170_),
    .Y(_0275_),
    .A2(_0274_),
    .A1(net147));
 sg13g2_inv_1 _0805_ (.Y(_0276_),
    .A(_0275_));
 sg13g2_o21ai_1 _0806_ (.B1(net147),
    .Y(_0277_),
    .A1(_0231_),
    .A2(_0264_));
 sg13g2_nand2_1 _0807_ (.Y(_0278_),
    .A(net158),
    .B(_0155_));
 sg13g2_nand2_1 _0808_ (.Y(_0279_),
    .A(net160),
    .B(_0175_));
 sg13g2_nand2_1 _0809_ (.Y(_0280_),
    .A(_0185_),
    .B(_0279_));
 sg13g2_nand2_1 _0810_ (.Y(_0281_),
    .A(_0275_),
    .B(_0277_));
 sg13g2_nand2_1 _0811_ (.Y(_0282_),
    .A(net146),
    .B(_0168_));
 sg13g2_a21o_1 _0812_ (.A2(_0274_),
    .A1(net164),
    .B1(_0184_),
    .X(_0283_));
 sg13g2_o21ai_1 _0813_ (.B1(_0152_),
    .Y(_0284_),
    .A1(_0163_),
    .A2(_0283_));
 sg13g2_nand4_1 _0814_ (.B(_0190_),
    .C(_0282_),
    .A(_0188_),
    .Y(_0285_),
    .D(_0284_));
 sg13g2_nor4_2 _0815_ (.A(_0273_),
    .B(_0280_),
    .C(_0281_),
    .Y(_0286_),
    .D(_0285_));
 sg13g2_and2_1 _0816_ (.A(_0270_),
    .B(_0286_),
    .X(_0287_));
 sg13g2_nand2_1 _0817_ (.Y(_0288_),
    .A(_0270_),
    .B(_0286_));
 sg13g2_nor2_2 _0818_ (.A(_0179_),
    .B(_0210_),
    .Y(_0289_));
 sg13g2_nand2_2 _0819_ (.Y(_0290_),
    .A(_0180_),
    .B(_0209_));
 sg13g2_nand2b_1 _0820_ (.Y(_0291_),
    .B(_0289_),
    .A_N(_0174_));
 sg13g2_and2_1 _0821_ (.A(_0195_),
    .B(_0261_),
    .X(_0292_));
 sg13g2_and3_1 _0822_ (.X(_0293_),
    .A(_0166_),
    .B(_0192_),
    .C(_0292_));
 sg13g2_nor2_2 _0823_ (.A(_0216_),
    .B(_0228_),
    .Y(_0294_));
 sg13g2_or2_1 _0824_ (.X(_0295_),
    .B(_0228_),
    .A(_0216_));
 sg13g2_nor4_1 _0825_ (.A(_0202_),
    .B(_0261_),
    .C(_0289_),
    .D(_0294_),
    .Y(_0296_));
 sg13g2_nor4_1 _0826_ (.A(\inval[4] ),
    .B(\inval[5] ),
    .C(\inval[6] ),
    .D(\inval[7] ),
    .Y(_0297_));
 sg13g2_nor4_1 _0827_ (.A(\inval[0] ),
    .B(\inval[1] ),
    .C(\inval[2] ),
    .D(\inval[3] ),
    .Y(_0298_));
 sg13g2_and2_1 _0828_ (.A(_0297_),
    .B(_0298_),
    .X(_0299_));
 sg13g2_a221oi_1 _0829_ (.B2(_0299_),
    .C1(_0296_),
    .B1(_0294_),
    .A1(_0172_),
    .Y(_0300_),
    .A2(_0293_));
 sg13g2_o21ai_1 _0830_ (.B1(_0300_),
    .Y(_0301_),
    .A1(_0288_),
    .A2(_0291_));
 sg13g2_nand2_1 _0831_ (.Y(_0302_),
    .A(net56),
    .B(net140));
 sg13g2_nor3_1 _0832_ (.A(net167),
    .B(_0206_),
    .C(_0216_),
    .Y(_0303_));
 sg13g2_nor3_1 _0833_ (.A(_0261_),
    .B(_0289_),
    .C(_0303_),
    .Y(_0304_));
 sg13g2_or2_2 _0834_ (.X(_0305_),
    .B(_0304_),
    .A(net140));
 sg13g2_or2_1 _0835_ (.X(_0306_),
    .B(_0231_),
    .A(_0171_));
 sg13g2_or2_1 _0836_ (.X(_0307_),
    .B(_0019_),
    .A(net151));
 sg13g2_nor2b_2 _0837_ (.A(net154),
    .B_N(net153),
    .Y(_0308_));
 sg13g2_nand2b_1 _0838_ (.Y(_0309_),
    .B(\counter[10] ),
    .A_N(net155));
 sg13g2_nor2_1 _0839_ (.A(net157),
    .B(net156),
    .Y(_0310_));
 sg13g2_or2_1 _0840_ (.X(_0311_),
    .B(net156),
    .A(net157));
 sg13g2_nand3_1 _0841_ (.B(_0308_),
    .C(_0310_),
    .A(_0307_),
    .Y(_0312_));
 sg13g2_nor2b_1 _0842_ (.A(net157),
    .B_N(\counter[8] ),
    .Y(_0313_));
 sg13g2_nand3_1 _0843_ (.B(\counter[10] ),
    .C(_0019_),
    .A(net155),
    .Y(_0314_));
 sg13g2_nand4_1 _0844_ (.B(net153),
    .C(_0019_),
    .A(net154),
    .Y(_0315_),
    .D(_0313_));
 sg13g2_nor2_1 _0845_ (.A(net154),
    .B(net153),
    .Y(_0316_));
 sg13g2_nand3_1 _0846_ (.B(_0313_),
    .C(_0316_),
    .A(net152),
    .Y(_0317_));
 sg13g2_nand4_1 _0847_ (.B(_0163_),
    .C(_0315_),
    .A(net161),
    .Y(_0318_),
    .D(_0317_));
 sg13g2_a21oi_1 _0848_ (.A1(_0112_),
    .A2(_0264_),
    .Y(_0319_),
    .B1(_0263_));
 sg13g2_nand2_1 _0849_ (.Y(_0320_),
    .A(_0318_),
    .B(_0319_));
 sg13g2_nand3_1 _0850_ (.B(_0315_),
    .C(_0317_),
    .A(_0274_),
    .Y(_0321_));
 sg13g2_nor2b_1 _0851_ (.A(net153),
    .B_N(net154),
    .Y(_0322_));
 sg13g2_and2_1 _0852_ (.A(net151),
    .B(_0322_),
    .X(_0323_));
 sg13g2_nand3b_1 _0853_ (.B(net152),
    .C(net154),
    .Y(_0324_),
    .A_N(net153));
 sg13g2_a21o_1 _0854_ (.A2(_0324_),
    .A1(_0314_),
    .B1(_0311_),
    .X(_0325_));
 sg13g2_nand3_1 _0855_ (.B(_0264_),
    .C(_0325_),
    .A(net163),
    .Y(_0326_));
 sg13g2_nor2b_1 _0856_ (.A(net156),
    .B_N(net157),
    .Y(_0327_));
 sg13g2_nand2b_1 _0857_ (.Y(_0328_),
    .B(net157),
    .A_N(\counter[8] ));
 sg13g2_nor3_1 _0858_ (.A(net152),
    .B(_0309_),
    .C(_0328_),
    .Y(_0329_));
 sg13g2_nand3b_1 _0859_ (.B(_0308_),
    .C(_0327_),
    .Y(_0330_),
    .A_N(net151));
 sg13g2_and2_1 _0860_ (.A(_0126_),
    .B(_0322_),
    .X(_0331_));
 sg13g2_a221oi_1 _0861_ (.B2(_0235_),
    .C1(_0329_),
    .B1(_0331_),
    .A1(_0321_),
    .Y(_0332_),
    .A2(_0326_));
 sg13g2_nand3b_1 _0862_ (.B(_0235_),
    .C(_0308_),
    .Y(_0333_),
    .A_N(net151));
 sg13g2_o21ai_1 _0863_ (.B1(_0333_),
    .Y(_0334_),
    .A1(_0164_),
    .A2(_0169_));
 sg13g2_nand3_1 _0864_ (.B(_0235_),
    .C(_0308_),
    .A(_0019_),
    .Y(_0335_));
 sg13g2_nand3_1 _0865_ (.B(_0312_),
    .C(_0335_),
    .A(_0168_),
    .Y(_0336_));
 sg13g2_nand2_1 _0866_ (.Y(_0337_),
    .A(_0334_),
    .B(_0336_));
 sg13g2_nand2_1 _0867_ (.Y(_0338_),
    .A(_0323_),
    .B(_0327_));
 sg13g2_nor2b_1 _0868_ (.A(net151),
    .B_N(_0236_),
    .Y(_0339_));
 sg13g2_nand3b_1 _0869_ (.B(net151),
    .C(_0316_),
    .Y(_0340_),
    .A_N(\counter[8] ));
 sg13g2_a21oi_1 _0870_ (.A1(_0126_),
    .A2(_0340_),
    .Y(_0341_),
    .B1(_0339_));
 sg13g2_o21ai_1 _0871_ (.B1(_0194_),
    .Y(_0342_),
    .A1(_0278_),
    .A2(_0341_));
 sg13g2_o21ai_1 _0872_ (.B1(_0324_),
    .Y(_0343_),
    .A1(net152),
    .A2(_0309_));
 sg13g2_nand2_1 _0873_ (.Y(_0344_),
    .A(_0313_),
    .B(_0343_));
 sg13g2_o21ai_1 _0874_ (.B1(_0325_),
    .Y(_0345_),
    .A1(_0150_),
    .A2(_0159_));
 sg13g2_and2_1 _0875_ (.A(_0235_),
    .B(_0323_),
    .X(_0346_));
 sg13g2_nand4_1 _0876_ (.B(_0315_),
    .C(_0317_),
    .A(_0184_),
    .Y(_0347_),
    .D(_0330_));
 sg13g2_o21ai_1 _0877_ (.B1(_0345_),
    .Y(_0348_),
    .A1(_0346_),
    .A2(_0347_));
 sg13g2_nor2_1 _0878_ (.A(_0314_),
    .B(_0328_),
    .Y(_0349_));
 sg13g2_nand3_1 _0879_ (.B(_0235_),
    .C(_0316_),
    .A(net151),
    .Y(_0350_));
 sg13g2_nor2b_1 _0880_ (.A(_0349_),
    .B_N(_0350_),
    .Y(_0351_));
 sg13g2_a221oi_1 _0881_ (.B2(_0344_),
    .C1(_0306_),
    .B1(_0342_),
    .A1(_0312_),
    .Y(_0352_),
    .A2(_0320_));
 sg13g2_a221oi_1 _0882_ (.B2(_0351_),
    .C1(_0332_),
    .B1(_0348_),
    .A1(_0337_),
    .Y(_0353_),
    .A2(_0338_));
 sg13g2_nand3_1 _0883_ (.B(_0317_),
    .C(_0340_),
    .A(_0126_),
    .Y(_0354_));
 sg13g2_nand2_1 _0884_ (.Y(_0355_),
    .A(_0315_),
    .B(_0339_));
 sg13g2_and2_1 _0885_ (.A(_0306_),
    .B(_0355_),
    .X(_0356_));
 sg13g2_a221oi_1 _0886_ (.B2(_0356_),
    .C1(\inval[6] ),
    .B1(_0354_),
    .A1(_0352_),
    .Y(_0357_),
    .A2(_0353_));
 sg13g2_o21ai_1 _0887_ (.B1(\inval[6] ),
    .Y(_0358_),
    .A1(net161),
    .A2(net156));
 sg13g2_a21oi_1 _0888_ (.A1(net161),
    .A2(net156),
    .Y(_0359_),
    .B1(_0358_));
 sg13g2_or2_1 _0889_ (.X(_0360_),
    .B(_0359_),
    .A(\inval[5] ));
 sg13g2_xnor2_1 _0890_ (.Y(_0361_),
    .A(net163),
    .B(net157));
 sg13g2_a21oi_1 _0891_ (.A1(\inval[5] ),
    .A2(_0361_),
    .Y(_0362_),
    .B1(\inval[4] ));
 sg13g2_o21ai_1 _0892_ (.B1(_0362_),
    .Y(_0363_),
    .A1(_0357_),
    .A2(_0360_));
 sg13g2_a21oi_1 _0893_ (.A1(_0111_),
    .A2(_0113_),
    .Y(_0364_),
    .B1(_0122_));
 sg13g2_o21ai_1 _0894_ (.B1(_0364_),
    .Y(_0365_),
    .A1(_0111_),
    .A2(_0113_));
 sg13g2_a21oi_1 _0895_ (.A1(_0363_),
    .A2(_0365_),
    .Y(_0366_),
    .B1(\inval[3] ));
 sg13g2_o21ai_1 _0896_ (.B1(_0119_),
    .Y(_0367_),
    .A1(_0121_),
    .A2(_0017_));
 sg13g2_a21oi_1 _0897_ (.A1(\inval[2] ),
    .A2(_0018_),
    .Y(_0368_),
    .B1(\inval[1] ));
 sg13g2_o21ai_1 _0898_ (.B1(_0368_),
    .Y(_0369_),
    .A1(_0366_),
    .A2(_0367_));
 sg13g2_a21oi_2 _0899_ (.B1(_0295_),
    .Y(_0370_),
    .A2(_0369_),
    .A1(_0118_));
 sg13g2_nand4_1 _0900_ (.B(_0270_),
    .C(_0272_),
    .A(_0160_),
    .Y(_0371_),
    .D(_0282_));
 sg13g2_o21ai_1 _0901_ (.B1(_0289_),
    .Y(_0372_),
    .A1(_0287_),
    .A2(_0371_));
 sg13g2_o21ai_1 _0902_ (.B1(_0372_),
    .Y(_0373_),
    .A1(_0162_),
    .A2(_0262_));
 sg13g2_nor2_1 _0903_ (.A(_0370_),
    .B(_0373_),
    .Y(_0374_));
 sg13g2_o21ai_1 _0904_ (.B1(_0302_),
    .Y(_0049_),
    .A1(_0305_),
    .A2(_0374_));
 sg13g2_nor4_1 _0905_ (.A(_0176_),
    .B(_0186_),
    .C(_0191_),
    .D(_0280_),
    .Y(_0375_));
 sg13g2_a21oi_1 _0906_ (.A1(_0271_),
    .A2(_0375_),
    .Y(_0376_),
    .B1(_0290_));
 sg13g2_nor4_1 _0907_ (.A(_0293_),
    .B(_0305_),
    .C(_0370_),
    .D(_0376_),
    .Y(_0377_));
 sg13g2_a21oi_1 _0908_ (.A1(_0106_),
    .A2(net140),
    .Y(_0050_),
    .B1(_0377_));
 sg13g2_nor2_1 _0909_ (.A(_0192_),
    .B(_0262_),
    .Y(_0378_));
 sg13g2_nor4_1 _0910_ (.A(_0175_),
    .B(_0267_),
    .C(_0273_),
    .D(_0276_),
    .Y(_0379_));
 sg13g2_nor2_1 _0911_ (.A(_0290_),
    .B(_0379_),
    .Y(_0380_));
 sg13g2_nor3_1 _0912_ (.A(_0370_),
    .B(_0378_),
    .C(_0380_),
    .Y(_0381_));
 sg13g2_nand2_1 _0913_ (.Y(_0382_),
    .A(net53),
    .B(_0301_));
 sg13g2_o21ai_1 _0914_ (.B1(_0382_),
    .Y(_0051_),
    .A1(_0305_),
    .A2(_0381_));
 sg13g2_nand4_1 _0915_ (.B(_0266_),
    .C(_0271_),
    .A(_0166_),
    .Y(_0383_),
    .D(_0279_));
 sg13g2_a21oi_1 _0916_ (.A1(_0289_),
    .A2(_0383_),
    .Y(_0384_),
    .B1(_0370_));
 sg13g2_nand2_1 _0917_ (.Y(_0385_),
    .A(net51),
    .B(net140));
 sg13g2_o21ai_1 _0918_ (.B1(_0385_),
    .Y(_0052_),
    .A1(_0305_),
    .A2(_0384_));
 sg13g2_nand4_1 _0919_ (.B(_0185_),
    .C(_0187_),
    .A(_0165_),
    .Y(_0386_),
    .D(_0266_));
 sg13g2_o21ai_1 _0920_ (.B1(_0289_),
    .Y(_0387_),
    .A1(_0287_),
    .A2(_0386_));
 sg13g2_o21ai_1 _0921_ (.B1(_0387_),
    .Y(_0388_),
    .A1(_0196_),
    .A2(_0262_));
 sg13g2_nor3_1 _0922_ (.A(_0305_),
    .B(_0370_),
    .C(_0388_),
    .Y(_0389_));
 sg13g2_a21oi_1 _0923_ (.A1(_0105_),
    .A2(net140),
    .Y(_0053_),
    .B1(_0389_));
 sg13g2_nor2_1 _0924_ (.A(_0266_),
    .B(_0290_),
    .Y(_0390_));
 sg13g2_nand3_1 _0925_ (.B(_0185_),
    .C(_0275_),
    .A(_0165_),
    .Y(_0391_));
 sg13g2_a221oi_1 _0926_ (.B2(_0289_),
    .C1(_0390_),
    .B1(_0391_),
    .A1(_0162_),
    .Y(_0392_),
    .A2(_0292_));
 sg13g2_nor2b_1 _0927_ (.A(_0370_),
    .B_N(_0392_),
    .Y(_0393_));
 sg13g2_nand2_1 _0928_ (.Y(_0394_),
    .A(net52),
    .B(net140));
 sg13g2_o21ai_1 _0929_ (.B1(_0394_),
    .Y(_0054_),
    .A1(_0305_),
    .A2(_0393_));
 sg13g2_and4_1 _0930_ (.A(_0151_),
    .B(_0161_),
    .C(_0266_),
    .D(_0279_),
    .X(_0395_));
 sg13g2_a21oi_1 _0931_ (.A1(_0282_),
    .A2(_0395_),
    .Y(_0396_),
    .B1(_0290_));
 sg13g2_nor3_1 _0932_ (.A(_0370_),
    .B(_0378_),
    .C(_0396_),
    .Y(_0397_));
 sg13g2_nand2_1 _0933_ (.Y(_0398_),
    .A(net49),
    .B(net140));
 sg13g2_o21ai_1 _0934_ (.B1(_0398_),
    .Y(_0055_),
    .A1(_0305_),
    .A2(_0397_));
 sg13g2_nor3_1 _0935_ (.A(_0370_),
    .B(_0378_),
    .C(_0390_),
    .Y(_0399_));
 sg13g2_nand2_1 _0936_ (.Y(_0400_),
    .A(net50),
    .B(net140));
 sg13g2_o21ai_1 _0937_ (.B1(_0400_),
    .Y(_0056_),
    .A1(_0305_),
    .A2(_0399_));
 sg13g2_nand2b_1 _0938_ (.Y(_0401_),
    .B(_0211_),
    .A_N(_0181_));
 sg13g2_nand2_2 _0939_ (.Y(_0402_),
    .A(_0229_),
    .B(_0401_));
 sg13g2_xnor2_1 _0940_ (.Y(_0403_),
    .A(\inval[1] ),
    .B(\inbuf[1] ));
 sg13g2_xnor2_1 _0941_ (.Y(_0404_),
    .A(\inval[6] ),
    .B(\inbuf[6] ));
 sg13g2_xnor2_1 _0942_ (.Y(_0405_),
    .A(\inval[3] ),
    .B(\inbuf[3] ));
 sg13g2_xnor2_1 _0943_ (.Y(_0406_),
    .A(\inval[5] ),
    .B(\inbuf[5] ));
 sg13g2_xnor2_1 _0944_ (.Y(_0407_),
    .A(\inval[7] ),
    .B(\inbuf[7] ));
 sg13g2_a22oi_1 _0945_ (.Y(_0408_),
    .B1(_0122_),
    .B2(\inbuf[4] ),
    .A2(_0120_),
    .A1(\inval[2] ));
 sg13g2_xnor2_1 _0946_ (.Y(_0409_),
    .A(\inval[0] ),
    .B(\inbuf[0] ));
 sg13g2_nand4_1 _0947_ (.B(_0406_),
    .C(_0408_),
    .A(_0404_),
    .Y(_0410_),
    .D(_0409_));
 sg13g2_a22oi_1 _0948_ (.Y(_0411_),
    .B1(\inval[4] ),
    .B2(_0123_),
    .A2(\inbuf[2] ),
    .A1(_0119_));
 sg13g2_nand4_1 _0949_ (.B(_0405_),
    .C(_0407_),
    .A(_0403_),
    .Y(_0412_),
    .D(_0411_));
 sg13g2_nor4_1 _0950_ (.A(\inbuf[4] ),
    .B(\inbuf[5] ),
    .C(\inbuf[6] ),
    .D(\inbuf[7] ),
    .Y(_0413_));
 sg13g2_nor4_1 _0951_ (.A(\inbuf[0] ),
    .B(\inbuf[1] ),
    .C(\inbuf[2] ),
    .D(\inbuf[3] ),
    .Y(_0414_));
 sg13g2_nand2_1 _0952_ (.Y(_0415_),
    .A(_0413_),
    .B(_0414_));
 sg13g2_o21ai_1 _0953_ (.B1(_0415_),
    .Y(_0416_),
    .A1(_0410_),
    .A2(_0412_));
 sg13g2_nand3_1 _0954_ (.B(_0203_),
    .C(_0416_),
    .A(_0201_),
    .Y(_0417_));
 sg13g2_nor2_2 _0955_ (.A(\spi.done ),
    .B(_0251_),
    .Y(_0418_));
 sg13g2_nand3_1 _0956_ (.B(_0205_),
    .C(_0211_),
    .A(net166),
    .Y(_0419_));
 sg13g2_nand2_1 _0957_ (.Y(_0420_),
    .A(_0257_),
    .B(_0419_));
 sg13g2_nor2_1 _0958_ (.A(_0253_),
    .B(_0418_),
    .Y(_0421_));
 sg13g2_o21ai_1 _0959_ (.B1(_0421_),
    .Y(_0422_),
    .A1(resetb),
    .A2(_0229_));
 sg13g2_a221oi_1 _0960_ (.B2(net9),
    .C1(_0422_),
    .B1(_0420_),
    .A1(\spi.done ),
    .Y(_0423_),
    .A2(_0247_));
 sg13g2_nand2_1 _0961_ (.Y(_0424_),
    .A(_0417_),
    .B(_0423_));
 sg13g2_a21oi_2 _0962_ (.B1(_0424_),
    .Y(_0425_),
    .A2(_0402_),
    .A1(_0240_));
 sg13g2_nor3_1 _0963_ (.A(\counter[12] ),
    .B(\counter[15] ),
    .C(\counter[14] ),
    .Y(_0426_));
 sg13g2_nand3_1 _0964_ (.B(_0114_),
    .C(_0426_),
    .A(_0113_),
    .Y(_0427_));
 sg13g2_nor4_2 _0965_ (.A(net155),
    .B(net153),
    .C(net152),
    .Y(_0428_),
    .D(_0311_));
 sg13g2_nand2b_2 _0966_ (.Y(_0429_),
    .B(_0428_),
    .A_N(_0427_));
 sg13g2_nor2_1 _0967_ (.A(_0195_),
    .B(_0429_),
    .Y(_0430_));
 sg13g2_o21ai_1 _0968_ (.B1(_0212_),
    .Y(_0431_),
    .A1(_0162_),
    .A2(_0429_));
 sg13g2_nor2_1 _0969_ (.A(_0430_),
    .B(_0431_),
    .Y(_0432_));
 sg13g2_nand2_1 _0970_ (.Y(_0433_),
    .A(_0152_),
    .B(_0231_));
 sg13g2_a21oi_1 _0971_ (.A1(\state[3] ),
    .A2(_0115_),
    .Y(_0434_),
    .B1(_0228_));
 sg13g2_nand3_1 _0972_ (.B(net166),
    .C(_0203_),
    .A(_0115_),
    .Y(_0435_));
 sg13g2_nand2_1 _0973_ (.Y(_0436_),
    .A(_0256_),
    .B(_0435_));
 sg13g2_or3_2 _0974_ (.A(_0237_),
    .B(_0427_),
    .C(_0433_),
    .X(_0437_));
 sg13g2_nor4_2 _0975_ (.A(net169),
    .B(net168),
    .C(_0207_),
    .Y(_0438_),
    .D(_0437_));
 sg13g2_or2_1 _0976_ (.X(_0439_),
    .B(_0438_),
    .A(_0432_));
 sg13g2_nor4_1 _0977_ (.A(_0182_),
    .B(_0434_),
    .C(_0436_),
    .D(_0439_),
    .Y(_0440_));
 sg13g2_nand2_1 _0978_ (.Y(_0441_),
    .A(_0246_),
    .B(_0440_));
 sg13g2_mux2_1 _0979_ (.A0(net169),
    .A1(_0441_),
    .S(_0425_),
    .X(_0057_));
 sg13g2_nand2_1 _0980_ (.Y(_0442_),
    .A(_0256_),
    .B(_0431_));
 sg13g2_a21oi_2 _0981_ (.B1(_0294_),
    .Y(_0443_),
    .A2(_0437_),
    .A1(_0250_));
 sg13g2_nand3_1 _0982_ (.B(_0249_),
    .C(_0419_),
    .A(_0224_),
    .Y(_0444_));
 sg13g2_o21ai_1 _0983_ (.B1(_0290_),
    .Y(_0445_),
    .A1(\state[2] ),
    .A2(_0228_));
 sg13g2_nand2_1 _0984_ (.Y(_0446_),
    .A(_0227_),
    .B(_0255_));
 sg13g2_nor3_1 _0985_ (.A(_0444_),
    .B(_0445_),
    .C(_0446_),
    .Y(_0447_));
 sg13g2_nand4_1 _0986_ (.B(_0431_),
    .C(_0443_),
    .A(_0256_),
    .Y(_0448_),
    .D(_0447_));
 sg13g2_mux2_1 _0987_ (.A0(net168),
    .A1(_0448_),
    .S(_0425_),
    .X(_0058_));
 sg13g2_nand2_1 _0988_ (.Y(_0449_),
    .A(_0245_),
    .B(_0262_));
 sg13g2_a21o_1 _0989_ (.A2(_0243_),
    .A1(net166),
    .B1(_0202_),
    .X(_0450_));
 sg13g2_nor2_1 _0990_ (.A(_0195_),
    .B(_0213_),
    .Y(_0451_));
 sg13g2_a21oi_1 _0991_ (.A1(_0170_),
    .A2(_0182_),
    .Y(_0452_),
    .B1(_0451_));
 sg13g2_nor2_1 _0992_ (.A(_0429_),
    .B(_0452_),
    .Y(_0453_));
 sg13g2_nor4_1 _0993_ (.A(_0444_),
    .B(_0449_),
    .C(_0450_),
    .D(_0453_),
    .Y(_0454_));
 sg13g2_nand2_1 _0994_ (.Y(_0455_),
    .A(_0443_),
    .B(_0454_));
 sg13g2_nand2_1 _0995_ (.Y(_0456_),
    .A(_0425_),
    .B(_0455_));
 sg13g2_o21ai_1 _0996_ (.B1(_0456_),
    .Y(_0059_),
    .A1(_0115_),
    .A2(_0425_));
 sg13g2_nand4_1 _0997_ (.B(_0224_),
    .C(_0401_),
    .A(_0179_),
    .Y(_0457_),
    .D(_0443_));
 sg13g2_mux2_1 _0998_ (.A0(net115),
    .A1(_0457_),
    .S(_0425_),
    .X(_0060_));
 sg13g2_o21ai_1 _0999_ (.B1(_0255_),
    .Y(_0458_),
    .A1(_0181_),
    .A2(_0216_));
 sg13g2_nor4_2 _1000_ (.A(_0438_),
    .B(_0442_),
    .C(_0449_),
    .Y(_0459_),
    .D(_0458_));
 sg13g2_nor2_1 _1001_ (.A(net89),
    .B(_0425_),
    .Y(_0460_));
 sg13g2_a21oi_1 _1002_ (.A1(_0425_),
    .A2(_0459_),
    .Y(_0061_),
    .B1(_0460_));
 sg13g2_nand2_2 _1003_ (.Y(_0461_),
    .A(_0204_),
    .B(_0227_));
 sg13g2_o21ai_1 _1004_ (.B1(_0224_),
    .Y(_0462_),
    .A1(_0206_),
    .A2(_0207_));
 sg13g2_nor2_2 _1005_ (.A(_0461_),
    .B(_0462_),
    .Y(_0463_));
 sg13g2_or2_2 _1006_ (.X(_0464_),
    .B(_0462_),
    .A(_0461_));
 sg13g2_nor3_1 _1007_ (.A(_0215_),
    .B(_0250_),
    .C(_0402_),
    .Y(_0465_));
 sg13g2_a21oi_2 _1008_ (.B1(_0418_),
    .Y(_0466_),
    .A2(_0465_),
    .A1(_0463_));
 sg13g2_a21o_1 _1009_ (.A2(_0465_),
    .A1(_0463_),
    .B1(_0418_),
    .X(_0467_));
 sg13g2_nand2_2 _1010_ (.Y(_0468_),
    .A(_0463_),
    .B(net141));
 sg13g2_a21oi_2 _1011_ (.B1(_0468_),
    .Y(_0469_),
    .A2(_0251_),
    .A1(_0239_));
 sg13g2_a22oi_1 _1012_ (.Y(_0470_),
    .B1(_0469_),
    .B2(net45),
    .A2(_0467_),
    .A1(net164));
 sg13g2_inv_1 _1013_ (.Y(_0062_),
    .A(net46));
 sg13g2_a21o_1 _1014_ (.A2(_0158_),
    .A1(_0148_),
    .B1(_0468_),
    .X(_0471_));
 sg13g2_o21ai_1 _1015_ (.B1(_0471_),
    .Y(_0063_),
    .A1(_0112_),
    .A2(net141));
 sg13g2_nand2b_1 _1016_ (.Y(_0472_),
    .B(net141),
    .A_N(_0183_));
 sg13g2_xor2_1 _1017_ (.B(_0472_),
    .A(net160),
    .X(_0473_));
 sg13g2_nor2_1 _1018_ (.A(_0464_),
    .B(_0473_),
    .Y(_0064_));
 sg13g2_nand2_2 _1019_ (.Y(_0474_),
    .A(_0238_),
    .B(_0402_));
 sg13g2_a21oi_1 _1020_ (.A1(_0239_),
    .A2(_0402_),
    .Y(_0475_),
    .B1(_0461_));
 sg13g2_nand2_1 _1021_ (.Y(_0476_),
    .A(_0463_),
    .B(_0474_));
 sg13g2_nor2_1 _1022_ (.A(net109),
    .B(_0472_),
    .Y(_0477_));
 sg13g2_xnor2_1 _1023_ (.Y(_0478_),
    .A(net159),
    .B(_0477_));
 sg13g2_nor2_1 _1024_ (.A(_0476_),
    .B(net110),
    .Y(_0065_));
 sg13g2_nand2b_1 _1025_ (.Y(_0479_),
    .B(_0463_),
    .A_N(_0232_));
 sg13g2_nand2_1 _1026_ (.Y(_0480_),
    .A(net141),
    .B(_0479_));
 sg13g2_a21oi_1 _1027_ (.A1(_0231_),
    .A2(net141),
    .Y(_0481_),
    .B1(net105));
 sg13g2_a21oi_1 _1028_ (.A1(net141),
    .A2(_0479_),
    .Y(_0066_),
    .B1(_0481_));
 sg13g2_nand2_1 _1029_ (.Y(_0482_),
    .A(net106),
    .B(_0480_));
 sg13g2_o21ai_1 _1030_ (.B1(_0482_),
    .Y(_0067_),
    .A1(_0433_),
    .A2(_0468_));
 sg13g2_nand3_1 _1031_ (.B(_0232_),
    .C(_0466_),
    .A(\counter[5] ),
    .Y(_0483_));
 sg13g2_nor2_1 _1032_ (.A(_0113_),
    .B(_0483_),
    .Y(_0484_));
 sg13g2_a21oi_1 _1033_ (.A1(_0113_),
    .A2(_0483_),
    .Y(_0485_),
    .B1(_0464_));
 sg13g2_nor2b_1 _1034_ (.A(_0484_),
    .B_N(net118),
    .Y(_0068_));
 sg13g2_xor2_1 _1035_ (.B(_0233_),
    .A(net92),
    .X(_0486_));
 sg13g2_a22oi_1 _1036_ (.Y(_0487_),
    .B1(_0469_),
    .B2(_0486_),
    .A2(_0467_),
    .A1(net157));
 sg13g2_inv_1 _1037_ (.Y(_0069_),
    .A(net93));
 sg13g2_nor2_1 _1038_ (.A(net156),
    .B(_0484_),
    .Y(_0488_));
 sg13g2_and2_1 _1039_ (.A(_0235_),
    .B(_0484_),
    .X(_0489_));
 sg13g2_nor4_1 _1040_ (.A(_0310_),
    .B(_0464_),
    .C(_0488_),
    .D(_0489_),
    .Y(_0070_));
 sg13g2_a21oi_1 _1041_ (.A1(net154),
    .A2(_0489_),
    .Y(_0490_),
    .B1(_0464_));
 sg13g2_o21ai_1 _1042_ (.B1(_0490_),
    .Y(_0491_),
    .A1(net154),
    .A2(_0489_));
 sg13g2_inv_1 _1043_ (.Y(_0071_),
    .A(_0491_));
 sg13g2_a21oi_1 _1044_ (.A1(net155),
    .A2(_0489_),
    .Y(_0492_),
    .B1(net72));
 sg13g2_a21oi_1 _1045_ (.A1(_0241_),
    .A2(net141),
    .Y(_0493_),
    .B1(_0464_));
 sg13g2_nor2b_1 _1046_ (.A(net73),
    .B_N(_0493_),
    .Y(_0072_));
 sg13g2_xnor2_1 _1047_ (.Y(_0494_),
    .A(_0019_),
    .B(_0241_));
 sg13g2_a22oi_1 _1048_ (.Y(_0495_),
    .B1(_0469_),
    .B2(_0494_),
    .A2(_0467_),
    .A1(net152));
 sg13g2_inv_1 _1049_ (.Y(_0073_),
    .A(net114));
 sg13g2_nor3_1 _1050_ (.A(_0113_),
    .B(_0237_),
    .C(_0483_),
    .Y(_0496_));
 sg13g2_nor2_1 _1051_ (.A(net97),
    .B(_0496_),
    .Y(_0497_));
 sg13g2_and2_1 _1052_ (.A(net97),
    .B(_0496_),
    .X(_0498_));
 sg13g2_nor3_1 _1053_ (.A(_0464_),
    .B(net98),
    .C(_0498_),
    .Y(_0074_));
 sg13g2_nor2_1 _1054_ (.A(net104),
    .B(_0498_),
    .Y(_0499_));
 sg13g2_and2_1 _1055_ (.A(net104),
    .B(_0498_),
    .X(_0500_));
 sg13g2_nor3_1 _1056_ (.A(_0464_),
    .B(_0499_),
    .C(_0500_),
    .Y(_0075_));
 sg13g2_or2_1 _1057_ (.X(_0501_),
    .B(_0500_),
    .A(net116));
 sg13g2_nand3_1 _1058_ (.B(net116),
    .C(_0498_),
    .A(net104),
    .Y(_0502_));
 sg13g2_and3_1 _1059_ (.X(_0076_),
    .A(_0463_),
    .B(_0501_),
    .C(_0502_));
 sg13g2_nand2_1 _1060_ (.Y(_0503_),
    .A(net101),
    .B(_0502_));
 sg13g2_nand2_1 _1061_ (.Y(_0504_),
    .A(_0239_),
    .B(net141));
 sg13g2_a21oi_1 _1062_ (.A1(net102),
    .A2(_0504_),
    .Y(_0077_),
    .B1(_0476_));
 sg13g2_nor2_1 _1063_ (.A(_0117_),
    .B(_0475_),
    .Y(_0505_));
 sg13g2_a21oi_1 _1064_ (.A1(_0117_),
    .A2(_0474_),
    .Y(_0078_),
    .B1(_0505_));
 sg13g2_nor2_1 _1065_ (.A(net90),
    .B(_0505_),
    .Y(_0506_));
 sg13g2_and2_1 _1066_ (.A(net90),
    .B(_0505_),
    .X(_0507_));
 sg13g2_nor3_1 _1067_ (.A(_0461_),
    .B(_0506_),
    .C(_0507_),
    .Y(_0079_));
 sg13g2_nor2_1 _1068_ (.A(net77),
    .B(_0507_),
    .Y(_0508_));
 sg13g2_and2_1 _1069_ (.A(net77),
    .B(_0507_),
    .X(_0509_));
 sg13g2_nor3_1 _1070_ (.A(_0461_),
    .B(net78),
    .C(_0509_),
    .Y(_0080_));
 sg13g2_xnor2_1 _1071_ (.Y(_0510_),
    .A(net75),
    .B(_0509_));
 sg13g2_nor2_1 _1072_ (.A(_0461_),
    .B(net76),
    .Y(_0081_));
 sg13g2_nor2b_2 _1073_ (.A(net144),
    .B_N(sck),
    .Y(_0511_));
 sg13g2_or2_2 _1074_ (.X(_0512_),
    .B(sck),
    .A(net144));
 sg13g2_nor2_1 _1075_ (.A(_0024_),
    .B(_0512_),
    .Y(_0513_));
 sg13g2_a221oi_1 _1076_ (.B2(_0511_),
    .C1(_0513_),
    .B1(\spi.treg[0] ),
    .A1(\spi.d_latched[0] ),
    .Y(_0082_),
    .A2(net143));
 sg13g2_nor2_1 _1077_ (.A(_0025_),
    .B(_0512_),
    .Y(_0514_));
 sg13g2_a221oi_1 _1078_ (.B2(_0511_),
    .C1(_0514_),
    .B1(\spi.treg[1] ),
    .A1(\spi.d_latched[1] ),
    .Y(_0083_),
    .A2(net143));
 sg13g2_nor2_1 _1079_ (.A(_0026_),
    .B(_0512_),
    .Y(_0515_));
 sg13g2_a221oi_1 _1080_ (.B2(_0511_),
    .C1(_0515_),
    .B1(\spi.treg[2] ),
    .A1(\spi.d_latched[2] ),
    .Y(_0084_),
    .A2(net143));
 sg13g2_nor2_1 _1081_ (.A(_0027_),
    .B(_0512_),
    .Y(_0516_));
 sg13g2_a221oi_1 _1082_ (.B2(_0511_),
    .C1(_0516_),
    .B1(\spi.treg[3] ),
    .A1(\spi.d_latched[3] ),
    .Y(_0085_),
    .A2(net143));
 sg13g2_nor2_1 _1083_ (.A(_0028_),
    .B(_0512_),
    .Y(_0517_));
 sg13g2_a221oi_1 _1084_ (.B2(_0511_),
    .C1(_0517_),
    .B1(\spi.treg[4] ),
    .A1(\spi.d_latched[4] ),
    .Y(_0086_),
    .A2(net144));
 sg13g2_nor2_1 _1085_ (.A(_0029_),
    .B(_0512_),
    .Y(_0518_));
 sg13g2_a221oi_1 _1086_ (.B2(_0511_),
    .C1(_0518_),
    .B1(\spi.treg[5] ),
    .A1(\spi.d_latched[5] ),
    .Y(_0087_),
    .A2(net143));
 sg13g2_nor2_1 _1087_ (.A(_0030_),
    .B(_0512_),
    .Y(_0519_));
 sg13g2_a221oi_1 _1088_ (.B2(_0511_),
    .C1(_0519_),
    .B1(\spi.treg[6] ),
    .A1(\spi.d_latched[6] ),
    .Y(_0088_),
    .A2(net143));
 sg13g2_nor2_1 _1089_ (.A(\spi.state[1] ),
    .B(\spi.state[3] ),
    .Y(_0520_));
 sg13g2_nor3_1 _1090_ (.A(\spi.state[0] ),
    .B(\spi.state[2] ),
    .C(_0520_),
    .Y(_0521_));
 sg13g2_a22oi_1 _1091_ (.Y(_0089_),
    .B1(_0521_),
    .B2(_0134_),
    .A2(_0135_),
    .A1(_0107_));
 sg13g2_nand2b_1 _1092_ (.Y(_0522_),
    .B(\spi.w_latched ),
    .A_N(\spi.d_latched[7] ));
 sg13g2_o21ai_1 _1093_ (.B1(_0522_),
    .Y(_0523_),
    .A1(mosi),
    .A2(_0512_));
 sg13g2_a21oi_1 _1094_ (.A1(_0125_),
    .A2(_0511_),
    .Y(_0090_),
    .B1(_0523_));
 sg13g2_nor3_1 _1095_ (.A(net144),
    .B(_0109_),
    .C(\spi.stream ),
    .Y(_0524_));
 sg13g2_nand2_1 _1096_ (.Y(_0525_),
    .A(\spi.state[3] ),
    .B(_0127_));
 sg13g2_nor2_1 _1097_ (.A(_0016_),
    .B(_0525_),
    .Y(_0526_));
 sg13g2_nor2_1 _1098_ (.A(\spi.state[0] ),
    .B(_0526_),
    .Y(_0527_));
 sg13g2_nand3_1 _1099_ (.B(_0109_),
    .C(_0525_),
    .A(_0032_),
    .Y(_0528_));
 sg13g2_o21ai_1 _1100_ (.B1(_0528_),
    .Y(_0091_),
    .A1(_0524_),
    .A2(_0527_));
 sg13g2_mux2_1 _1101_ (.A0(net148),
    .A1(net47),
    .S(_0138_),
    .X(_0092_));
 sg13g2_nand2b_1 _1102_ (.Y(_0529_),
    .B(\spi.done ),
    .A_N(\spi.stream ));
 sg13g2_and2_1 _1103_ (.A(net54),
    .B(_0529_),
    .X(_0093_));
 sg13g2_or3_1 _1104_ (.A(\spi.state[0] ),
    .B(_0110_),
    .C(\spi.state[2] ),
    .X(_0530_));
 sg13g2_and2_1 _1105_ (.A(_0135_),
    .B(_0530_),
    .X(_0531_));
 sg13g2_nand2_1 _1106_ (.Y(_0532_),
    .A(\spi.nbit[0] ),
    .B(_0531_));
 sg13g2_o21ai_1 _1107_ (.B1(_0532_),
    .Y(_0094_),
    .A1(\spi.nbit[0] ),
    .A2(_0530_));
 sg13g2_nand2_1 _1108_ (.Y(_0533_),
    .A(\spi.nbit[1] ),
    .B(_0531_));
 sg13g2_xnor2_1 _1109_ (.Y(_0534_),
    .A(\spi.nbit[0] ),
    .B(\spi.nbit[1] ));
 sg13g2_o21ai_1 _1110_ (.B1(_0533_),
    .Y(_0095_),
    .A1(_0530_),
    .A2(_0534_));
 sg13g2_and2_1 _1111_ (.A(_0013_),
    .B(_0133_),
    .X(_0535_));
 sg13g2_nor4_1 _1112_ (.A(\spi.state[0] ),
    .B(\spi.state[2] ),
    .C(_0134_),
    .D(_0535_),
    .Y(_0536_));
 sg13g2_a21o_1 _1113_ (.A2(_0531_),
    .A1(\spi.nbit[2] ),
    .B1(_0536_),
    .X(_0096_));
 sg13g2_inv_1 _1115__3 (.Y(net30),
    .A(clknet_1_1__leaf_clk));
 sg13g2_inv_1 _1116__4 (.Y(net31),
    .A(clknet_1_1__leaf_clk));
 sg13g2_inv_1 _1117__5 (.Y(net32),
    .A(clknet_1_1__leaf_clk));
 sg13g2_inv_1 _1118__6 (.Y(net33),
    .A(clknet_1_0__leaf_clk));
 sg13g2_inv_1 _1119__7 (.Y(net34),
    .A(clknet_1_1__leaf_clk));
 sg13g2_inv_1 _1120__8 (.Y(net35),
    .A(clknet_1_0__leaf_clk));
 sg13g2_inv_1 _1121__9 (.Y(net36),
    .A(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_dfrbp_1 _1122_ (.CLK(net150),
    .RESET_B(net175),
    .D(_0033_),
    .Q_N(\spi.state[0] ),
    .Q(_0020_));
 sg13g2_dfrbp_1 _1123_ (.CLK(net149),
    .RESET_B(net174),
    .D(\spi.state[2] ),
    .Q_N(_0580_),
    .Q(\spi.state[1] ));
 sg13g2_dfrbp_1 _1124_ (.CLK(net149),
    .RESET_B(net174),
    .D(_0001_),
    .Q_N(_0581_),
    .Q(\spi.state[2] ));
 sg13g2_dfrbp_1 _1125_ (.CLK(net149),
    .RESET_B(net175),
    .D(_0000_),
    .Q_N(_0579_),
    .Q(\spi.state[3] ));
 sg13g2_dfrbp_1 _1126_ (.CLK(net148),
    .RESET_B(net174),
    .D(_0043_),
    .Q_N(\spi.treg[0] ),
    .Q(_0021_));
 sg13g2_dfrbp_1 _1127_ (.CLK(net28),
    .RESET_B(net174),
    .D(_0044_),
    .Q_N(_0578_),
    .Q(\spi.w_latched ));
 sg13g2_dfrbp_1 _1128_ (.CLK(clknet_4_6_0_clk_regs),
    .RESET_B(net177),
    .D(_0045_),
    .Q_N(dcb),
    .Q(_0022_));
 sg13g2_dfrbp_1 _1129_ (.CLK(clknet_4_5_0_clk_regs),
    .RESET_B(net176),
    .D(_0046_),
    .Q_N(resetb),
    .Q(_0023_));
 sg13g2_dfrbp_1 _1130_ (.CLK(clknet_4_5_0_clk_regs),
    .RESET_B(net174),
    .D(_0047_),
    .Q_N(_0015_),
    .Q(\spi.reg_dat_we ));
 sg13g2_dfrbp_1 _1131_ (.CLK(clknet_4_6_0_clk_regs),
    .RESET_B(net176),
    .D(_0048_),
    .Q_N(_0577_),
    .Q(stream));
 sg13g2_dfrbp_1 _1132_ (.CLK(clknet_4_5_0_clk_regs),
    .RESET_B(net175),
    .D(_0049_),
    .Q_N(_0576_),
    .Q(\data_out[0] ));
 sg13g2_dfrbp_1 _1133_ (.CLK(clknet_4_4_0_clk_regs),
    .RESET_B(net173),
    .D(_0050_),
    .Q_N(_0575_),
    .Q(\data_out[1] ));
 sg13g2_dfrbp_1 _1134_ (.CLK(clknet_4_6_0_clk_regs),
    .RESET_B(net173),
    .D(_0051_),
    .Q_N(_0574_),
    .Q(\data_out[2] ));
 sg13g2_dfrbp_1 _1135_ (.CLK(clknet_4_2_0_clk_regs),
    .RESET_B(net173),
    .D(_0052_),
    .Q_N(_0573_),
    .Q(\data_out[3] ));
 sg13g2_dfrbp_1 _1136_ (.CLK(clknet_4_2_0_clk_regs),
    .RESET_B(net170),
    .D(_0053_),
    .Q_N(_0572_),
    .Q(\data_out[4] ));
 sg13g2_dfrbp_1 _1137_ (.CLK(clknet_4_4_0_clk_regs),
    .RESET_B(net173),
    .D(_0054_),
    .Q_N(_0571_),
    .Q(\data_out[5] ));
 sg13g2_dfrbp_1 _1138_ (.CLK(clknet_4_4_0_clk_regs),
    .RESET_B(net172),
    .D(_0055_),
    .Q_N(_0570_),
    .Q(\data_out[6] ));
 sg13g2_dfrbp_1 _1139_ (.CLK(clknet_4_4_0_clk_regs),
    .RESET_B(net177),
    .D(_0056_),
    .Q_N(_0569_),
    .Q(\data_out[7] ));
 sg13g2_dfrbp_1 _1140_ (.CLK(clknet_4_7_0_clk_regs),
    .RESET_B(net183),
    .D(_0057_),
    .Q_N(_0568_),
    .Q(\state[0] ));
 sg13g2_dfrbp_1 _1141_ (.CLK(clknet_4_7_0_clk_regs),
    .RESET_B(net183),
    .D(_0058_),
    .Q_N(_0567_),
    .Q(\state[1] ));
 sg13g2_dfrbp_1 _1142_ (.CLK(clknet_4_7_0_clk_regs),
    .RESET_B(net176),
    .D(_0059_),
    .Q_N(_0566_),
    .Q(\state[2] ));
 sg13g2_dfrbp_1 _1143_ (.CLK(clknet_4_7_0_clk_regs),
    .RESET_B(net183),
    .D(_0060_),
    .Q_N(_0565_),
    .Q(\state[3] ));
 sg13g2_dfrbp_1 _1144_ (.CLK(clknet_4_6_0_clk_regs),
    .RESET_B(net176),
    .D(_0061_),
    .Q_N(_0012_),
    .Q(\state[4] ));
 sg13g2_dfrbp_1 _1145_ (.CLK(clknet_4_8_0_clk_regs),
    .RESET_B(net182),
    .D(_0062_),
    .Q_N(_0017_),
    .Q(\counter[0] ));
 sg13g2_dfrbp_1 _1146_ (.CLK(clknet_4_3_0_clk_regs),
    .RESET_B(net178),
    .D(_0063_),
    .Q_N(_0564_),
    .Q(\counter[1] ));
 sg13g2_dfrbp_1 _1147_ (.CLK(clknet_4_2_0_clk_regs),
    .RESET_B(net179),
    .D(_0064_),
    .Q_N(_0014_),
    .Q(\counter[2] ));
 sg13g2_dfrbp_1 _1148_ (.CLK(clknet_4_3_0_clk_regs),
    .RESET_B(net179),
    .D(_0065_),
    .Q_N(_0563_),
    .Q(\counter[3] ));
 sg13g2_dfrbp_1 _1149_ (.CLK(clknet_4_3_0_clk_regs),
    .RESET_B(net179),
    .D(_0066_),
    .Q_N(_0562_),
    .Q(\counter[4] ));
 sg13g2_dfrbp_1 _1150_ (.CLK(clknet_4_10_0_clk_regs),
    .RESET_B(net178),
    .D(net107),
    .Q_N(_0561_),
    .Q(\counter[5] ));
 sg13g2_dfrbp_1 _1151_ (.CLK(clknet_4_11_0_clk_regs),
    .RESET_B(net178),
    .D(_0068_),
    .Q_N(_0560_),
    .Q(\counter[6] ));
 sg13g2_dfrbp_1 _1152_ (.CLK(clknet_4_15_0_clk_regs),
    .RESET_B(net182),
    .D(_0069_),
    .Q_N(_0018_),
    .Q(\counter[7] ));
 sg13g2_dfrbp_1 _1153_ (.CLK(clknet_4_11_0_clk_regs),
    .RESET_B(net179),
    .D(net122),
    .Q_N(_0559_),
    .Q(\counter[8] ));
 sg13g2_dfrbp_1 _1154_ (.CLK(clknet_4_11_0_clk_regs),
    .RESET_B(net178),
    .D(_0071_),
    .Q_N(_0558_),
    .Q(\counter[9] ));
 sg13g2_dfrbp_1 _1155_ (.CLK(clknet_4_11_0_clk_regs),
    .RESET_B(net178),
    .D(_0072_),
    .Q_N(_0557_),
    .Q(\counter[10] ));
 sg13g2_dfrbp_1 _1156_ (.CLK(clknet_4_8_0_clk_regs),
    .RESET_B(net182),
    .D(_0073_),
    .Q_N(_0019_),
    .Q(\counter[11] ));
 sg13g2_dfrbp_1 _1157_ (.CLK(clknet_4_10_0_clk_regs),
    .RESET_B(net178),
    .D(_0074_),
    .Q_N(_0556_),
    .Q(\counter[12] ));
 sg13g2_dfrbp_1 _1158_ (.CLK(clknet_4_10_0_clk_regs),
    .RESET_B(net178),
    .D(_0075_),
    .Q_N(_0555_),
    .Q(\counter[13] ));
 sg13g2_dfrbp_1 _1159_ (.CLK(clknet_4_10_0_clk_regs),
    .RESET_B(net178),
    .D(_0076_),
    .Q_N(_0554_),
    .Q(\counter[14] ));
 sg13g2_dfrbp_1 _1160_ (.CLK(clknet_4_3_0_clk_regs),
    .RESET_B(net179),
    .D(net103),
    .Q_N(_0582_),
    .Q(\counter[15] ));
 sg13g2_dfrbp_1 _1161_ (.CLK(clknet_4_14_0_clk_regs),
    .RESET_B(net181),
    .D(net1),
    .Q_N(_0583_),
    .Q(\inbuf[0] ));
 sg13g2_dfrbp_1 _1162_ (.CLK(clknet_4_13_0_clk_regs),
    .RESET_B(net181),
    .D(net2),
    .Q_N(_0584_),
    .Q(\inbuf[1] ));
 sg13g2_dfrbp_1 _1163_ (.CLK(clknet_4_13_0_clk_regs),
    .RESET_B(net180),
    .D(net3),
    .Q_N(_0585_),
    .Q(\inbuf[2] ));
 sg13g2_dfrbp_1 _1164_ (.CLK(clknet_4_13_0_clk_regs),
    .RESET_B(net180),
    .D(net4),
    .Q_N(_0586_),
    .Q(\inbuf[3] ));
 sg13g2_dfrbp_1 _1165_ (.CLK(clknet_4_14_0_clk_regs),
    .RESET_B(net181),
    .D(net5),
    .Q_N(_0587_),
    .Q(\inbuf[4] ));
 sg13g2_dfrbp_1 _1166_ (.CLK(clknet_4_9_0_clk_regs),
    .RESET_B(net180),
    .D(net6),
    .Q_N(_0588_),
    .Q(\inbuf[5] ));
 sg13g2_dfrbp_1 _1167_ (.CLK(clknet_4_9_0_clk_regs),
    .RESET_B(net180),
    .D(net7),
    .Q_N(_0589_),
    .Q(\inbuf[6] ));
 sg13g2_dfrbp_1 _1168_ (.CLK(clknet_4_9_0_clk_regs),
    .RESET_B(net180),
    .D(net8),
    .Q_N(_0590_),
    .Q(\inbuf[7] ));
 sg13g2_dfrbp_1 _1169_ (.CLK(clknet_4_15_0_clk_regs),
    .RESET_B(net181),
    .D(net43),
    .Q_N(_0591_),
    .Q(\inval[0] ));
 sg13g2_dfrbp_1 _1170_ (.CLK(clknet_4_13_0_clk_regs),
    .RESET_B(net181),
    .D(net42),
    .Q_N(_0592_),
    .Q(\inval[1] ));
 sg13g2_dfrbp_1 _1171_ (.CLK(clknet_4_15_0_clk_regs),
    .RESET_B(net182),
    .D(net44),
    .Q_N(_0593_),
    .Q(\inval[2] ));
 sg13g2_dfrbp_1 _1172_ (.CLK(clknet_4_14_0_clk_regs),
    .RESET_B(net181),
    .D(net40),
    .Q_N(_0594_),
    .Q(\inval[3] ));
 sg13g2_dfrbp_1 _1173_ (.CLK(clknet_4_14_0_clk_regs),
    .RESET_B(net182),
    .D(net41),
    .Q_N(_0595_),
    .Q(\inval[4] ));
 sg13g2_dfrbp_1 _1174_ (.CLK(clknet_4_8_0_clk_regs),
    .RESET_B(net180),
    .D(net38),
    .Q_N(_0596_),
    .Q(\inval[5] ));
 sg13g2_dfrbp_1 _1175_ (.CLK(clknet_4_8_0_clk_regs),
    .RESET_B(net180),
    .D(net37),
    .Q_N(_0597_),
    .Q(\inval[6] ));
 sg13g2_dfrbp_1 _1176_ (.CLK(clknet_4_9_0_clk_regs),
    .RESET_B(net180),
    .D(net39),
    .Q_N(_0553_),
    .Q(\inval[7] ));
 sg13g2_dfrbp_1 _1177_ (.CLK(clknet_4_12_0_clk_regs),
    .RESET_B(net183),
    .D(net71),
    .Q_N(_0552_),
    .Q(\timer[0] ));
 sg13g2_dfrbp_1 _1178_ (.CLK(clknet_4_12_0_clk_regs),
    .RESET_B(net183),
    .D(_0079_),
    .Q_N(_0551_),
    .Q(\timer[1] ));
 sg13g2_dfrbp_1 _1179_ (.CLK(clknet_4_12_0_clk_regs),
    .RESET_B(net183),
    .D(net79),
    .Q_N(_0550_),
    .Q(\timer[2] ));
 sg13g2_dfrbp_1 _1180_ (.CLK(clknet_4_12_0_clk_regs),
    .RESET_B(net183),
    .D(_0081_),
    .Q_N(_0549_),
    .Q(\timer[3] ));
 sg13g2_dfrbp_1 _1181_ (.CLK(net148),
    .RESET_B(net172),
    .D(_0082_),
    .Q_N(\spi.treg[1] ),
    .Q(_0024_));
 sg13g2_dfrbp_1 _1182_ (.CLK(net148),
    .RESET_B(net172),
    .D(_0083_),
    .Q_N(\spi.treg[2] ),
    .Q(_0025_));
 sg13g2_dfrbp_1 _1183_ (.CLK(net148),
    .RESET_B(net170),
    .D(_0084_),
    .Q_N(\spi.treg[3] ),
    .Q(_0026_));
 sg13g2_dfrbp_1 _1184_ (.CLK(net150),
    .RESET_B(net171),
    .D(_0085_),
    .Q_N(\spi.treg[4] ),
    .Q(_0027_));
 sg13g2_dfrbp_1 _1185_ (.CLK(net148),
    .RESET_B(net172),
    .D(_0086_),
    .Q_N(\spi.treg[5] ),
    .Q(_0028_));
 sg13g2_dfrbp_1 _1186_ (.CLK(net148),
    .RESET_B(net172),
    .D(_0087_),
    .Q_N(\spi.treg[6] ),
    .Q(_0029_));
 sg13g2_dfrbp_1 _1187_ (.CLK(net148),
    .RESET_B(net174),
    .D(_0088_),
    .Q_N(\spi.treg[7] ),
    .Q(_0030_));
 sg13g2_dfrbp_1 _1188_ (.CLK(net150),
    .RESET_B(net174),
    .D(_0089_),
    .Q_N(\spi.done ),
    .Q(_0031_));
 sg13g2_dfrbp_1 _1189_ (.CLK(net149),
    .RESET_B(net175),
    .D(_0010_),
    .Q_N(_0548_),
    .Q(sck));
 sg13g2_dfrbp_1 _1190_ (.CLK(net150),
    .RESET_B(net174),
    .D(_0090_),
    .Q_N(_0547_),
    .Q(mosi));
 sg13g2_dfrbp_1 _1191_ (.CLK(net149),
    .RESET_B(net175),
    .D(_0091_),
    .Q_N(csb),
    .Q(_0032_));
 sg13g2_dfrbp_1 _1192_ (.CLK(clknet_4_0_0_clk_regs),
    .RESET_B(net173),
    .D(net48),
    .Q_N(_0011_),
    .Q(\spi.hsck ));
 sg13g2_dfrbp_1 _1193_ (.CLK(clknet_4_5_0_clk_regs),
    .RESET_B(net175),
    .D(net55),
    .Q_N(_0016_),
    .Q(\spi.stream ));
 sg13g2_dfrbp_1 _1194_ (.CLK(net149),
    .RESET_B(net176),
    .D(_0094_),
    .Q_N(_0546_),
    .Q(\spi.nbit[0] ));
 sg13g2_dfrbp_1 _1195_ (.CLK(net149),
    .RESET_B(net176),
    .D(_0095_),
    .Q_N(_0545_),
    .Q(\spi.nbit[1] ));
 sg13g2_dfrbp_1 _1196_ (.CLK(net149),
    .RESET_B(net176),
    .D(_0096_),
    .Q_N(_0013_),
    .Q(\spi.nbit[2] ));
 sg13g2_dfrbp_1 _1197_ (.CLK(net29),
    .RESET_B(net175),
    .D(net100),
    .Q_N(_0544_),
    .Q(\spi.d_latched[0] ));
 sg13g2_dfrbp_1 _1198_ (.CLK(net30),
    .RESET_B(net177),
    .D(_0098_),
    .Q_N(_0543_),
    .Q(\spi.d_latched[1] ));
 sg13g2_dfrbp_1 _1199_ (.CLK(net31),
    .RESET_B(net177),
    .D(_0099_),
    .Q_N(_0542_),
    .Q(\spi.d_latched[2] ));
 sg13g2_dfrbp_1 _1200_ (.CLK(net32),
    .RESET_B(net173),
    .D(_0100_),
    .Q_N(_0541_),
    .Q(\spi.d_latched[3] ));
 sg13g2_dfrbp_1 _1201_ (.CLK(net33),
    .RESET_B(net171),
    .D(_0101_),
    .Q_N(_0540_),
    .Q(\spi.d_latched[4] ));
 sg13g2_dfrbp_1 _1202_ (.CLK(net34),
    .RESET_B(net173),
    .D(_0102_),
    .Q_N(_0539_),
    .Q(\spi.d_latched[5] ));
 sg13g2_dfrbp_1 _1203_ (.CLK(net35),
    .RESET_B(net172),
    .D(net81),
    .Q_N(_0538_),
    .Q(\spi.d_latched[6] ));
 sg13g2_dfrbp_1 _1204_ (.CLK(net36),
    .RESET_B(net177),
    .D(_0104_),
    .Q_N(_0598_),
    .Q(\spi.d_latched[7] ));
 sg13g2_dfrbp_1 _1205_ (.CLK(clknet_4_0_0_clk_regs),
    .RESET_B(net170),
    .D(net63),
    .Q_N(_0599_),
    .Q(\spi.count[0] ));
 sg13g2_dfrbp_1 _1206_ (.CLK(clknet_4_1_0_clk_regs),
    .RESET_B(net170),
    .D(net96),
    .Q_N(_0600_),
    .Q(\spi.count[1] ));
 sg13g2_dfrbp_1 _1207_ (.CLK(clknet_4_0_0_clk_regs),
    .RESET_B(net170),
    .D(_0004_),
    .Q_N(_0601_),
    .Q(\spi.count[2] ));
 sg13g2_dfrbp_1 _1208_ (.CLK(clknet_4_0_0_clk_regs),
    .RESET_B(net170),
    .D(net85),
    .Q_N(_0602_),
    .Q(\spi.count[3] ));
 sg13g2_dfrbp_1 _1209_ (.CLK(clknet_4_2_0_clk_regs),
    .RESET_B(net171),
    .D(net87),
    .Q_N(_0603_),
    .Q(\spi.count[4] ));
 sg13g2_dfrbp_1 _1210_ (.CLK(clknet_4_1_0_clk_regs),
    .RESET_B(net170),
    .D(_0007_),
    .Q_N(_0604_),
    .Q(\spi.count[5] ));
 sg13g2_dfrbp_1 _1211_ (.CLK(clknet_4_1_0_clk_regs),
    .RESET_B(net170),
    .D(net69),
    .Q_N(_0605_),
    .Q(\spi.count[6] ));
 sg13g2_dfrbp_1 _1212_ (.CLK(clknet_4_1_0_clk_regs),
    .RESET_B(net171),
    .D(net60),
    .Q_N(_0537_),
    .Q(\spi.count[7] ));
 sg13g2_tiehi tt_um_rte_eink_driver_23 (.L_HI(net23));
 sg13g2_tiehi tt_um_rte_eink_driver_24 (.L_HI(net24));
 sg13g2_tiehi tt_um_rte_eink_driver_25 (.L_HI(net25));
 sg13g2_tiehi tt_um_rte_eink_driver_26 (.L_HI(net26));
 sg13g2_tiehi tt_um_rte_eink_driver_27 (.L_HI(net27));
 sg13g2_inv_1 _0629__1 (.Y(net28),
    .A(clknet_1_0__leaf_clk));
 sg13g2_tielo tt_um_rte_eink_driver_11 (.L_LO(net11));
 sg13g2_tielo tt_um_rte_eink_driver_12 (.L_LO(net12));
 sg13g2_tielo tt_um_rte_eink_driver_13 (.L_LO(net13));
 sg13g2_tielo tt_um_rte_eink_driver_14 (.L_LO(net14));
 sg13g2_tielo tt_um_rte_eink_driver_15 (.L_LO(net15));
 sg13g2_tielo tt_um_rte_eink_driver_16 (.L_LO(net16));
 sg13g2_tielo tt_um_rte_eink_driver_17 (.L_LO(net17));
 sg13g2_tielo tt_um_rte_eink_driver_18 (.L_LO(net18));
 sg13g2_tielo tt_um_rte_eink_driver_19 (.L_LO(net19));
 sg13g2_tielo tt_um_rte_eink_driver_20 (.L_LO(net20));
 sg13g2_tielo tt_um_rte_eink_driver_21 (.L_LO(net21));
 sg13g2_tiehi tt_um_rte_eink_driver_22 (.L_HI(net22));
 sg13g2_buf_1 _1231_ (.A(csb),
    .X(uio_out[0]));
 sg13g2_buf_2 _1232_ (.A(mosi),
    .X(uio_out[1]));
 sg13g2_buf_1 _1233_ (.A(sck),
    .X(uio_out[3]));
 sg13g2_buf_1 _1234_ (.A(resetb),
    .X(uio_out[5]));
 sg13g2_buf_1 _1235_ (.A(dcb),
    .X(uio_out[7]));
 sg13g2_buf_2 fanout140 (.A(_0301_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_0466_),
    .X(net141));
 sg13g2_buf_4 fanout142 (.X(net142),
    .A(_0129_));
 sg13g2_buf_2 fanout143 (.A(net144),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(net124),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_0152_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(net147),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_0147_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(net150),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(net150),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(\spi.hsck ),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(net152),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(net113),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(\counter[10] ),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(net123),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(\counter[9] ),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(net121),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(\counter[7] ),
    .X(net157));
 sg13g2_buf_4 fanout158 (.X(net158),
    .A(net159));
 sg13g2_buf_2 fanout159 (.A(\counter[3] ),
    .X(net159));
 sg13g2_buf_4 fanout160 (.X(net160),
    .A(net161));
 sg13g2_buf_2 fanout161 (.A(\counter[2] ),
    .X(net161));
 sg13g2_buf_4 fanout162 (.X(net162),
    .A(net163));
 sg13g2_buf_2 fanout163 (.A(\counter[1] ),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(\counter[0] ),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(\counter[0] ),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(net82),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(\state[4] ),
    .X(net167));
 sg13g2_buf_4 fanout168 (.X(net168),
    .A(net120));
 sg13g2_buf_2 fanout169 (.A(net125),
    .X(net169));
 sg13g2_buf_4 fanout170 (.X(net170),
    .A(net172));
 sg13g2_buf_2 fanout171 (.A(net172),
    .X(net171));
 sg13g2_buf_4 fanout172 (.X(net172),
    .A(net173));
 sg13g2_buf_4 fanout173 (.X(net173),
    .A(net177));
 sg13g2_buf_4 fanout174 (.X(net174),
    .A(net175));
 sg13g2_buf_4 fanout175 (.X(net175),
    .A(net176));
 sg13g2_buf_4 fanout176 (.X(net176),
    .A(net177));
 sg13g2_buf_4 fanout177 (.X(net177),
    .A(rst_n));
 sg13g2_buf_4 fanout178 (.X(net178),
    .A(net179));
 sg13g2_buf_4 fanout179 (.X(net179),
    .A(rst_n));
 sg13g2_buf_4 fanout180 (.X(net180),
    .A(net182));
 sg13g2_buf_4 fanout181 (.X(net181),
    .A(net182));
 sg13g2_buf_4 fanout182 (.X(net182),
    .A(net183));
 sg13g2_buf_4 fanout183 (.X(net183),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[6]),
    .X(net9));
 sg13g2_tielo tt_um_rte_eink_driver_10 (.L_LO(net10));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(delaynet_0_clk));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_1_1__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_0_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_0_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_1_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_1_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_2_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_2_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_3_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_3_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_4_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_4_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_5_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_5_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_6_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_6_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_7_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_7_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_8_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_8_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_9_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_9_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_10_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_10_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_11_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_11_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_12_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_12_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_13_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_13_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_14_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_14_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_15_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_15_0_clk_regs));
 sg13g2_inv_1 clkload1 (.A(clknet_4_15_0_clk_regs));
 sg13g2_buf_2 delaybuf_0_clk (.A(delaynet_0_clk),
    .X(clknet_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\inbuf[6] ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold2 (.A(\inbuf[5] ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold3 (.A(\inbuf[7] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold4 (.A(\inbuf[3] ),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold5 (.A(\inbuf[4] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold6 (.A(\inbuf[1] ),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold7 (.A(\inbuf[0] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold8 (.A(\inbuf[2] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0017_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0470_),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0011_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0092_),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold13 (.A(\data_out[6] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold14 (.A(\data_out[7] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold15 (.A(\data_out[3] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold16 (.A(\data_out[5] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold17 (.A(\data_out[2] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold18 (.A(stream),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0093_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold20 (.A(\data_out[0] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0023_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0242_),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold23 (.A(\spi.count[7] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0009_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0022_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold26 (.A(\spi.count[0] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0002_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold28 (.A(\spi.d_latched[1] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold29 (.A(\spi.d_latched[4] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold30 (.A(\data_out[4] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold31 (.A(\data_out[1] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold32 (.A(\spi.count[6] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0008_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold34 (.A(\timer[0] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0078_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold36 (.A(\counter[10] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0492_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold38 (.A(\spi.d_latched[7] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold39 (.A(\timer[3] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0510_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold41 (.A(\timer[2] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0508_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0080_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold44 (.A(\spi.d_latched[6] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0103_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0012_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0244_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold48 (.A(\spi.count[3] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0005_),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold50 (.A(\spi.count[4] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0006_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold52 (.A(\spi.d_latched[5] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold53 (.A(\state[4] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold54 (.A(\timer[1] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold55 (.A(\spi.d_latched[3] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0018_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0487_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold58 (.A(\spi.d_latched[2] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold59 (.A(\spi.count[1] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0003_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold61 (.A(\counter[12] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0497_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold63 (.A(\spi.d_latched[0] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0097_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold65 (.A(\counter[15] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0503_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0077_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold68 (.A(\counter[13] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold69 (.A(\counter[4] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold70 (.A(\counter[5] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0067_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold72 (.A(\spi.reg_dat_we ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0014_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0478_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold75 (.A(\spi.count[2] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold76 (.A(\spi.count[5] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold77 (.A(\counter[11] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0495_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold79 (.A(\state[3] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold80 (.A(\counter[14] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold81 (.A(\counter[6] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0485_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold83 (.A(\state[2] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold84 (.A(\state[1] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold85 (.A(\counter[8] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0070_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold87 (.A(\counter[9] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold88 (.A(\spi.w_latched ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold89 (.A(\state[0] ),
    .X(net125));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_fill_2 FILLER_12_70 ();
 sg13g2_fill_1 FILLER_12_72 ();
 sg13g2_fill_2 FILLER_12_79 ();
 sg13g2_fill_1 FILLER_12_81 ();
 sg13g2_decap_4 FILLER_12_87 ();
 sg13g2_fill_1 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_101 ();
 sg13g2_decap_8 FILLER_12_108 ();
 sg13g2_decap_8 FILLER_12_115 ();
 sg13g2_decap_8 FILLER_12_122 ();
 sg13g2_decap_8 FILLER_12_129 ();
 sg13g2_decap_8 FILLER_12_136 ();
 sg13g2_decap_8 FILLER_12_143 ();
 sg13g2_decap_8 FILLER_12_150 ();
 sg13g2_decap_8 FILLER_12_157 ();
 sg13g2_decap_8 FILLER_12_164 ();
 sg13g2_decap_8 FILLER_12_171 ();
 sg13g2_decap_8 FILLER_12_178 ();
 sg13g2_decap_8 FILLER_12_185 ();
 sg13g2_decap_8 FILLER_12_192 ();
 sg13g2_decap_8 FILLER_12_199 ();
 sg13g2_decap_8 FILLER_12_206 ();
 sg13g2_decap_8 FILLER_12_213 ();
 sg13g2_decap_8 FILLER_12_220 ();
 sg13g2_decap_8 FILLER_12_227 ();
 sg13g2_decap_8 FILLER_12_234 ();
 sg13g2_decap_8 FILLER_12_241 ();
 sg13g2_decap_8 FILLER_12_248 ();
 sg13g2_decap_8 FILLER_12_255 ();
 sg13g2_decap_8 FILLER_12_262 ();
 sg13g2_decap_8 FILLER_12_269 ();
 sg13g2_decap_8 FILLER_12_276 ();
 sg13g2_decap_8 FILLER_12_283 ();
 sg13g2_decap_8 FILLER_12_290 ();
 sg13g2_decap_8 FILLER_12_297 ();
 sg13g2_decap_8 FILLER_12_304 ();
 sg13g2_decap_8 FILLER_12_311 ();
 sg13g2_decap_8 FILLER_12_318 ();
 sg13g2_decap_8 FILLER_12_325 ();
 sg13g2_decap_8 FILLER_12_332 ();
 sg13g2_decap_8 FILLER_12_339 ();
 sg13g2_decap_8 FILLER_12_346 ();
 sg13g2_decap_8 FILLER_12_353 ();
 sg13g2_decap_8 FILLER_12_360 ();
 sg13g2_decap_8 FILLER_12_367 ();
 sg13g2_decap_8 FILLER_12_374 ();
 sg13g2_decap_8 FILLER_12_381 ();
 sg13g2_decap_8 FILLER_12_388 ();
 sg13g2_decap_8 FILLER_12_395 ();
 sg13g2_decap_8 FILLER_12_402 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_fill_2 FILLER_13_14 ();
 sg13g2_fill_1 FILLER_13_54 ();
 sg13g2_decap_8 FILLER_13_127 ();
 sg13g2_decap_8 FILLER_13_134 ();
 sg13g2_decap_8 FILLER_13_141 ();
 sg13g2_decap_8 FILLER_13_148 ();
 sg13g2_decap_8 FILLER_13_155 ();
 sg13g2_decap_8 FILLER_13_162 ();
 sg13g2_decap_8 FILLER_13_169 ();
 sg13g2_decap_8 FILLER_13_176 ();
 sg13g2_decap_8 FILLER_13_183 ();
 sg13g2_decap_8 FILLER_13_190 ();
 sg13g2_decap_8 FILLER_13_197 ();
 sg13g2_decap_8 FILLER_13_204 ();
 sg13g2_decap_8 FILLER_13_211 ();
 sg13g2_decap_8 FILLER_13_218 ();
 sg13g2_decap_8 FILLER_13_225 ();
 sg13g2_decap_8 FILLER_13_232 ();
 sg13g2_decap_8 FILLER_13_239 ();
 sg13g2_decap_8 FILLER_13_246 ();
 sg13g2_decap_8 FILLER_13_253 ();
 sg13g2_decap_8 FILLER_13_260 ();
 sg13g2_decap_8 FILLER_13_267 ();
 sg13g2_decap_8 FILLER_13_274 ();
 sg13g2_decap_8 FILLER_13_281 ();
 sg13g2_decap_8 FILLER_13_288 ();
 sg13g2_decap_8 FILLER_13_295 ();
 sg13g2_decap_8 FILLER_13_302 ();
 sg13g2_decap_8 FILLER_13_309 ();
 sg13g2_decap_8 FILLER_13_316 ();
 sg13g2_decap_8 FILLER_13_323 ();
 sg13g2_decap_8 FILLER_13_330 ();
 sg13g2_decap_8 FILLER_13_337 ();
 sg13g2_decap_8 FILLER_13_344 ();
 sg13g2_decap_8 FILLER_13_351 ();
 sg13g2_decap_8 FILLER_13_358 ();
 sg13g2_decap_8 FILLER_13_365 ();
 sg13g2_decap_8 FILLER_13_372 ();
 sg13g2_decap_8 FILLER_13_379 ();
 sg13g2_decap_8 FILLER_13_386 ();
 sg13g2_decap_8 FILLER_13_393 ();
 sg13g2_decap_8 FILLER_13_400 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_4 FILLER_14_21 ();
 sg13g2_fill_2 FILLER_14_25 ();
 sg13g2_fill_1 FILLER_14_70 ();
 sg13g2_decap_4 FILLER_14_92 ();
 sg13g2_decap_8 FILLER_14_131 ();
 sg13g2_decap_8 FILLER_14_138 ();
 sg13g2_decap_8 FILLER_14_145 ();
 sg13g2_decap_8 FILLER_14_152 ();
 sg13g2_decap_8 FILLER_14_159 ();
 sg13g2_decap_8 FILLER_14_166 ();
 sg13g2_decap_8 FILLER_14_173 ();
 sg13g2_decap_8 FILLER_14_180 ();
 sg13g2_decap_8 FILLER_14_187 ();
 sg13g2_decap_8 FILLER_14_194 ();
 sg13g2_decap_8 FILLER_14_201 ();
 sg13g2_decap_8 FILLER_14_208 ();
 sg13g2_decap_8 FILLER_14_215 ();
 sg13g2_decap_8 FILLER_14_222 ();
 sg13g2_decap_8 FILLER_14_229 ();
 sg13g2_decap_8 FILLER_14_236 ();
 sg13g2_decap_8 FILLER_14_243 ();
 sg13g2_decap_8 FILLER_14_250 ();
 sg13g2_decap_8 FILLER_14_257 ();
 sg13g2_decap_8 FILLER_14_264 ();
 sg13g2_decap_8 FILLER_14_271 ();
 sg13g2_decap_8 FILLER_14_278 ();
 sg13g2_decap_8 FILLER_14_285 ();
 sg13g2_decap_8 FILLER_14_292 ();
 sg13g2_decap_8 FILLER_14_299 ();
 sg13g2_decap_8 FILLER_14_306 ();
 sg13g2_decap_8 FILLER_14_313 ();
 sg13g2_decap_8 FILLER_14_320 ();
 sg13g2_decap_8 FILLER_14_327 ();
 sg13g2_decap_8 FILLER_14_334 ();
 sg13g2_decap_8 FILLER_14_341 ();
 sg13g2_decap_8 FILLER_14_348 ();
 sg13g2_decap_8 FILLER_14_355 ();
 sg13g2_decap_8 FILLER_14_362 ();
 sg13g2_decap_8 FILLER_14_369 ();
 sg13g2_decap_8 FILLER_14_376 ();
 sg13g2_decap_8 FILLER_14_383 ();
 sg13g2_decap_8 FILLER_14_390 ();
 sg13g2_decap_8 FILLER_14_397 ();
 sg13g2_decap_4 FILLER_14_404 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_37 ();
 sg13g2_fill_1 FILLER_15_39 ();
 sg13g2_decap_4 FILLER_15_49 ();
 sg13g2_fill_2 FILLER_15_76 ();
 sg13g2_decap_8 FILLER_15_121 ();
 sg13g2_decap_8 FILLER_15_128 ();
 sg13g2_decap_8 FILLER_15_135 ();
 sg13g2_decap_8 FILLER_15_142 ();
 sg13g2_decap_8 FILLER_15_149 ();
 sg13g2_decap_8 FILLER_15_156 ();
 sg13g2_decap_8 FILLER_15_163 ();
 sg13g2_decap_8 FILLER_15_170 ();
 sg13g2_decap_8 FILLER_15_177 ();
 sg13g2_decap_8 FILLER_15_184 ();
 sg13g2_decap_8 FILLER_15_191 ();
 sg13g2_decap_8 FILLER_15_198 ();
 sg13g2_decap_8 FILLER_15_205 ();
 sg13g2_decap_8 FILLER_15_212 ();
 sg13g2_decap_8 FILLER_15_219 ();
 sg13g2_decap_8 FILLER_15_226 ();
 sg13g2_decap_8 FILLER_15_233 ();
 sg13g2_decap_8 FILLER_15_240 ();
 sg13g2_decap_8 FILLER_15_247 ();
 sg13g2_decap_8 FILLER_15_254 ();
 sg13g2_decap_8 FILLER_15_261 ();
 sg13g2_decap_8 FILLER_15_268 ();
 sg13g2_decap_8 FILLER_15_275 ();
 sg13g2_decap_8 FILLER_15_282 ();
 sg13g2_decap_8 FILLER_15_289 ();
 sg13g2_decap_8 FILLER_15_296 ();
 sg13g2_decap_8 FILLER_15_303 ();
 sg13g2_decap_8 FILLER_15_310 ();
 sg13g2_decap_8 FILLER_15_317 ();
 sg13g2_decap_8 FILLER_15_324 ();
 sg13g2_decap_8 FILLER_15_331 ();
 sg13g2_decap_8 FILLER_15_338 ();
 sg13g2_decap_8 FILLER_15_345 ();
 sg13g2_decap_8 FILLER_15_352 ();
 sg13g2_decap_8 FILLER_15_359 ();
 sg13g2_decap_8 FILLER_15_366 ();
 sg13g2_decap_8 FILLER_15_373 ();
 sg13g2_decap_8 FILLER_15_380 ();
 sg13g2_decap_8 FILLER_15_387 ();
 sg13g2_decap_8 FILLER_15_394 ();
 sg13g2_decap_8 FILLER_15_401 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_4 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_20 ();
 sg13g2_fill_1 FILLER_16_27 ();
 sg13g2_fill_1 FILLER_16_102 ();
 sg13g2_decap_8 FILLER_16_129 ();
 sg13g2_decap_8 FILLER_16_136 ();
 sg13g2_decap_8 FILLER_16_143 ();
 sg13g2_decap_8 FILLER_16_150 ();
 sg13g2_decap_8 FILLER_16_157 ();
 sg13g2_decap_8 FILLER_16_164 ();
 sg13g2_decap_8 FILLER_16_171 ();
 sg13g2_decap_8 FILLER_16_178 ();
 sg13g2_decap_8 FILLER_16_185 ();
 sg13g2_decap_8 FILLER_16_192 ();
 sg13g2_decap_8 FILLER_16_199 ();
 sg13g2_decap_8 FILLER_16_206 ();
 sg13g2_decap_8 FILLER_16_213 ();
 sg13g2_decap_8 FILLER_16_220 ();
 sg13g2_decap_8 FILLER_16_227 ();
 sg13g2_decap_8 FILLER_16_234 ();
 sg13g2_decap_8 FILLER_16_241 ();
 sg13g2_decap_8 FILLER_16_248 ();
 sg13g2_decap_8 FILLER_16_255 ();
 sg13g2_decap_8 FILLER_16_262 ();
 sg13g2_decap_8 FILLER_16_269 ();
 sg13g2_decap_8 FILLER_16_276 ();
 sg13g2_decap_8 FILLER_16_283 ();
 sg13g2_decap_8 FILLER_16_290 ();
 sg13g2_decap_8 FILLER_16_297 ();
 sg13g2_decap_8 FILLER_16_304 ();
 sg13g2_decap_8 FILLER_16_311 ();
 sg13g2_decap_8 FILLER_16_318 ();
 sg13g2_decap_8 FILLER_16_325 ();
 sg13g2_decap_4 FILLER_16_332 ();
 sg13g2_fill_2 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_342 ();
 sg13g2_decap_8 FILLER_16_349 ();
 sg13g2_decap_8 FILLER_16_356 ();
 sg13g2_decap_8 FILLER_16_363 ();
 sg13g2_decap_8 FILLER_16_370 ();
 sg13g2_decap_8 FILLER_16_377 ();
 sg13g2_decap_8 FILLER_16_384 ();
 sg13g2_decap_8 FILLER_16_391 ();
 sg13g2_decap_8 FILLER_16_398 ();
 sg13g2_decap_4 FILLER_16_405 ();
 sg13g2_decap_4 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_4 ();
 sg13g2_decap_4 FILLER_17_47 ();
 sg13g2_decap_8 FILLER_17_59 ();
 sg13g2_decap_8 FILLER_17_66 ();
 sg13g2_decap_8 FILLER_17_73 ();
 sg13g2_decap_8 FILLER_17_80 ();
 sg13g2_fill_2 FILLER_17_87 ();
 sg13g2_fill_1 FILLER_17_89 ();
 sg13g2_decap_4 FILLER_17_95 ();
 sg13g2_fill_1 FILLER_17_99 ();
 sg13g2_fill_2 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_123 ();
 sg13g2_decap_4 FILLER_17_130 ();
 sg13g2_fill_2 FILLER_17_134 ();
 sg13g2_decap_8 FILLER_17_145 ();
 sg13g2_decap_4 FILLER_17_152 ();
 sg13g2_fill_1 FILLER_17_156 ();
 sg13g2_decap_8 FILLER_17_160 ();
 sg13g2_fill_2 FILLER_17_167 ();
 sg13g2_decap_8 FILLER_17_172 ();
 sg13g2_decap_8 FILLER_17_179 ();
 sg13g2_decap_8 FILLER_17_186 ();
 sg13g2_decap_8 FILLER_17_193 ();
 sg13g2_decap_8 FILLER_17_200 ();
 sg13g2_decap_8 FILLER_17_207 ();
 sg13g2_decap_8 FILLER_17_214 ();
 sg13g2_decap_8 FILLER_17_221 ();
 sg13g2_decap_8 FILLER_17_228 ();
 sg13g2_decap_4 FILLER_17_235 ();
 sg13g2_fill_1 FILLER_17_239 ();
 sg13g2_decap_8 FILLER_17_244 ();
 sg13g2_decap_8 FILLER_17_251 ();
 sg13g2_decap_4 FILLER_17_258 ();
 sg13g2_decap_8 FILLER_17_276 ();
 sg13g2_decap_8 FILLER_17_283 ();
 sg13g2_fill_2 FILLER_17_290 ();
 sg13g2_fill_1 FILLER_17_292 ();
 sg13g2_fill_2 FILLER_17_324 ();
 sg13g2_fill_1 FILLER_17_326 ();
 sg13g2_fill_1 FILLER_17_353 ();
 sg13g2_decap_8 FILLER_17_362 ();
 sg13g2_decap_8 FILLER_17_369 ();
 sg13g2_decap_8 FILLER_17_376 ();
 sg13g2_decap_8 FILLER_17_383 ();
 sg13g2_decap_8 FILLER_17_390 ();
 sg13g2_decap_8 FILLER_17_397 ();
 sg13g2_decap_4 FILLER_17_404 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_37 ();
 sg13g2_fill_2 FILLER_18_129 ();
 sg13g2_fill_1 FILLER_18_131 ();
 sg13g2_fill_2 FILLER_18_162 ();
 sg13g2_decap_8 FILLER_18_190 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_4 FILLER_18_231 ();
 sg13g2_decap_4 FILLER_18_310 ();
 sg13g2_decap_4 FILLER_18_319 ();
 sg13g2_fill_2 FILLER_18_342 ();
 sg13g2_fill_2 FILLER_18_353 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_4 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_4 ();
 sg13g2_decap_8 FILLER_19_52 ();
 sg13g2_decap_4 FILLER_19_59 ();
 sg13g2_fill_1 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_76 ();
 sg13g2_fill_2 FILLER_19_83 ();
 sg13g2_fill_2 FILLER_19_116 ();
 sg13g2_fill_1 FILLER_19_118 ();
 sg13g2_fill_2 FILLER_19_157 ();
 sg13g2_fill_1 FILLER_19_169 ();
 sg13g2_fill_1 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_216 ();
 sg13g2_decap_8 FILLER_19_223 ();
 sg13g2_decap_4 FILLER_19_230 ();
 sg13g2_fill_1 FILLER_19_234 ();
 sg13g2_fill_2 FILLER_19_260 ();
 sg13g2_fill_2 FILLER_19_270 ();
 sg13g2_fill_1 FILLER_19_272 ();
 sg13g2_decap_8 FILLER_19_278 ();
 sg13g2_decap_8 FILLER_19_285 ();
 sg13g2_fill_1 FILLER_19_303 ();
 sg13g2_fill_1 FILLER_19_316 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_fill_1 FILLER_20_70 ();
 sg13g2_fill_1 FILLER_20_75 ();
 sg13g2_decap_4 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_97 ();
 sg13g2_fill_1 FILLER_20_104 ();
 sg13g2_decap_8 FILLER_20_120 ();
 sg13g2_fill_2 FILLER_20_127 ();
 sg13g2_fill_1 FILLER_20_173 ();
 sg13g2_fill_2 FILLER_20_239 ();
 sg13g2_fill_2 FILLER_20_268 ();
 sg13g2_decap_4 FILLER_20_316 ();
 sg13g2_fill_2 FILLER_20_320 ();
 sg13g2_decap_4 FILLER_20_330 ();
 sg13g2_fill_2 FILLER_20_334 ();
 sg13g2_decap_4 FILLER_20_346 ();
 sg13g2_decap_8 FILLER_20_376 ();
 sg13g2_fill_1 FILLER_20_383 ();
 sg13g2_decap_4 FILLER_20_389 ();
 sg13g2_fill_2 FILLER_20_393 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_7 ();
 sg13g2_fill_2 FILLER_21_43 ();
 sg13g2_fill_1 FILLER_21_45 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_fill_2 FILLER_21_84 ();
 sg13g2_fill_2 FILLER_21_116 ();
 sg13g2_decap_8 FILLER_21_183 ();
 sg13g2_fill_2 FILLER_21_202 ();
 sg13g2_decap_4 FILLER_21_209 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_fill_1 FILLER_21_231 ();
 sg13g2_fill_1 FILLER_21_256 ();
 sg13g2_fill_2 FILLER_21_269 ();
 sg13g2_decap_4 FILLER_21_276 ();
 sg13g2_fill_2 FILLER_21_299 ();
 sg13g2_fill_1 FILLER_21_301 ();
 sg13g2_fill_1 FILLER_21_328 ();
 sg13g2_fill_1 FILLER_21_339 ();
 sg13g2_fill_1 FILLER_21_345 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_4 FILLER_21_371 ();
 sg13g2_fill_2 FILLER_21_375 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_fill_2 FILLER_22_40 ();
 sg13g2_fill_2 FILLER_22_68 ();
 sg13g2_fill_1 FILLER_22_70 ();
 sg13g2_fill_1 FILLER_22_100 ();
 sg13g2_fill_2 FILLER_22_110 ();
 sg13g2_fill_1 FILLER_22_112 ();
 sg13g2_decap_4 FILLER_22_118 ();
 sg13g2_fill_1 FILLER_22_122 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_fill_1 FILLER_22_140 ();
 sg13g2_fill_1 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_160 ();
 sg13g2_fill_2 FILLER_22_171 ();
 sg13g2_fill_1 FILLER_22_184 ();
 sg13g2_decap_8 FILLER_22_190 ();
 sg13g2_decap_8 FILLER_22_197 ();
 sg13g2_decap_8 FILLER_22_227 ();
 sg13g2_decap_8 FILLER_22_234 ();
 sg13g2_decap_8 FILLER_22_241 ();
 sg13g2_fill_2 FILLER_22_248 ();
 sg13g2_fill_1 FILLER_22_250 ();
 sg13g2_fill_1 FILLER_22_275 ();
 sg13g2_fill_2 FILLER_22_283 ();
 sg13g2_fill_1 FILLER_22_285 ();
 sg13g2_fill_2 FILLER_22_309 ();
 sg13g2_fill_1 FILLER_22_311 ();
 sg13g2_fill_2 FILLER_22_321 ();
 sg13g2_decap_8 FILLER_22_328 ();
 sg13g2_fill_2 FILLER_22_379 ();
 sg13g2_fill_1 FILLER_22_381 ();
 sg13g2_decap_4 FILLER_22_396 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_4 ();
 sg13g2_decap_8 FILLER_23_41 ();
 sg13g2_decap_8 FILLER_23_48 ();
 sg13g2_fill_2 FILLER_23_55 ();
 sg13g2_fill_1 FILLER_23_57 ();
 sg13g2_fill_2 FILLER_23_78 ();
 sg13g2_fill_1 FILLER_23_80 ();
 sg13g2_decap_8 FILLER_23_121 ();
 sg13g2_decap_4 FILLER_23_146 ();
 sg13g2_fill_1 FILLER_23_150 ();
 sg13g2_fill_2 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_178 ();
 sg13g2_decap_4 FILLER_23_195 ();
 sg13g2_fill_2 FILLER_23_199 ();
 sg13g2_fill_2 FILLER_23_208 ();
 sg13g2_decap_4 FILLER_23_233 ();
 sg13g2_fill_2 FILLER_23_237 ();
 sg13g2_decap_8 FILLER_23_244 ();
 sg13g2_decap_8 FILLER_23_251 ();
 sg13g2_decap_4 FILLER_23_258 ();
 sg13g2_fill_1 FILLER_23_262 ();
 sg13g2_decap_4 FILLER_23_271 ();
 sg13g2_fill_1 FILLER_23_275 ();
 sg13g2_fill_1 FILLER_23_299 ();
 sg13g2_decap_8 FILLER_23_331 ();
 sg13g2_fill_1 FILLER_23_338 ();
 sg13g2_fill_2 FILLER_23_363 ();
 sg13g2_decap_4 FILLER_23_370 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_4 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_62 ();
 sg13g2_decap_8 FILLER_24_69 ();
 sg13g2_decap_8 FILLER_24_76 ();
 sg13g2_decap_4 FILLER_24_83 ();
 sg13g2_fill_2 FILLER_24_87 ();
 sg13g2_fill_2 FILLER_24_112 ();
 sg13g2_fill_1 FILLER_24_114 ();
 sg13g2_decap_8 FILLER_24_146 ();
 sg13g2_fill_2 FILLER_24_153 ();
 sg13g2_fill_1 FILLER_24_155 ();
 sg13g2_decap_4 FILLER_24_160 ();
 sg13g2_fill_2 FILLER_24_164 ();
 sg13g2_decap_8 FILLER_24_174 ();
 sg13g2_decap_4 FILLER_24_194 ();
 sg13g2_fill_1 FILLER_24_198 ();
 sg13g2_fill_2 FILLER_24_215 ();
 sg13g2_decap_4 FILLER_24_233 ();
 sg13g2_fill_1 FILLER_24_237 ();
 sg13g2_decap_4 FILLER_24_250 ();
 sg13g2_fill_2 FILLER_24_272 ();
 sg13g2_fill_1 FILLER_24_274 ();
 sg13g2_decap_8 FILLER_24_281 ();
 sg13g2_decap_8 FILLER_24_298 ();
 sg13g2_decap_8 FILLER_24_305 ();
 sg13g2_decap_8 FILLER_24_312 ();
 sg13g2_fill_1 FILLER_24_319 ();
 sg13g2_decap_8 FILLER_24_325 ();
 sg13g2_fill_2 FILLER_24_353 ();
 sg13g2_fill_1 FILLER_24_355 ();
 sg13g2_decap_8 FILLER_24_385 ();
 sg13g2_fill_1 FILLER_24_392 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_50 ();
 sg13g2_decap_8 FILLER_25_57 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_4 FILLER_25_84 ();
 sg13g2_fill_1 FILLER_25_97 ();
 sg13g2_fill_2 FILLER_25_121 ();
 sg13g2_fill_1 FILLER_25_123 ();
 sg13g2_fill_1 FILLER_25_134 ();
 sg13g2_decap_4 FILLER_25_149 ();
 sg13g2_fill_1 FILLER_25_153 ();
 sg13g2_fill_1 FILLER_25_179 ();
 sg13g2_fill_2 FILLER_25_196 ();
 sg13g2_fill_1 FILLER_25_198 ();
 sg13g2_decap_8 FILLER_25_215 ();
 sg13g2_decap_8 FILLER_25_228 ();
 sg13g2_fill_2 FILLER_25_235 ();
 sg13g2_fill_2 FILLER_25_260 ();
 sg13g2_decap_8 FILLER_25_267 ();
 sg13g2_fill_2 FILLER_25_274 ();
 sg13g2_decap_8 FILLER_25_281 ();
 sg13g2_fill_1 FILLER_25_288 ();
 sg13g2_fill_2 FILLER_25_306 ();
 sg13g2_fill_1 FILLER_25_308 ();
 sg13g2_decap_4 FILLER_25_323 ();
 sg13g2_fill_2 FILLER_25_327 ();
 sg13g2_fill_1 FILLER_25_334 ();
 sg13g2_decap_8 FILLER_25_357 ();
 sg13g2_decap_4 FILLER_25_364 ();
 sg13g2_fill_1 FILLER_25_368 ();
 sg13g2_decap_8 FILLER_25_374 ();
 sg13g2_fill_2 FILLER_25_381 ();
 sg13g2_decap_4 FILLER_25_388 ();
 sg13g2_decap_8 FILLER_25_402 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_fill_1 FILLER_26_14 ();
 sg13g2_fill_1 FILLER_26_41 ();
 sg13g2_fill_1 FILLER_26_52 ();
 sg13g2_fill_2 FILLER_26_124 ();
 sg13g2_decap_8 FILLER_26_156 ();
 sg13g2_fill_1 FILLER_26_163 ();
 sg13g2_decap_4 FILLER_26_180 ();
 sg13g2_fill_1 FILLER_26_184 ();
 sg13g2_fill_1 FILLER_26_190 ();
 sg13g2_decap_4 FILLER_26_201 ();
 sg13g2_fill_2 FILLER_26_205 ();
 sg13g2_decap_4 FILLER_26_229 ();
 sg13g2_decap_8 FILLER_26_249 ();
 sg13g2_decap_4 FILLER_26_256 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_fill_1 FILLER_26_273 ();
 sg13g2_decap_8 FILLER_26_291 ();
 sg13g2_fill_2 FILLER_26_298 ();
 sg13g2_fill_1 FILLER_26_300 ();
 sg13g2_fill_1 FILLER_26_306 ();
 sg13g2_fill_2 FILLER_26_322 ();
 sg13g2_fill_1 FILLER_26_324 ();
 sg13g2_fill_1 FILLER_26_331 ();
 sg13g2_fill_2 FILLER_26_357 ();
 sg13g2_fill_1 FILLER_26_379 ();
 sg13g2_decap_4 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_fill_2 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_47 ();
 sg13g2_decap_8 FILLER_27_62 ();
 sg13g2_decap_4 FILLER_27_69 ();
 sg13g2_fill_1 FILLER_27_73 ();
 sg13g2_decap_4 FILLER_27_77 ();
 sg13g2_fill_1 FILLER_27_81 ();
 sg13g2_fill_1 FILLER_27_91 ();
 sg13g2_fill_1 FILLER_27_104 ();
 sg13g2_fill_2 FILLER_27_129 ();
 sg13g2_decap_8 FILLER_27_134 ();
 sg13g2_fill_2 FILLER_27_141 ();
 sg13g2_fill_1 FILLER_27_143 ();
 sg13g2_decap_8 FILLER_27_148 ();
 sg13g2_decap_8 FILLER_27_155 ();
 sg13g2_fill_2 FILLER_27_162 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_decap_4 FILLER_27_182 ();
 sg13g2_fill_1 FILLER_27_186 ();
 sg13g2_fill_2 FILLER_27_191 ();
 sg13g2_fill_1 FILLER_27_201 ();
 sg13g2_fill_2 FILLER_27_213 ();
 sg13g2_fill_1 FILLER_27_215 ();
 sg13g2_decap_8 FILLER_27_221 ();
 sg13g2_fill_2 FILLER_27_228 ();
 sg13g2_fill_1 FILLER_27_230 ();
 sg13g2_fill_1 FILLER_27_238 ();
 sg13g2_fill_2 FILLER_27_249 ();
 sg13g2_fill_1 FILLER_27_251 ();
 sg13g2_decap_4 FILLER_27_257 ();
 sg13g2_fill_2 FILLER_27_261 ();
 sg13g2_decap_8 FILLER_27_274 ();
 sg13g2_decap_8 FILLER_27_303 ();
 sg13g2_fill_2 FILLER_27_310 ();
 sg13g2_decap_8 FILLER_27_320 ();
 sg13g2_decap_8 FILLER_27_327 ();
 sg13g2_fill_2 FILLER_27_334 ();
 sg13g2_fill_1 FILLER_27_336 ();
 sg13g2_decap_4 FILLER_27_352 ();
 sg13g2_fill_1 FILLER_27_356 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_fill_1 FILLER_27_385 ();
 sg13g2_fill_1 FILLER_27_391 ();
 sg13g2_decap_8 FILLER_27_397 ();
 sg13g2_decap_4 FILLER_27_404 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_4 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_16 ();
 sg13g2_fill_1 FILLER_28_23 ();
 sg13g2_decap_4 FILLER_28_80 ();
 sg13g2_fill_2 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_178 ();
 sg13g2_fill_2 FILLER_28_185 ();
 sg13g2_fill_1 FILLER_28_187 ();
 sg13g2_decap_8 FILLER_28_197 ();
 sg13g2_decap_8 FILLER_28_204 ();
 sg13g2_decap_8 FILLER_28_215 ();
 sg13g2_decap_4 FILLER_28_222 ();
 sg13g2_fill_2 FILLER_28_226 ();
 sg13g2_decap_8 FILLER_28_233 ();
 sg13g2_decap_4 FILLER_28_240 ();
 sg13g2_decap_4 FILLER_28_255 ();
 sg13g2_fill_1 FILLER_28_259 ();
 sg13g2_decap_8 FILLER_28_280 ();
 sg13g2_decap_4 FILLER_28_287 ();
 sg13g2_fill_2 FILLER_28_304 ();
 sg13g2_fill_1 FILLER_28_306 ();
 sg13g2_decap_4 FILLER_28_315 ();
 sg13g2_fill_1 FILLER_28_319 ();
 sg13g2_decap_8 FILLER_28_345 ();
 sg13g2_decap_4 FILLER_28_352 ();
 sg13g2_decap_8 FILLER_28_370 ();
 sg13g2_decap_4 FILLER_28_377 ();
 sg13g2_fill_2 FILLER_28_381 ();
 sg13g2_fill_2 FILLER_28_389 ();
 sg13g2_decap_4 FILLER_28_403 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_4 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_45 ();
 sg13g2_fill_2 FILLER_29_52 ();
 sg13g2_decap_4 FILLER_29_59 ();
 sg13g2_fill_1 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_93 ();
 sg13g2_decap_4 FILLER_29_100 ();
 sg13g2_fill_2 FILLER_29_114 ();
 sg13g2_fill_1 FILLER_29_116 ();
 sg13g2_decap_4 FILLER_29_122 ();
 sg13g2_fill_2 FILLER_29_136 ();
 sg13g2_fill_1 FILLER_29_138 ();
 sg13g2_decap_8 FILLER_29_148 ();
 sg13g2_decap_8 FILLER_29_155 ();
 sg13g2_fill_1 FILLER_29_162 ();
 sg13g2_fill_2 FILLER_29_172 ();
 sg13g2_fill_1 FILLER_29_174 ();
 sg13g2_decap_8 FILLER_29_180 ();
 sg13g2_fill_1 FILLER_29_187 ();
 sg13g2_decap_4 FILLER_29_201 ();
 sg13g2_decap_4 FILLER_29_222 ();
 sg13g2_decap_8 FILLER_29_245 ();
 sg13g2_decap_8 FILLER_29_252 ();
 sg13g2_fill_1 FILLER_29_259 ();
 sg13g2_fill_2 FILLER_29_266 ();
 sg13g2_fill_1 FILLER_29_268 ();
 sg13g2_decap_8 FILLER_29_273 ();
 sg13g2_decap_4 FILLER_29_280 ();
 sg13g2_fill_1 FILLER_29_284 ();
 sg13g2_decap_4 FILLER_29_297 ();
 sg13g2_decap_8 FILLER_29_311 ();
 sg13g2_fill_2 FILLER_29_318 ();
 sg13g2_fill_1 FILLER_29_320 ();
 sg13g2_decap_4 FILLER_29_331 ();
 sg13g2_fill_1 FILLER_29_335 ();
 sg13g2_decap_8 FILLER_29_341 ();
 sg13g2_decap_8 FILLER_29_351 ();
 sg13g2_fill_2 FILLER_29_358 ();
 sg13g2_fill_1 FILLER_29_360 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_7 ();
 sg13g2_fill_1 FILLER_30_9 ();
 sg13g2_decap_4 FILLER_30_40 ();
 sg13g2_fill_1 FILLER_30_59 ();
 sg13g2_decap_4 FILLER_30_64 ();
 sg13g2_fill_2 FILLER_30_68 ();
 sg13g2_decap_8 FILLER_30_75 ();
 sg13g2_decap_4 FILLER_30_82 ();
 sg13g2_fill_1 FILLER_30_86 ();
 sg13g2_fill_1 FILLER_30_139 ();
 sg13g2_fill_2 FILLER_30_146 ();
 sg13g2_fill_1 FILLER_30_159 ();
 sg13g2_fill_1 FILLER_30_172 ();
 sg13g2_fill_1 FILLER_30_179 ();
 sg13g2_fill_1 FILLER_30_203 ();
 sg13g2_fill_1 FILLER_30_214 ();
 sg13g2_decap_4 FILLER_30_220 ();
 sg13g2_fill_1 FILLER_30_224 ();
 sg13g2_decap_8 FILLER_30_235 ();
 sg13g2_fill_2 FILLER_30_242 ();
 sg13g2_fill_1 FILLER_30_244 ();
 sg13g2_fill_1 FILLER_30_256 ();
 sg13g2_decap_8 FILLER_30_278 ();
 sg13g2_fill_2 FILLER_30_285 ();
 sg13g2_fill_1 FILLER_30_287 ();
 sg13g2_fill_2 FILLER_30_291 ();
 sg13g2_decap_8 FILLER_30_313 ();
 sg13g2_fill_1 FILLER_30_348 ();
 sg13g2_fill_2 FILLER_30_363 ();
 sg13g2_fill_2 FILLER_30_383 ();
 sg13g2_decap_4 FILLER_30_390 ();
 sg13g2_fill_1 FILLER_30_394 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_fill_1 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_29 ();
 sg13g2_fill_1 FILLER_31_36 ();
 sg13g2_fill_2 FILLER_31_45 ();
 sg13g2_fill_2 FILLER_31_73 ();
 sg13g2_fill_2 FILLER_31_91 ();
 sg13g2_fill_1 FILLER_31_93 ();
 sg13g2_decap_8 FILLER_31_108 ();
 sg13g2_decap_8 FILLER_31_115 ();
 sg13g2_decap_8 FILLER_31_122 ();
 sg13g2_fill_2 FILLER_31_134 ();
 sg13g2_fill_2 FILLER_31_145 ();
 sg13g2_fill_1 FILLER_31_147 ();
 sg13g2_decap_4 FILLER_31_157 ();
 sg13g2_fill_1 FILLER_31_167 ();
 sg13g2_decap_4 FILLER_31_181 ();
 sg13g2_fill_2 FILLER_31_185 ();
 sg13g2_decap_8 FILLER_31_196 ();
 sg13g2_decap_8 FILLER_31_209 ();
 sg13g2_decap_8 FILLER_31_216 ();
 sg13g2_decap_8 FILLER_31_223 ();
 sg13g2_decap_8 FILLER_31_239 ();
 sg13g2_decap_8 FILLER_31_246 ();
 sg13g2_fill_2 FILLER_31_253 ();
 sg13g2_fill_1 FILLER_31_255 ();
 sg13g2_fill_1 FILLER_31_264 ();
 sg13g2_decap_8 FILLER_31_271 ();
 sg13g2_fill_2 FILLER_31_278 ();
 sg13g2_fill_1 FILLER_31_283 ();
 sg13g2_decap_8 FILLER_31_319 ();
 sg13g2_fill_1 FILLER_31_326 ();
 sg13g2_fill_2 FILLER_31_332 ();
 sg13g2_fill_1 FILLER_31_334 ();
 sg13g2_fill_2 FILLER_31_353 ();
 sg13g2_fill_1 FILLER_31_355 ();
 sg13g2_decap_8 FILLER_31_391 ();
 sg13g2_decap_8 FILLER_31_398 ();
 sg13g2_decap_4 FILLER_31_405 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_52 ();
 sg13g2_decap_8 FILLER_32_59 ();
 sg13g2_fill_1 FILLER_32_66 ();
 sg13g2_fill_1 FILLER_32_93 ();
 sg13g2_fill_2 FILLER_32_133 ();
 sg13g2_fill_1 FILLER_32_164 ();
 sg13g2_fill_2 FILLER_32_194 ();
 sg13g2_decap_4 FILLER_32_218 ();
 sg13g2_fill_2 FILLER_32_222 ();
 sg13g2_decap_8 FILLER_32_241 ();
 sg13g2_decap_4 FILLER_32_248 ();
 sg13g2_fill_2 FILLER_32_252 ();
 sg13g2_fill_2 FILLER_32_270 ();
 sg13g2_fill_2 FILLER_32_280 ();
 sg13g2_fill_1 FILLER_32_299 ();
 sg13g2_fill_2 FILLER_32_342 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_4 FILLER_33_28 ();
 sg13g2_fill_1 FILLER_33_32 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_64 ();
 sg13g2_decap_4 FILLER_33_71 ();
 sg13g2_fill_1 FILLER_33_75 ();
 sg13g2_fill_2 FILLER_33_90 ();
 sg13g2_fill_1 FILLER_33_92 ();
 sg13g2_decap_8 FILLER_33_102 ();
 sg13g2_decap_8 FILLER_33_109 ();
 sg13g2_decap_8 FILLER_33_116 ();
 sg13g2_fill_1 FILLER_33_123 ();
 sg13g2_fill_2 FILLER_33_138 ();
 sg13g2_fill_1 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_151 ();
 sg13g2_fill_2 FILLER_33_158 ();
 sg13g2_decap_8 FILLER_33_179 ();
 sg13g2_decap_8 FILLER_33_186 ();
 sg13g2_fill_2 FILLER_33_193 ();
 sg13g2_fill_1 FILLER_33_195 ();
 sg13g2_decap_8 FILLER_33_206 ();
 sg13g2_decap_8 FILLER_33_213 ();
 sg13g2_decap_4 FILLER_33_220 ();
 sg13g2_decap_8 FILLER_33_238 ();
 sg13g2_fill_2 FILLER_33_245 ();
 sg13g2_fill_1 FILLER_33_247 ();
 sg13g2_decap_8 FILLER_33_252 ();
 sg13g2_fill_2 FILLER_33_259 ();
 sg13g2_fill_2 FILLER_33_304 ();
 sg13g2_fill_1 FILLER_33_306 ();
 sg13g2_decap_8 FILLER_33_312 ();
 sg13g2_decap_4 FILLER_33_319 ();
 sg13g2_fill_2 FILLER_33_336 ();
 sg13g2_fill_2 FILLER_33_352 ();
 sg13g2_fill_2 FILLER_33_380 ();
 sg13g2_fill_1 FILLER_33_382 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_fill_2 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_44 ();
 sg13g2_decap_4 FILLER_34_51 ();
 sg13g2_fill_2 FILLER_34_55 ();
 sg13g2_decap_8 FILLER_34_83 ();
 sg13g2_decap_8 FILLER_34_90 ();
 sg13g2_decap_8 FILLER_34_97 ();
 sg13g2_decap_8 FILLER_34_104 ();
 sg13g2_decap_8 FILLER_34_111 ();
 sg13g2_fill_1 FILLER_34_118 ();
 sg13g2_fill_1 FILLER_34_123 ();
 sg13g2_decap_8 FILLER_34_141 ();
 sg13g2_fill_1 FILLER_34_148 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_4 FILLER_34_161 ();
 sg13g2_decap_4 FILLER_34_176 ();
 sg13g2_fill_2 FILLER_34_180 ();
 sg13g2_fill_1 FILLER_34_188 ();
 sg13g2_decap_8 FILLER_34_211 ();
 sg13g2_fill_2 FILLER_34_218 ();
 sg13g2_fill_1 FILLER_34_220 ();
 sg13g2_decap_8 FILLER_34_227 ();
 sg13g2_fill_1 FILLER_34_234 ();
 sg13g2_fill_1 FILLER_34_284 ();
 sg13g2_decap_8 FILLER_34_293 ();
 sg13g2_fill_2 FILLER_34_300 ();
 sg13g2_fill_1 FILLER_34_351 ();
 sg13g2_fill_1 FILLER_34_360 ();
 sg13g2_decap_8 FILLER_34_367 ();
 sg13g2_decap_8 FILLER_34_374 ();
 sg13g2_fill_2 FILLER_34_381 ();
 sg13g2_decap_4 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_4 ();
 sg13g2_decap_4 FILLER_35_31 ();
 sg13g2_decap_8 FILLER_35_61 ();
 sg13g2_decap_8 FILLER_35_68 ();
 sg13g2_fill_1 FILLER_35_75 ();
 sg13g2_decap_8 FILLER_35_83 ();
 sg13g2_decap_8 FILLER_35_90 ();
 sg13g2_fill_2 FILLER_35_97 ();
 sg13g2_fill_2 FILLER_35_125 ();
 sg13g2_fill_1 FILLER_35_136 ();
 sg13g2_fill_2 FILLER_35_162 ();
 sg13g2_fill_1 FILLER_35_183 ();
 sg13g2_decap_8 FILLER_35_204 ();
 sg13g2_decap_8 FILLER_35_211 ();
 sg13g2_fill_1 FILLER_35_218 ();
 sg13g2_fill_1 FILLER_35_224 ();
 sg13g2_fill_2 FILLER_35_261 ();
 sg13g2_fill_1 FILLER_35_263 ();
 sg13g2_fill_1 FILLER_35_325 ();
 sg13g2_decap_4 FILLER_35_334 ();
 sg13g2_decap_8 FILLER_35_364 ();
 sg13g2_decap_8 FILLER_35_371 ();
 sg13g2_fill_2 FILLER_35_378 ();
 sg13g2_fill_1 FILLER_35_380 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_fill_1 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_34 ();
 sg13g2_decap_8 FILLER_36_41 ();
 sg13g2_decap_8 FILLER_36_48 ();
 sg13g2_decap_8 FILLER_36_55 ();
 sg13g2_decap_8 FILLER_36_62 ();
 sg13g2_decap_8 FILLER_36_69 ();
 sg13g2_decap_8 FILLER_36_76 ();
 sg13g2_decap_8 FILLER_36_83 ();
 sg13g2_decap_8 FILLER_36_90 ();
 sg13g2_decap_8 FILLER_36_97 ();
 sg13g2_decap_8 FILLER_36_104 ();
 sg13g2_decap_4 FILLER_36_111 ();
 sg13g2_fill_2 FILLER_36_115 ();
 sg13g2_fill_2 FILLER_36_149 ();
 sg13g2_fill_1 FILLER_36_160 ();
 sg13g2_decap_4 FILLER_36_177 ();
 sg13g2_fill_1 FILLER_36_181 ();
 sg13g2_fill_1 FILLER_36_186 ();
 sg13g2_fill_1 FILLER_36_191 ();
 sg13g2_fill_2 FILLER_36_209 ();
 sg13g2_fill_1 FILLER_36_246 ();
 sg13g2_fill_1 FILLER_36_256 ();
 sg13g2_decap_8 FILLER_36_281 ();
 sg13g2_decap_8 FILLER_36_288 ();
 sg13g2_decap_8 FILLER_36_295 ();
 sg13g2_fill_1 FILLER_36_302 ();
 sg13g2_decap_8 FILLER_36_329 ();
 sg13g2_decap_8 FILLER_36_340 ();
 sg13g2_decap_8 FILLER_36_388 ();
 sg13g2_decap_4 FILLER_36_395 ();
 sg13g2_fill_1 FILLER_36_399 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_4 FILLER_37_112 ();
 sg13g2_fill_1 FILLER_37_116 ();
 sg13g2_fill_2 FILLER_37_179 ();
 sg13g2_fill_1 FILLER_37_181 ();
 sg13g2_fill_2 FILLER_37_210 ();
 sg13g2_fill_2 FILLER_37_220 ();
 sg13g2_fill_1 FILLER_37_222 ();
 sg13g2_fill_1 FILLER_37_231 ();
 sg13g2_fill_1 FILLER_37_258 ();
 sg13g2_decap_8 FILLER_37_316 ();
 sg13g2_decap_4 FILLER_37_323 ();
 sg13g2_fill_1 FILLER_37_327 ();
 sg13g2_decap_4 FILLER_37_354 ();
 sg13g2_fill_1 FILLER_37_358 ();
 sg13g2_decap_8 FILLER_37_385 ();
 sg13g2_decap_4 FILLER_37_392 ();
 sg13g2_fill_1 FILLER_37_396 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_8 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_107 ();
 sg13g2_fill_1 FILLER_38_111 ();
 sg13g2_decap_8 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_123 ();
 sg13g2_fill_1 FILLER_38_127 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_fill_2 FILLER_38_136 ();
 sg13g2_decap_4 FILLER_38_155 ();
 sg13g2_fill_1 FILLER_38_159 ();
 sg13g2_decap_8 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_171 ();
 sg13g2_fill_1 FILLER_38_297 ();
 sg13g2_decap_4 FILLER_38_307 ();
 sg13g2_fill_1 FILLER_38_311 ();
 sg13g2_decap_4 FILLER_38_316 ();
 sg13g2_fill_2 FILLER_38_324 ();
 sg13g2_fill_1 FILLER_38_368 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net22;
 assign uio_oe[2] = net10;
 assign uio_oe[3] = net23;
 assign uio_oe[4] = net24;
 assign uio_oe[5] = net25;
 assign uio_oe[6] = net11;
 assign uio_oe[7] = net26;
 assign uio_out[2] = net12;
 assign uio_out[4] = net27;
 assign uio_out[6] = net13;
 assign uo_out[0] = net14;
 assign uo_out[1] = net15;
 assign uo_out[2] = net16;
 assign uo_out[3] = net17;
 assign uo_out[4] = net18;
 assign uo_out[5] = net19;
 assign uo_out[6] = net20;
 assign uo_out[7] = net21;
endmodule
