module tt_um_wokwi_434917577229968385 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire params_ready;
 wire spike_out;
 wire \system_inst.leak_cycles[0] ;
 wire \system_inst.leak_cycles[1] ;
 wire \system_inst.leak_cycles[2] ;
 wire \system_inst.leak_cycles[3] ;
 wire \system_inst.leak_rate[0] ;
 wire \system_inst.leak_rate[1] ;
 wire \system_inst.leak_rate[2] ;
 wire \system_inst.leak_rate[3] ;
 wire \system_inst.leak_rate[4] ;
 wire \system_inst.leak_rate[5] ;
 wire \system_inst.leak_rate[6] ;
 wire \system_inst.leak_rate[7] ;
 wire \system_inst.loader.bit_count[0] ;
 wire \system_inst.loader.bit_count[1] ;
 wire \system_inst.loader.bit_count[2] ;
 wire \system_inst.loader.current_state[0] ;
 wire \system_inst.loader.current_state[1] ;
 wire \system_inst.loader.current_state[2] ;
 wire \system_inst.loader.current_state[4] ;
 wire \system_inst.loader.current_state[5] ;
 wire \system_inst.loader.current_state[6] ;
 wire \system_inst.loader.shift_reg[0] ;
 wire \system_inst.loader.shift_reg[1] ;
 wire \system_inst.loader.shift_reg[2] ;
 wire \system_inst.loader.shift_reg[3] ;
 wire \system_inst.loader.shift_reg[4] ;
 wire \system_inst.loader.shift_reg[5] ;
 wire \system_inst.loader.shift_reg[6] ;
 wire \system_inst.loader.threshold[0] ;
 wire \system_inst.loader.threshold[1] ;
 wire \system_inst.loader.threshold[2] ;
 wire \system_inst.loader.threshold[3] ;
 wire \system_inst.loader.threshold[4] ;
 wire \system_inst.loader.threshold[5] ;
 wire \system_inst.loader.threshold[6] ;
 wire \system_inst.loader.threshold[7] ;
 wire \system_inst.loader.weight_a[0] ;
 wire \system_inst.loader.weight_a[1] ;
 wire \system_inst.loader.weight_a[2] ;
 wire \system_inst.loader.weight_b[0] ;
 wire \system_inst.loader.weight_b[1] ;
 wire \system_inst.loader.weight_b[2] ;
 wire \system_inst.neuron.leak_counter[0] ;
 wire \system_inst.neuron.leak_counter[1] ;
 wire \system_inst.neuron.leak_counter[2] ;
 wire \system_inst.neuron.leak_counter[3] ;
 wire \system_inst.neuron.refr_cnt[0] ;
 wire \system_inst.neuron.refr_cnt[1] ;
 wire \system_inst.neuron.refr_cnt[2] ;
 wire \system_inst.neuron.refr_cnt[3] ;
 wire \system_inst.neuron.v_mem[0] ;
 wire \system_inst.neuron.v_mem[1] ;
 wire \system_inst.neuron.v_mem[2] ;
 wire \system_inst.neuron.v_mem[3] ;
 wire \system_inst.neuron.v_mem[4] ;
 wire \system_inst.neuron.v_mem[5] ;
 wire \system_inst.neuron.v_mem[6] ;
 wire \system_inst.neuron.v_mem[7] ;
 wire \system_inst.neuron.v_mem[8] ;
 wire clknet_0_clk;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;

 sg13g2_inv_1 _0534_ (.Y(_0066_),
    .A(net138));
 sg13g2_inv_1 _0535_ (.Y(_0067_),
    .A(net127));
 sg13g2_inv_1 _0536_ (.Y(_0068_),
    .A(net148));
 sg13g2_inv_1 _0537_ (.Y(_0069_),
    .A(net125));
 sg13g2_inv_1 _0538_ (.Y(_0070_),
    .A(net137));
 sg13g2_inv_1 _0539_ (.Y(_0071_),
    .A(net133));
 sg13g2_inv_2 _0540_ (.Y(_0072_),
    .A(net168));
 sg13g2_inv_1 _0541_ (.Y(_0073_),
    .A(\system_inst.loader.shift_reg[0] ));
 sg13g2_inv_1 _0542_ (.Y(_0074_),
    .A(\system_inst.leak_cycles[2] ));
 sg13g2_inv_1 _0543_ (.Y(_0075_),
    .A(net121));
 sg13g2_inv_2 _0544_ (.Y(_0076_),
    .A(net4));
 sg13g2_inv_1 _0545_ (.Y(_0077_),
    .A(net144));
 sg13g2_inv_1 _0546_ (.Y(_0078_),
    .A(net142));
 sg13g2_inv_1 _0547_ (.Y(_0079_),
    .A(\system_inst.leak_rate[2] ));
 sg13g2_inv_1 _0548_ (.Y(_0080_),
    .A(net150));
 sg13g2_inv_1 _0549_ (.Y(_0081_),
    .A(net118));
 sg13g2_inv_1 _0550_ (.Y(_0082_),
    .A(net193));
 sg13g2_inv_1 _0551_ (.Y(_0083_),
    .A(net189));
 sg13g2_inv_1 _0552_ (.Y(_0084_),
    .A(net195));
 sg13g2_inv_1 _0553_ (.Y(_0085_),
    .A(_0007_));
 sg13g2_inv_1 _0554_ (.Y(_0086_),
    .A(_0008_));
 sg13g2_inv_1 _0555_ (.Y(_0087_),
    .A(net101));
 sg13g2_inv_1 _0556_ (.Y(_0088_),
    .A(net124));
 sg13g2_inv_1 _0557_ (.Y(_0089_),
    .A(\system_inst.loader.current_state[0] ));
 sg13g2_nand2b_1 _0558_ (.Y(_0090_),
    .B(net99),
    .A_N(net1));
 sg13g2_nand2_1 _0559_ (.Y(_0091_),
    .A(net169),
    .B(net138));
 sg13g2_nor2_1 _0560_ (.A(_0009_),
    .B(_0091_),
    .Y(_0092_));
 sg13g2_inv_1 _0561_ (.Y(_0093_),
    .A(net91));
 sg13g2_and2_2 _0562_ (.A(net3),
    .B(net1),
    .X(_0094_));
 sg13g2_nand2_1 _0563_ (.Y(_0095_),
    .A(net101),
    .B(_0094_));
 sg13g2_o21ai_1 _0564_ (.B1(_0090_),
    .Y(_0096_),
    .A1(net91),
    .A2(_0095_));
 sg13g2_and3_1 _0565_ (.X(_0097_),
    .A(net139),
    .B(_0092_),
    .C(_0094_));
 sg13g2_a22oi_1 _0566_ (.Y(_0098_),
    .B1(_0097_),
    .B2(net101),
    .A2(_0096_),
    .A1(net163));
 sg13g2_inv_1 _0567_ (.Y(_0001_),
    .A(net164));
 sg13g2_nand3_1 _0568_ (.B(net91),
    .C(_0094_),
    .A(net141),
    .Y(_0099_));
 sg13g2_inv_2 _0569_ (.Y(_0100_),
    .A(_0099_));
 sg13g2_a22oi_1 _0570_ (.Y(_0101_),
    .B1(_0100_),
    .B2(net101),
    .A2(_0096_),
    .A1(net139));
 sg13g2_inv_1 _0571_ (.Y(_0005_),
    .A(net140));
 sg13g2_nor2_1 _0572_ (.A(net123),
    .B(_0090_),
    .Y(_0102_));
 sg13g2_a21oi_1 _0573_ (.A1(net99),
    .A2(_0094_),
    .Y(_0000_),
    .B1(_0102_));
 sg13g2_nand3_1 _0574_ (.B(net91),
    .C(_0094_),
    .A(net116),
    .Y(_0103_));
 sg13g2_inv_2 _0575_ (.Y(_0104_),
    .A(_0103_));
 sg13g2_a22oi_1 _0576_ (.Y(_0105_),
    .B1(_0104_),
    .B2(net101),
    .A2(_0096_),
    .A1(net141));
 sg13g2_inv_1 _0577_ (.Y(_0002_),
    .A(_0105_));
 sg13g2_nand2_1 _0578_ (.Y(_0106_),
    .A(net116),
    .B(_0096_));
 sg13g2_o21ai_1 _0579_ (.B1(_0106_),
    .Y(_0003_),
    .A1(_0089_),
    .A2(_0095_));
 sg13g2_and3_1 _0580_ (.X(_0107_),
    .A(\system_inst.loader.current_state[1] ),
    .B(_0092_),
    .C(_0094_));
 sg13g2_nand3_1 _0581_ (.B(net91),
    .C(_0094_),
    .A(\system_inst.loader.current_state[1] ),
    .Y(_0108_));
 sg13g2_a22oi_1 _0582_ (.Y(_0109_),
    .B1(net88),
    .B2(net100),
    .A2(_0096_),
    .A1(net124));
 sg13g2_inv_1 _0583_ (.Y(_0004_),
    .A(_0109_));
 sg13g2_nor2b_1 _0584_ (.A(net92),
    .B_N(\system_inst.neuron.v_mem[0] ),
    .Y(uo_out[1]));
 sg13g2_nor2b_1 _0585_ (.A(net92),
    .B_N(\system_inst.neuron.v_mem[1] ),
    .Y(uo_out[2]));
 sg13g2_nor2b_1 _0586_ (.A(net92),
    .B_N(\system_inst.neuron.v_mem[2] ),
    .Y(uo_out[3]));
 sg13g2_nor2b_1 _0587_ (.A(net92),
    .B_N(\system_inst.neuron.v_mem[3] ),
    .Y(uo_out[4]));
 sg13g2_nor2b_1 _0588_ (.A(\system_inst.neuron.v_mem[8] ),
    .B_N(\system_inst.neuron.v_mem[4] ),
    .Y(uo_out[5]));
 sg13g2_nor2b_1 _0589_ (.A(net92),
    .B_N(\system_inst.neuron.v_mem[5] ),
    .Y(uo_out[6]));
 sg13g2_nor2b_1 _0590_ (.A(net92),
    .B_N(\system_inst.neuron.v_mem[6] ),
    .Y(uo_out[7]));
 sg13g2_nor2_1 _0591_ (.A(net197),
    .B(\system_inst.neuron.refr_cnt[0] ),
    .Y(_0110_));
 sg13g2_nor4_2 _0592_ (.A(net112),
    .B(\system_inst.neuron.refr_cnt[2] ),
    .C(\system_inst.neuron.refr_cnt[1] ),
    .Y(_0111_),
    .D(\system_inst.neuron.refr_cnt[0] ));
 sg13g2_nand2_2 _0593_ (.Y(_0112_),
    .A(net170),
    .B(net1));
 sg13g2_inv_1 _0594_ (.Y(_0113_),
    .A(_0112_));
 sg13g2_nand2_1 _0595_ (.Y(_0114_),
    .A(net2),
    .B(_0113_));
 sg13g2_nand3_1 _0596_ (.B(_0111_),
    .C(_0113_),
    .A(net2),
    .Y(_0115_));
 sg13g2_nand2_1 _0597_ (.Y(_0116_),
    .A(\system_inst.loader.weight_a[1] ),
    .B(net6));
 sg13g2_nand3_1 _0598_ (.B(net7),
    .C(_0116_),
    .A(\system_inst.loader.weight_a[2] ),
    .Y(_0117_));
 sg13g2_nand2_1 _0599_ (.Y(_0118_),
    .A(\system_inst.loader.weight_a[2] ),
    .B(net6));
 sg13g2_and4_1 _0600_ (.A(\system_inst.loader.weight_a[2] ),
    .B(\system_inst.loader.weight_a[1] ),
    .C(net5),
    .D(net6),
    .X(_0119_));
 sg13g2_nand4_1 _0601_ (.B(\system_inst.loader.weight_a[1] ),
    .C(net5),
    .A(\system_inst.loader.weight_a[2] ),
    .Y(_0120_),
    .D(net6));
 sg13g2_nand2_1 _0602_ (.Y(_0121_),
    .A(\system_inst.loader.weight_a[0] ),
    .B(net7));
 sg13g2_a22oi_1 _0603_ (.Y(_0122_),
    .B1(net6),
    .B2(\system_inst.loader.weight_a[1] ),
    .A2(net5),
    .A1(\system_inst.loader.weight_a[2] ));
 sg13g2_or3_1 _0604_ (.A(_0119_),
    .B(_0121_),
    .C(_0122_),
    .X(_0123_));
 sg13g2_o21ai_1 _0605_ (.B1(_0120_),
    .Y(_0124_),
    .A1(_0121_),
    .A2(_0122_));
 sg13g2_nand2_1 _0606_ (.Y(_0125_),
    .A(\system_inst.loader.weight_a[1] ),
    .B(net7));
 sg13g2_xor2_1 _0607_ (.B(_0125_),
    .A(_0118_),
    .X(_0126_));
 sg13g2_nand2_1 _0608_ (.Y(_0127_),
    .A(_0124_),
    .B(_0126_));
 sg13g2_nand2_1 _0609_ (.Y(_0128_),
    .A(\system_inst.loader.weight_a[0] ),
    .B(net5));
 sg13g2_and4_1 _0610_ (.A(\system_inst.loader.weight_a[1] ),
    .B(\system_inst.loader.weight_a[0] ),
    .C(net5),
    .D(net6),
    .X(_0129_));
 sg13g2_o21ai_1 _0611_ (.B1(_0121_),
    .Y(_0130_),
    .A1(_0119_),
    .A2(_0122_));
 sg13g2_nand3_1 _0612_ (.B(_0129_),
    .C(_0130_),
    .A(_0123_),
    .Y(_0131_));
 sg13g2_xnor2_1 _0613_ (.Y(_0132_),
    .A(_0124_),
    .B(_0126_));
 sg13g2_o21ai_1 _0614_ (.B1(_0127_),
    .Y(_0133_),
    .A1(_0131_),
    .A2(_0132_));
 sg13g2_nand2b_1 _0615_ (.Y(_0134_),
    .B(_0133_),
    .A_N(_0117_));
 sg13g2_xnor2_1 _0616_ (.Y(_0135_),
    .A(_0117_),
    .B(_0133_));
 sg13g2_nand2_1 _0617_ (.Y(_0136_),
    .A(\system_inst.neuron.v_mem[4] ),
    .B(_0135_));
 sg13g2_nand2_2 _0618_ (.Y(_0137_),
    .A(\system_inst.loader.weight_b[1] ),
    .B(net8));
 sg13g2_nand2_1 _0619_ (.Y(_0138_),
    .A(\system_inst.loader.weight_b[2] ),
    .B(net9));
 sg13g2_nand2b_1 _0620_ (.Y(_0139_),
    .B(_0137_),
    .A_N(_0138_));
 sg13g2_nand2_1 _0621_ (.Y(_0140_),
    .A(\system_inst.loader.weight_b[2] ),
    .B(net8));
 sg13g2_nand2_1 _0622_ (.Y(_0141_),
    .A(\system_inst.loader.weight_b[1] ),
    .B(net9));
 sg13g2_xor2_1 _0623_ (.B(_0141_),
    .A(_0140_),
    .X(_0142_));
 sg13g2_a22oi_1 _0624_ (.Y(_0143_),
    .B1(net9),
    .B2(\system_inst.loader.weight_b[0] ),
    .A2(net10),
    .A1(\system_inst.loader.weight_b[2] ));
 sg13g2_nand2_2 _0625_ (.Y(_0144_),
    .A(\system_inst.loader.weight_b[0] ),
    .B(net10));
 sg13g2_nand4_1 _0626_ (.B(\system_inst.loader.weight_b[0] ),
    .C(net10),
    .A(\system_inst.loader.weight_b[2] ),
    .Y(_0145_),
    .D(net9));
 sg13g2_o21ai_1 _0627_ (.B1(_0145_),
    .Y(_0146_),
    .A1(_0137_),
    .A2(_0143_));
 sg13g2_nor2b_1 _0628_ (.A(_0143_),
    .B_N(_0145_),
    .Y(_0147_));
 sg13g2_nor3_1 _0629_ (.A(_0137_),
    .B(_0144_),
    .C(_0147_),
    .Y(_0148_));
 sg13g2_xnor2_1 _0630_ (.Y(_0149_),
    .A(_0142_),
    .B(_0146_));
 sg13g2_nor4_1 _0631_ (.A(_0137_),
    .B(_0144_),
    .C(_0147_),
    .D(_0149_),
    .Y(_0150_));
 sg13g2_a21oi_2 _0632_ (.B1(_0150_),
    .Y(_0151_),
    .A2(_0146_),
    .A1(_0142_));
 sg13g2_xor2_1 _0633_ (.B(_0151_),
    .A(_0139_),
    .X(_0152_));
 sg13g2_xnor2_1 _0634_ (.Y(_0153_),
    .A(\system_inst.neuron.v_mem[4] ),
    .B(_0135_));
 sg13g2_o21ai_1 _0635_ (.B1(_0136_),
    .Y(_0154_),
    .A1(_0152_),
    .A2(_0153_));
 sg13g2_a21oi_2 _0636_ (.B1(_0138_),
    .Y(_0155_),
    .A2(_0151_),
    .A1(_0137_));
 sg13g2_o21ai_1 _0637_ (.B1(_0134_),
    .Y(_0156_),
    .A1(_0118_),
    .A2(_0125_));
 sg13g2_xor2_1 _0638_ (.B(_0156_),
    .A(\system_inst.neuron.v_mem[5] ),
    .X(_0157_));
 sg13g2_nor2b_1 _0639_ (.A(_0155_),
    .B_N(_0157_),
    .Y(_0158_));
 sg13g2_xnor2_1 _0640_ (.Y(_0159_),
    .A(_0155_),
    .B(_0157_));
 sg13g2_nand2_1 _0641_ (.Y(_0160_),
    .A(_0154_),
    .B(_0159_));
 sg13g2_xor2_1 _0642_ (.B(_0132_),
    .A(_0131_),
    .X(_0161_));
 sg13g2_xor2_1 _0643_ (.B(_0149_),
    .A(_0148_),
    .X(_0162_));
 sg13g2_xnor2_1 _0644_ (.Y(_0163_),
    .A(\system_inst.neuron.v_mem[3] ),
    .B(_0161_));
 sg13g2_nor2b_1 _0645_ (.A(_0163_),
    .B_N(_0162_),
    .Y(_0164_));
 sg13g2_a21o_1 _0646_ (.A2(_0161_),
    .A1(\system_inst.neuron.v_mem[3] ),
    .B1(_0164_),
    .X(_0165_));
 sg13g2_xor2_1 _0647_ (.B(_0153_),
    .A(_0152_),
    .X(_0166_));
 sg13g2_and2_1 _0648_ (.A(_0165_),
    .B(_0166_),
    .X(_0167_));
 sg13g2_a21o_1 _0649_ (.A2(_0130_),
    .A1(_0123_),
    .B1(_0129_),
    .X(_0168_));
 sg13g2_nand3_1 _0650_ (.B(_0131_),
    .C(_0168_),
    .A(\system_inst.neuron.v_mem[2] ),
    .Y(_0169_));
 sg13g2_a21o_1 _0651_ (.A2(_0168_),
    .A1(_0131_),
    .B1(\system_inst.neuron.v_mem[2] ),
    .X(_0170_));
 sg13g2_nor2b_1 _0652_ (.A(_0137_),
    .B_N(_0144_),
    .Y(_0171_));
 sg13g2_xnor2_1 _0653_ (.Y(_0172_),
    .A(_0147_),
    .B(_0171_));
 sg13g2_nand3_1 _0654_ (.B(_0170_),
    .C(_0172_),
    .A(_0169_),
    .Y(_0173_));
 sg13g2_nand2_1 _0655_ (.Y(_0174_),
    .A(_0169_),
    .B(_0173_));
 sg13g2_xor2_1 _0656_ (.B(_0163_),
    .A(_0162_),
    .X(_0175_));
 sg13g2_nor2b_1 _0657_ (.A(_0175_),
    .B_N(_0174_),
    .Y(_0176_));
 sg13g2_a22oi_1 _0658_ (.Y(_0177_),
    .B1(net6),
    .B2(\system_inst.loader.weight_a[0] ),
    .A2(net5),
    .A1(\system_inst.loader.weight_a[1] ));
 sg13g2_nor2_1 _0659_ (.A(_0129_),
    .B(_0177_),
    .Y(_0178_));
 sg13g2_a22oi_1 _0660_ (.Y(_0179_),
    .B1(net8),
    .B2(\system_inst.loader.weight_b[0] ),
    .A2(net10),
    .A1(\system_inst.loader.weight_b[1] ));
 sg13g2_inv_1 _0661_ (.Y(_0180_),
    .A(_0179_));
 sg13g2_o21ai_1 _0662_ (.B1(_0180_),
    .Y(_0181_),
    .A1(_0137_),
    .A2(_0144_));
 sg13g2_xnor2_1 _0663_ (.Y(_0182_),
    .A(\system_inst.neuron.v_mem[1] ),
    .B(_0178_));
 sg13g2_nor2b_1 _0664_ (.A(_0182_),
    .B_N(_0181_),
    .Y(_0183_));
 sg13g2_a21o_1 _0665_ (.A2(_0178_),
    .A1(\system_inst.neuron.v_mem[1] ),
    .B1(_0183_),
    .X(_0184_));
 sg13g2_a21o_1 _0666_ (.A2(_0170_),
    .A1(_0169_),
    .B1(_0172_),
    .X(_0185_));
 sg13g2_and3_1 _0667_ (.X(_0186_),
    .A(_0173_),
    .B(_0184_),
    .C(_0185_));
 sg13g2_nand3_1 _0668_ (.B(_0184_),
    .C(_0185_),
    .A(_0173_),
    .Y(_0187_));
 sg13g2_nor2_1 _0669_ (.A(\system_inst.neuron.v_mem[0] ),
    .B(_0144_),
    .Y(_0188_));
 sg13g2_xnor2_1 _0670_ (.Y(_0189_),
    .A(_0181_),
    .B(_0182_));
 sg13g2_nor2b_1 _0671_ (.A(_0188_),
    .B_N(_0189_),
    .Y(_0190_));
 sg13g2_xor2_1 _0672_ (.B(_0144_),
    .A(\system_inst.neuron.v_mem[0] ),
    .X(_0191_));
 sg13g2_nor2_1 _0673_ (.A(_0128_),
    .B(_0191_),
    .Y(_0192_));
 sg13g2_xnor2_1 _0674_ (.Y(_0193_),
    .A(_0188_),
    .B(_0189_));
 sg13g2_a21oi_1 _0675_ (.A1(_0192_),
    .A2(_0193_),
    .Y(_0194_),
    .B1(_0190_));
 sg13g2_a21oi_1 _0676_ (.A1(_0173_),
    .A2(_0185_),
    .Y(_0195_),
    .B1(_0184_));
 sg13g2_or3_1 _0677_ (.A(_0186_),
    .B(_0194_),
    .C(_0195_),
    .X(_0196_));
 sg13g2_o21ai_1 _0678_ (.B1(_0187_),
    .Y(_0197_),
    .A1(_0194_),
    .A2(_0195_));
 sg13g2_xnor2_1 _0679_ (.Y(_0198_),
    .A(_0174_),
    .B(_0175_));
 sg13g2_a21o_1 _0680_ (.A2(_0198_),
    .A1(_0197_),
    .B1(_0176_),
    .X(_0199_));
 sg13g2_xor2_1 _0681_ (.B(_0166_),
    .A(_0165_),
    .X(_0200_));
 sg13g2_a21oi_1 _0682_ (.A1(_0199_),
    .A2(_0200_),
    .Y(_0201_),
    .B1(_0167_));
 sg13g2_xnor2_1 _0683_ (.Y(_0202_),
    .A(_0154_),
    .B(_0159_));
 sg13g2_o21ai_1 _0684_ (.B1(_0160_),
    .Y(_0203_),
    .A1(_0201_),
    .A2(_0202_));
 sg13g2_a21o_1 _0685_ (.A2(_0156_),
    .A1(\system_inst.neuron.v_mem[5] ),
    .B1(_0158_),
    .X(_0204_));
 sg13g2_xor2_1 _0686_ (.B(_0156_),
    .A(\system_inst.neuron.v_mem[6] ),
    .X(_0205_));
 sg13g2_nor2b_1 _0687_ (.A(_0155_),
    .B_N(_0205_),
    .Y(_0206_));
 sg13g2_xnor2_1 _0688_ (.Y(_0207_),
    .A(_0155_),
    .B(_0205_));
 sg13g2_and2_1 _0689_ (.A(_0204_),
    .B(_0207_),
    .X(_0208_));
 sg13g2_or2_1 _0690_ (.X(_0209_),
    .B(_0207_),
    .A(_0204_));
 sg13g2_xor2_1 _0691_ (.B(_0207_),
    .A(_0204_),
    .X(_0210_));
 sg13g2_xnor2_1 _0692_ (.Y(_0211_),
    .A(_0203_),
    .B(_0210_));
 sg13g2_or2_1 _0693_ (.X(_0212_),
    .B(_0211_),
    .A(\system_inst.leak_rate[6] ));
 sg13g2_and2_1 _0694_ (.A(\system_inst.leak_rate[6] ),
    .B(_0211_),
    .X(_0213_));
 sg13g2_xor2_1 _0695_ (.B(_0211_),
    .A(\system_inst.leak_rate[6] ),
    .X(_0214_));
 sg13g2_xnor2_1 _0696_ (.Y(_0215_),
    .A(_0201_),
    .B(_0202_));
 sg13g2_nor2_1 _0697_ (.A(\system_inst.leak_rate[5] ),
    .B(_0215_),
    .Y(_0216_));
 sg13g2_xnor2_1 _0698_ (.Y(_0217_),
    .A(_0199_),
    .B(_0200_));
 sg13g2_or2_1 _0699_ (.X(_0218_),
    .B(_0217_),
    .A(\system_inst.leak_rate[4] ));
 sg13g2_and2_1 _0700_ (.A(\system_inst.leak_rate[4] ),
    .B(_0217_),
    .X(_0219_));
 sg13g2_xor2_1 _0701_ (.B(_0217_),
    .A(\system_inst.leak_rate[4] ),
    .X(_0220_));
 sg13g2_xnor2_1 _0702_ (.Y(_0221_),
    .A(_0197_),
    .B(_0198_));
 sg13g2_nor2_1 _0703_ (.A(\system_inst.leak_rate[3] ),
    .B(_0221_),
    .Y(_0222_));
 sg13g2_xor2_1 _0704_ (.B(_0221_),
    .A(\system_inst.leak_rate[3] ),
    .X(_0223_));
 sg13g2_o21ai_1 _0705_ (.B1(_0194_),
    .Y(_0224_),
    .A1(_0186_),
    .A2(_0195_));
 sg13g2_and2_1 _0706_ (.A(_0196_),
    .B(_0224_),
    .X(_0225_));
 sg13g2_nand3_1 _0707_ (.B(_0196_),
    .C(_0224_),
    .A(_0079_),
    .Y(_0226_));
 sg13g2_a21oi_1 _0708_ (.A1(_0196_),
    .A2(_0224_),
    .Y(_0227_),
    .B1(_0079_));
 sg13g2_xnor2_1 _0709_ (.Y(_0228_),
    .A(_0079_),
    .B(_0225_));
 sg13g2_xnor2_1 _0710_ (.Y(_0229_),
    .A(_0192_),
    .B(_0193_));
 sg13g2_nor2_1 _0711_ (.A(\system_inst.leak_rate[1] ),
    .B(_0229_),
    .Y(_0230_));
 sg13g2_xnor2_1 _0712_ (.Y(_0231_),
    .A(_0128_),
    .B(_0191_));
 sg13g2_nand2_1 _0713_ (.Y(_0232_),
    .A(\system_inst.leak_rate[0] ),
    .B(_0231_));
 sg13g2_xnor2_1 _0714_ (.Y(_0233_),
    .A(_0080_),
    .B(_0229_));
 sg13g2_a21oi_1 _0715_ (.A1(_0232_),
    .A2(_0233_),
    .Y(_0234_),
    .B1(_0230_));
 sg13g2_o21ai_1 _0716_ (.B1(_0226_),
    .Y(_0235_),
    .A1(_0227_),
    .A2(_0234_));
 sg13g2_a21oi_2 _0717_ (.B1(_0222_),
    .Y(_0236_),
    .A2(_0235_),
    .A1(_0223_));
 sg13g2_o21ai_1 _0718_ (.B1(_0218_),
    .Y(_0237_),
    .A1(_0219_),
    .A2(_0236_));
 sg13g2_xor2_1 _0719_ (.B(_0215_),
    .A(\system_inst.leak_rate[5] ),
    .X(_0238_));
 sg13g2_a21oi_1 _0720_ (.A1(_0237_),
    .A2(_0238_),
    .Y(_0239_),
    .B1(_0216_));
 sg13g2_o21ai_1 _0721_ (.B1(_0212_),
    .Y(_0240_),
    .A1(_0213_),
    .A2(_0239_));
 sg13g2_a21oi_1 _0722_ (.A1(_0203_),
    .A2(_0209_),
    .Y(_0241_),
    .B1(_0208_));
 sg13g2_a21o_1 _0723_ (.A2(_0156_),
    .A1(\system_inst.neuron.v_mem[6] ),
    .B1(_0206_),
    .X(_0242_));
 sg13g2_nand2_1 _0724_ (.Y(_0243_),
    .A(\system_inst.neuron.v_mem[7] ),
    .B(_0155_));
 sg13g2_nor2_1 _0725_ (.A(\system_inst.neuron.v_mem[7] ),
    .B(_0155_),
    .Y(_0244_));
 sg13g2_xor2_1 _0726_ (.B(_0155_),
    .A(\system_inst.neuron.v_mem[7] ),
    .X(_0245_));
 sg13g2_xnor2_1 _0727_ (.Y(_0246_),
    .A(_0156_),
    .B(_0245_));
 sg13g2_nand2_1 _0728_ (.Y(_0247_),
    .A(_0242_),
    .B(_0246_));
 sg13g2_xnor2_1 _0729_ (.Y(_0248_),
    .A(_0242_),
    .B(_0246_));
 sg13g2_xnor2_1 _0730_ (.Y(_0249_),
    .A(_0241_),
    .B(_0248_));
 sg13g2_xor2_1 _0731_ (.B(_0249_),
    .A(\system_inst.leak_rate[7] ),
    .X(_0250_));
 sg13g2_nand2b_1 _0732_ (.Y(_0251_),
    .B(\system_inst.neuron.leak_counter[3] ),
    .A_N(\system_inst.leak_cycles[3] ));
 sg13g2_a22oi_1 _0733_ (.Y(_0252_),
    .B1(_0082_),
    .B2(\system_inst.leak_cycles[0] ),
    .A2(_0081_),
    .A1(\system_inst.leak_cycles[1] ));
 sg13g2_a221oi_1 _0734_ (.B2(_0075_),
    .C1(_0252_),
    .B1(\system_inst.neuron.leak_counter[1] ),
    .A1(_0074_),
    .Y(_0253_),
    .A2(\system_inst.neuron.leak_counter[2] ));
 sg13g2_nand2b_1 _0735_ (.Y(_0254_),
    .B(\system_inst.leak_cycles[3] ),
    .A_N(\system_inst.neuron.leak_counter[3] ));
 sg13g2_o21ai_1 _0736_ (.B1(_0254_),
    .Y(_0255_),
    .A1(_0074_),
    .A2(\system_inst.neuron.leak_counter[2] ));
 sg13g2_o21ai_1 _0737_ (.B1(_0251_),
    .Y(_0256_),
    .A1(_0253_),
    .A2(_0255_));
 sg13g2_o21ai_1 _0738_ (.B1(net83),
    .Y(_0257_),
    .A1(\system_inst.leak_rate[7] ),
    .A2(_0249_));
 sg13g2_a21oi_2 _0739_ (.B1(_0257_),
    .Y(_0258_),
    .A2(_0250_),
    .A1(_0240_));
 sg13g2_o21ai_1 _0740_ (.B1(_0247_),
    .Y(_0259_),
    .A1(_0241_),
    .A2(_0248_));
 sg13g2_o21ai_1 _0741_ (.B1(_0243_),
    .Y(_0260_),
    .A1(_0156_),
    .A2(_0244_));
 sg13g2_xnor2_1 _0742_ (.Y(_0261_),
    .A(net92),
    .B(_0260_));
 sg13g2_xor2_1 _0743_ (.B(_0261_),
    .A(_0259_),
    .X(_0262_));
 sg13g2_xor2_1 _0744_ (.B(_0262_),
    .A(_0258_),
    .X(_0263_));
 sg13g2_xnor2_1 _0745_ (.Y(_0264_),
    .A(_0258_),
    .B(_0262_));
 sg13g2_xnor2_1 _0746_ (.Y(_0265_),
    .A(_0237_),
    .B(_0238_));
 sg13g2_mux2_1 _0747_ (.A0(_0215_),
    .A1(_0265_),
    .S(net83),
    .X(_0266_));
 sg13g2_nand2b_1 _0748_ (.Y(_0267_),
    .B(net80),
    .A_N(_0266_));
 sg13g2_or3_1 _0749_ (.A(\system_inst.loader.threshold[5] ),
    .B(_0263_),
    .C(_0266_),
    .X(_0268_));
 sg13g2_xnor2_1 _0750_ (.Y(_0269_),
    .A(_0214_),
    .B(_0239_));
 sg13g2_nand2_1 _0751_ (.Y(_0270_),
    .A(net83),
    .B(_0269_));
 sg13g2_o21ai_1 _0752_ (.B1(_0270_),
    .Y(_0271_),
    .A1(_0211_),
    .A2(net83));
 sg13g2_nand2_1 _0753_ (.Y(_0272_),
    .A(net80),
    .B(_0271_));
 sg13g2_nand3b_1 _0754_ (.B(net80),
    .C(_0271_),
    .Y(_0273_),
    .A_N(\system_inst.loader.threshold[6] ));
 sg13g2_nand2_1 _0755_ (.Y(_0274_),
    .A(_0268_),
    .B(_0273_));
 sg13g2_xnor2_1 _0756_ (.Y(_0275_),
    .A(_0240_),
    .B(_0250_));
 sg13g2_nor2b_1 _0757_ (.A(net83),
    .B_N(_0249_),
    .Y(_0276_));
 sg13g2_a21oi_1 _0758_ (.A1(net83),
    .A2(_0275_),
    .Y(_0277_),
    .B1(_0276_));
 sg13g2_nand2_1 _0759_ (.Y(_0278_),
    .A(net80),
    .B(_0277_));
 sg13g2_nand3_1 _0760_ (.B(net80),
    .C(_0277_),
    .A(_0007_),
    .Y(_0279_));
 sg13g2_xnor2_1 _0761_ (.Y(_0280_),
    .A(_0220_),
    .B(_0236_));
 sg13g2_nand2_1 _0762_ (.Y(_0281_),
    .A(net83),
    .B(_0280_));
 sg13g2_o21ai_1 _0763_ (.B1(_0281_),
    .Y(_0282_),
    .A1(_0217_),
    .A2(net83));
 sg13g2_nand2_1 _0764_ (.Y(_0283_),
    .A(net80),
    .B(_0282_));
 sg13g2_nand3_1 _0765_ (.B(net80),
    .C(_0282_),
    .A(_0008_),
    .Y(_0284_));
 sg13g2_and3_1 _0766_ (.X(_0285_),
    .A(_0268_),
    .B(_0273_),
    .C(_0279_));
 sg13g2_a22oi_1 _0767_ (.Y(_0286_),
    .B1(_0283_),
    .B2(_0086_),
    .A2(_0267_),
    .A1(\system_inst.loader.threshold[5] ));
 sg13g2_a22oi_1 _0768_ (.Y(_0287_),
    .B1(_0278_),
    .B2(_0085_),
    .A2(_0272_),
    .A1(\system_inst.loader.threshold[6] ));
 sg13g2_and4_1 _0769_ (.A(_0284_),
    .B(_0285_),
    .C(_0286_),
    .D(_0287_),
    .X(_0288_));
 sg13g2_xnor2_1 _0770_ (.Y(_0289_),
    .A(_0228_),
    .B(_0234_));
 sg13g2_nor2_1 _0771_ (.A(_0225_),
    .B(net84),
    .Y(_0290_));
 sg13g2_a21oi_1 _0772_ (.A1(net84),
    .A2(_0289_),
    .Y(_0291_),
    .B1(_0290_));
 sg13g2_inv_1 _0773_ (.Y(_0292_),
    .A(_0291_));
 sg13g2_o21ai_1 _0774_ (.B1(\system_inst.loader.threshold[2] ),
    .Y(_0293_),
    .A1(_0263_),
    .A2(_0292_));
 sg13g2_xor2_1 _0775_ (.B(_0235_),
    .A(_0223_),
    .X(_0294_));
 sg13g2_nand2_1 _0776_ (.Y(_0295_),
    .A(net84),
    .B(_0294_));
 sg13g2_o21ai_1 _0777_ (.B1(_0295_),
    .Y(_0296_),
    .A1(_0221_),
    .A2(net84));
 sg13g2_nand2_1 _0778_ (.Y(_0297_),
    .A(_0264_),
    .B(_0296_));
 sg13g2_a21o_1 _0779_ (.A2(_0296_),
    .A1(_0264_),
    .B1(_0006_),
    .X(_0298_));
 sg13g2_nand3_1 _0780_ (.B(net79),
    .C(_0291_),
    .A(_0077_),
    .Y(_0299_));
 sg13g2_and3_1 _0781_ (.X(_0300_),
    .A(_0006_),
    .B(net79),
    .C(_0296_));
 sg13g2_nand3_1 _0782_ (.B(net79),
    .C(_0296_),
    .A(_0006_),
    .Y(_0301_));
 sg13g2_nand4_1 _0783_ (.B(_0298_),
    .C(_0299_),
    .A(_0293_),
    .Y(_0302_),
    .D(_0301_));
 sg13g2_xnor2_1 _0784_ (.Y(_0303_),
    .A(_0232_),
    .B(_0233_));
 sg13g2_nor2b_1 _0785_ (.A(net84),
    .B_N(_0229_),
    .Y(_0304_));
 sg13g2_a21oi_2 _0786_ (.B1(_0304_),
    .Y(_0305_),
    .A2(_0303_),
    .A1(net84));
 sg13g2_nand2_1 _0787_ (.Y(_0306_),
    .A(net79),
    .B(_0305_));
 sg13g2_a21oi_1 _0788_ (.A1(net79),
    .A2(_0305_),
    .Y(_0307_),
    .B1(_0078_));
 sg13g2_nand3_1 _0789_ (.B(net79),
    .C(_0305_),
    .A(_0078_),
    .Y(_0308_));
 sg13g2_nand2_1 _0790_ (.Y(_0309_),
    .A(\system_inst.leak_rate[0] ),
    .B(net84));
 sg13g2_xor2_1 _0791_ (.B(_0309_),
    .A(_0231_),
    .X(_0310_));
 sg13g2_nand2_1 _0792_ (.Y(_0311_),
    .A(net79),
    .B(_0310_));
 sg13g2_nand3b_1 _0793_ (.B(net79),
    .C(_0310_),
    .Y(_0312_),
    .A_N(\system_inst.loader.threshold[0] ));
 sg13g2_nand2_1 _0794_ (.Y(_0313_),
    .A(_0308_),
    .B(_0312_));
 sg13g2_a21oi_1 _0795_ (.A1(_0308_),
    .A2(_0312_),
    .Y(_0314_),
    .B1(_0307_));
 sg13g2_a21o_1 _0796_ (.A2(_0298_),
    .A1(_0293_),
    .B1(_0300_),
    .X(_0315_));
 sg13g2_o21ai_1 _0797_ (.B1(_0315_),
    .Y(_0316_),
    .A1(_0302_),
    .A2(_0314_));
 sg13g2_o21ai_1 _0798_ (.B1(_0287_),
    .Y(_0317_),
    .A1(_0274_),
    .A2(_0286_));
 sg13g2_a22oi_1 _0799_ (.Y(_0318_),
    .B1(_0317_),
    .B2(_0279_),
    .A2(_0316_),
    .A1(_0288_));
 sg13g2_and2_1 _0800_ (.A(\system_inst.loader.threshold[0] ),
    .B(_0311_),
    .X(_0319_));
 sg13g2_nor4_1 _0801_ (.A(_0302_),
    .B(_0307_),
    .C(_0313_),
    .D(_0319_),
    .Y(_0320_));
 sg13g2_a21oi_2 _0802_ (.B1(_0318_),
    .Y(_0321_),
    .A2(_0320_),
    .A1(_0288_));
 sg13g2_nor2_1 _0803_ (.A(_0115_),
    .B(_0311_),
    .Y(_0322_));
 sg13g2_a22oi_1 _0804_ (.Y(_0323_),
    .B1(net78),
    .B2(_0322_),
    .A2(net86),
    .A1(net179));
 sg13g2_nor2_1 _0805_ (.A(net93),
    .B(_0323_),
    .Y(_0011_));
 sg13g2_nor2_1 _0806_ (.A(net86),
    .B(_0306_),
    .Y(_0324_));
 sg13g2_a22oi_1 _0807_ (.Y(_0325_),
    .B1(net78),
    .B2(_0324_),
    .A2(_0115_),
    .A1(net174));
 sg13g2_nor2_1 _0808_ (.A(net93),
    .B(_0325_),
    .Y(_0012_));
 sg13g2_nor3_1 _0809_ (.A(net86),
    .B(_0263_),
    .C(_0292_),
    .Y(_0326_));
 sg13g2_a22oi_1 _0810_ (.Y(_0327_),
    .B1(net78),
    .B2(_0326_),
    .A2(net86),
    .A1(net147));
 sg13g2_nor2_1 _0811_ (.A(net94),
    .B(_0327_),
    .Y(_0013_));
 sg13g2_nor2_1 _0812_ (.A(net86),
    .B(_0297_),
    .Y(_0328_));
 sg13g2_a22oi_1 _0813_ (.Y(_0329_),
    .B1(_0321_),
    .B2(_0328_),
    .A2(_0115_),
    .A1(net162));
 sg13g2_nor2_1 _0814_ (.A(net93),
    .B(_0329_),
    .Y(_0014_));
 sg13g2_nor2_1 _0815_ (.A(net85),
    .B(_0283_),
    .Y(_0330_));
 sg13g2_a22oi_1 _0816_ (.Y(_0331_),
    .B1(net78),
    .B2(_0330_),
    .A2(net86),
    .A1(net161));
 sg13g2_nor2_1 _0817_ (.A(net93),
    .B(_0331_),
    .Y(_0015_));
 sg13g2_nor2_1 _0818_ (.A(net85),
    .B(_0267_),
    .Y(_0332_));
 sg13g2_a22oi_1 _0819_ (.Y(_0333_),
    .B1(net78),
    .B2(_0332_),
    .A2(net86),
    .A1(net165));
 sg13g2_nor2_1 _0820_ (.A(net93),
    .B(_0333_),
    .Y(_0016_));
 sg13g2_nor2_1 _0821_ (.A(net85),
    .B(_0272_),
    .Y(_0334_));
 sg13g2_a22oi_1 _0822_ (.Y(_0335_),
    .B1(net78),
    .B2(_0334_),
    .A2(net85),
    .A1(net160));
 sg13g2_nor2_1 _0823_ (.A(net93),
    .B(_0335_),
    .Y(_0017_));
 sg13g2_nor2_1 _0824_ (.A(net85),
    .B(_0278_),
    .Y(_0336_));
 sg13g2_a22oi_1 _0825_ (.Y(_0337_),
    .B1(net78),
    .B2(_0336_),
    .A2(net85),
    .A1(net159));
 sg13g2_nor2_1 _0826_ (.A(net93),
    .B(_0337_),
    .Y(_0018_));
 sg13g2_and3_1 _0827_ (.X(_0019_),
    .A(net92),
    .B(net98),
    .C(net85));
 sg13g2_or2_1 _0828_ (.X(_0338_),
    .B(_0112_),
    .A(_0111_));
 sg13g2_o21ai_1 _0829_ (.B1(_0338_),
    .Y(_0339_),
    .A1(_0114_),
    .A2(_0321_));
 sg13g2_o21ai_1 _0830_ (.B1(_0339_),
    .Y(_0340_),
    .A1(net191),
    .A2(_0111_));
 sg13g2_o21ai_1 _0831_ (.B1(net100),
    .Y(_0341_),
    .A1(net191),
    .A2(_0339_));
 sg13g2_nor2b_1 _0832_ (.A(_0341_),
    .B_N(_0340_),
    .Y(_0020_));
 sg13g2_xnor2_1 _0833_ (.Y(_0342_),
    .A(net195),
    .B(\system_inst.neuron.refr_cnt[0] ));
 sg13g2_nand2b_1 _0834_ (.Y(_0343_),
    .B(_0342_),
    .A_N(_0338_));
 sg13g2_o21ai_1 _0835_ (.B1(_0343_),
    .Y(_0344_),
    .A1(_0084_),
    .A2(_0339_));
 sg13g2_and2_1 _0836_ (.A(net100),
    .B(net196),
    .X(_0021_));
 sg13g2_nand3_1 _0837_ (.B(_0110_),
    .C(_0339_),
    .A(_0083_),
    .Y(_0345_));
 sg13g2_a21o_1 _0838_ (.A2(_0339_),
    .A1(net198),
    .B1(_0083_),
    .X(_0346_));
 sg13g2_a21oi_1 _0839_ (.A1(net190),
    .A2(_0346_),
    .Y(_0022_),
    .B1(_0087_));
 sg13g2_and3_1 _0840_ (.X(_0023_),
    .A(net112),
    .B(net100),
    .C(_0345_));
 sg13g2_a21o_1 _0841_ (.A2(net84),
    .A1(_0113_),
    .B1(net95),
    .X(_0347_));
 sg13g2_xnor2_1 _0842_ (.Y(_0348_),
    .A(_0082_),
    .B(_0112_));
 sg13g2_nor2_1 _0843_ (.A(_0347_),
    .B(_0348_),
    .Y(_0024_));
 sg13g2_nor3_2 _0844_ (.A(_0081_),
    .B(_0082_),
    .C(_0112_),
    .Y(_0349_));
 sg13g2_a21oi_1 _0845_ (.A1(\system_inst.neuron.leak_counter[0] ),
    .A2(_0113_),
    .Y(_0350_),
    .B1(net118));
 sg13g2_nor3_1 _0846_ (.A(_0347_),
    .B(_0349_),
    .C(net119),
    .Y(_0025_));
 sg13g2_nand2_1 _0847_ (.Y(_0351_),
    .A(\system_inst.neuron.leak_counter[2] ),
    .B(_0349_));
 sg13g2_xnor2_1 _0848_ (.Y(_0352_),
    .A(net175),
    .B(_0349_));
 sg13g2_nor2_1 _0849_ (.A(_0347_),
    .B(net176),
    .Y(_0026_));
 sg13g2_xor2_1 _0850_ (.B(_0351_),
    .A(net172),
    .X(_0353_));
 sg13g2_nor2_1 _0851_ (.A(_0347_),
    .B(net173),
    .Y(_0027_));
 sg13g2_nor4_2 _0852_ (.A(\system_inst.loader.current_state[1] ),
    .B(\system_inst.loader.current_state[6] ),
    .C(\system_inst.loader.current_state[2] ),
    .Y(_0354_),
    .D(net116));
 sg13g2_nand2_1 _0853_ (.Y(_0355_),
    .A(net149),
    .B(_0354_));
 sg13g2_nor2_1 _0854_ (.A(net123),
    .B(_0355_),
    .Y(_0356_));
 sg13g2_o21ai_1 _0855_ (.B1(net1),
    .Y(_0357_),
    .A1(net3),
    .A2(_0089_));
 sg13g2_nor2_2 _0856_ (.A(_0356_),
    .B(_0357_),
    .Y(_0358_));
 sg13g2_and2_1 _0857_ (.A(_0088_),
    .B(_0354_),
    .X(_0359_));
 sg13g2_nand2_1 _0858_ (.Y(_0360_),
    .A(_0088_),
    .B(_0354_));
 sg13g2_o21ai_1 _0859_ (.B1(_0354_),
    .Y(_0361_),
    .A1(_0088_),
    .A2(net91));
 sg13g2_nand2_1 _0860_ (.Y(_0362_),
    .A(net3),
    .B(_0361_));
 sg13g2_nand2_1 _0861_ (.Y(_0363_),
    .A(_0358_),
    .B(_0362_));
 sg13g2_a21oi_1 _0862_ (.A1(net170),
    .A2(_0363_),
    .Y(_0364_),
    .B1(net95));
 sg13g2_o21ai_1 _0863_ (.B1(_0364_),
    .Y(_0028_),
    .A1(_0359_),
    .A2(_0363_));
 sg13g2_o21ai_1 _0864_ (.B1(net101),
    .Y(_0365_),
    .A1(net184),
    .A2(_0104_));
 sg13g2_a21oi_1 _0865_ (.A1(_0076_),
    .A2(_0104_),
    .Y(_0029_),
    .B1(_0365_));
 sg13g2_a21oi_1 _0866_ (.A1(net180),
    .A2(_0103_),
    .Y(_0366_),
    .B1(net95));
 sg13g2_o21ai_1 _0867_ (.B1(_0366_),
    .Y(_0030_),
    .A1(_0073_),
    .A2(_0103_));
 sg13g2_o21ai_1 _0868_ (.B1(net101),
    .Y(_0367_),
    .A1(net187),
    .A2(_0104_));
 sg13g2_a21oi_1 _0869_ (.A1(_0072_),
    .A2(_0104_),
    .Y(_0031_),
    .B1(_0367_));
 sg13g2_o21ai_1 _0870_ (.B1(net102),
    .Y(_0368_),
    .A1(net188),
    .A2(_0100_));
 sg13g2_a21oi_1 _0871_ (.A1(_0076_),
    .A2(_0100_),
    .Y(_0032_),
    .B1(_0368_));
 sg13g2_a21oi_1 _0872_ (.A1(net182),
    .A2(_0099_),
    .Y(_0369_),
    .B1(net95));
 sg13g2_o21ai_1 _0873_ (.B1(_0369_),
    .Y(_0033_),
    .A1(_0073_),
    .A2(_0099_));
 sg13g2_o21ai_1 _0874_ (.B1(net101),
    .Y(_0370_),
    .A1(net185),
    .A2(_0100_));
 sg13g2_a21oi_1 _0875_ (.A1(_0072_),
    .A2(_0100_),
    .Y(_0034_),
    .B1(_0370_));
 sg13g2_o21ai_1 _0876_ (.B1(net102),
    .Y(_0371_),
    .A1(net167),
    .A2(net89));
 sg13g2_a21oi_1 _0877_ (.A1(_0076_),
    .A2(net89),
    .Y(_0035_),
    .B1(_0371_));
 sg13g2_a21oi_1 _0878_ (.A1(\system_inst.loader.shift_reg[0] ),
    .A2(net89),
    .Y(_0372_),
    .B1(net95));
 sg13g2_o21ai_1 _0879_ (.B1(_0372_),
    .Y(_0036_),
    .A1(_0080_),
    .A2(net89));
 sg13g2_o21ai_1 _0880_ (.B1(net99),
    .Y(_0373_),
    .A1(net152),
    .A2(net89));
 sg13g2_a21oi_1 _0881_ (.A1(_0072_),
    .A2(net89),
    .Y(_0037_),
    .B1(_0373_));
 sg13g2_o21ai_1 _0882_ (.B1(net97),
    .Y(_0374_),
    .A1(net177),
    .A2(net89));
 sg13g2_a21oi_1 _0883_ (.A1(_0071_),
    .A2(net89),
    .Y(_0038_),
    .B1(_0374_));
 sg13g2_o21ai_1 _0884_ (.B1(net97),
    .Y(_0375_),
    .A1(net146),
    .A2(net90));
 sg13g2_a21oi_1 _0885_ (.A1(_0070_),
    .A2(net90),
    .Y(_0039_),
    .B1(_0375_));
 sg13g2_o21ai_1 _0886_ (.B1(net96),
    .Y(_0376_),
    .A1(\system_inst.leak_rate[5] ),
    .A2(net90));
 sg13g2_a21oi_1 _0887_ (.A1(_0069_),
    .A2(net90),
    .Y(_0040_),
    .B1(_0376_));
 sg13g2_o21ai_1 _0888_ (.B1(net96),
    .Y(_0377_),
    .A1(net154),
    .A2(net90));
 sg13g2_a21oi_1 _0889_ (.A1(_0068_),
    .A2(net90),
    .Y(_0041_),
    .B1(_0377_));
 sg13g2_o21ai_1 _0890_ (.B1(net98),
    .Y(_0378_),
    .A1(\system_inst.leak_rate[7] ),
    .A2(net90));
 sg13g2_a21oi_1 _0891_ (.A1(_0067_),
    .A2(net90),
    .Y(_0042_),
    .B1(_0378_));
 sg13g2_o21ai_1 _0892_ (.B1(net99),
    .Y(_0379_),
    .A1(net178),
    .A2(net88));
 sg13g2_a21oi_1 _0893_ (.A1(_0076_),
    .A2(net88),
    .Y(_0043_),
    .B1(_0379_));
 sg13g2_a21oi_1 _0894_ (.A1(\system_inst.loader.shift_reg[0] ),
    .A2(net88),
    .Y(_0380_),
    .B1(net94));
 sg13g2_o21ai_1 _0895_ (.B1(_0380_),
    .Y(_0044_),
    .A1(_0078_),
    .A2(net88));
 sg13g2_a21oi_1 _0896_ (.A1(\system_inst.loader.shift_reg[1] ),
    .A2(net87),
    .Y(_0381_),
    .B1(net94));
 sg13g2_o21ai_1 _0897_ (.B1(_0381_),
    .Y(_0045_),
    .A1(_0077_),
    .A2(net87));
 sg13g2_a21oi_1 _0898_ (.A1(net135),
    .A2(_0108_),
    .Y(_0382_),
    .B1(net94));
 sg13g2_o21ai_1 _0899_ (.B1(_0382_),
    .Y(_0046_),
    .A1(_0071_),
    .A2(_0108_));
 sg13g2_a21oi_1 _0900_ (.A1(net131),
    .A2(_0108_),
    .Y(_0383_),
    .B1(net94));
 sg13g2_o21ai_1 _0901_ (.B1(_0383_),
    .Y(_0047_),
    .A1(_0070_),
    .A2(_0108_));
 sg13g2_o21ai_1 _0902_ (.B1(net96),
    .Y(_0384_),
    .A1(net130),
    .A2(net87));
 sg13g2_a21oi_1 _0903_ (.A1(_0069_),
    .A2(net87),
    .Y(_0048_),
    .B1(_0384_));
 sg13g2_o21ai_1 _0904_ (.B1(net96),
    .Y(_0385_),
    .A1(net157),
    .A2(net87));
 sg13g2_a21oi_1 _0905_ (.A1(_0068_),
    .A2(net87),
    .Y(_0049_),
    .B1(_0385_));
 sg13g2_o21ai_1 _0906_ (.B1(net98),
    .Y(_0386_),
    .A1(net129),
    .A2(net87));
 sg13g2_a21oi_1 _0907_ (.A1(_0067_),
    .A2(net87),
    .Y(_0050_),
    .B1(_0386_));
 sg13g2_and3_2 _0908_ (.X(_0387_),
    .A(net124),
    .B(net91),
    .C(_0094_));
 sg13g2_o21ai_1 _0909_ (.B1(net99),
    .Y(_0388_),
    .A1(net158),
    .A2(_0387_));
 sg13g2_a21oi_1 _0910_ (.A1(_0076_),
    .A2(_0387_),
    .Y(_0051_),
    .B1(_0388_));
 sg13g2_a21oi_1 _0911_ (.A1(\system_inst.loader.shift_reg[0] ),
    .A2(_0387_),
    .Y(_0389_),
    .B1(net95));
 sg13g2_o21ai_1 _0912_ (.B1(_0389_),
    .Y(_0052_),
    .A1(_0075_),
    .A2(_0387_));
 sg13g2_o21ai_1 _0913_ (.B1(net99),
    .Y(_0390_),
    .A1(net155),
    .A2(_0387_));
 sg13g2_a21oi_1 _0914_ (.A1(_0072_),
    .A2(_0387_),
    .Y(_0053_),
    .B1(_0390_));
 sg13g2_o21ai_1 _0915_ (.B1(net99),
    .Y(_0391_),
    .A1(net166),
    .A2(_0387_));
 sg13g2_a21oi_1 _0916_ (.A1(_0071_),
    .A2(_0387_),
    .Y(_0054_),
    .B1(_0391_));
 sg13g2_nand2b_1 _0917_ (.Y(_0392_),
    .B(_0360_),
    .A_N(net3));
 sg13g2_and2_1 _0918_ (.A(_0358_),
    .B(_0392_),
    .X(_0393_));
 sg13g2_nand2_1 _0919_ (.Y(_0394_),
    .A(_0358_),
    .B(_0392_));
 sg13g2_a21oi_2 _0920_ (.B1(_0359_),
    .Y(_0395_),
    .A2(net91),
    .A1(_0088_));
 sg13g2_a21oi_1 _0921_ (.A1(net4),
    .A2(_0395_),
    .Y(_0396_),
    .B1(_0394_));
 sg13g2_o21ai_1 _0922_ (.B1(net99),
    .Y(_0397_),
    .A1(net186),
    .A2(_0393_));
 sg13g2_nor2_1 _0923_ (.A(_0396_),
    .B(_0397_),
    .Y(_0055_));
 sg13g2_a21oi_1 _0924_ (.A1(net186),
    .A2(_0395_),
    .Y(_0398_),
    .B1(net81));
 sg13g2_o21ai_1 _0925_ (.B1(net97),
    .Y(_0399_),
    .A1(net168),
    .A2(net82));
 sg13g2_nor2_1 _0926_ (.A(_0398_),
    .B(_0399_),
    .Y(_0056_));
 sg13g2_a21oi_1 _0927_ (.A1(net168),
    .A2(_0395_),
    .Y(_0400_),
    .B1(net81));
 sg13g2_o21ai_1 _0928_ (.B1(net97),
    .Y(_0401_),
    .A1(net133),
    .A2(net82));
 sg13g2_nor2_1 _0929_ (.A(_0400_),
    .B(_0401_),
    .Y(_0057_));
 sg13g2_a21oi_1 _0930_ (.A1(net133),
    .A2(_0395_),
    .Y(_0402_),
    .B1(net81));
 sg13g2_o21ai_1 _0931_ (.B1(net96),
    .Y(_0403_),
    .A1(\system_inst.loader.shift_reg[3] ),
    .A2(net82));
 sg13g2_nor2_1 _0932_ (.A(_0402_),
    .B(_0403_),
    .Y(_0058_));
 sg13g2_a21oi_1 _0933_ (.A1(net137),
    .A2(_0395_),
    .Y(_0404_),
    .B1(net81));
 sg13g2_o21ai_1 _0934_ (.B1(net96),
    .Y(_0405_),
    .A1(net125),
    .A2(net82));
 sg13g2_nor2_1 _0935_ (.A(_0404_),
    .B(_0405_),
    .Y(_0059_));
 sg13g2_a21oi_1 _0936_ (.A1(net125),
    .A2(_0395_),
    .Y(_0406_),
    .B1(net81));
 sg13g2_o21ai_1 _0937_ (.B1(net96),
    .Y(_0407_),
    .A1(net148),
    .A2(net82));
 sg13g2_nor2_1 _0938_ (.A(_0406_),
    .B(_0407_),
    .Y(_0060_));
 sg13g2_a21oi_1 _0939_ (.A1(net148),
    .A2(_0395_),
    .Y(_0408_),
    .B1(net81));
 sg13g2_o21ai_1 _0940_ (.B1(net96),
    .Y(_0409_),
    .A1(net127),
    .A2(net82));
 sg13g2_nor2_1 _0941_ (.A(_0408_),
    .B(_0409_),
    .Y(_0061_));
 sg13g2_nand3_1 _0942_ (.B(_0358_),
    .C(_0360_),
    .A(net3),
    .Y(_0410_));
 sg13g2_o21ai_1 _0943_ (.B1(net100),
    .Y(_0411_),
    .A1(_0066_),
    .A2(net81));
 sg13g2_a21oi_1 _0944_ (.A1(_0066_),
    .A2(_0410_),
    .Y(_0062_),
    .B1(_0411_));
 sg13g2_a21oi_1 _0945_ (.A1(net138),
    .A2(net82),
    .Y(_0412_),
    .B1(net169));
 sg13g2_nand3_1 _0946_ (.B(_0355_),
    .C(_0360_),
    .A(_0091_),
    .Y(_0413_));
 sg13g2_nand2b_1 _0947_ (.Y(_0414_),
    .B(net100),
    .A_N(_0412_));
 sg13g2_a21oi_1 _0948_ (.A1(net82),
    .A2(_0413_),
    .Y(_0063_),
    .B1(_0414_));
 sg13g2_a221oi_1 _0949_ (.B2(_0010_),
    .C1(_0410_),
    .B1(_0354_),
    .A1(_0009_),
    .Y(_0415_),
    .A2(_0091_));
 sg13g2_a22oi_1 _0950_ (.Y(_0416_),
    .B1(_0415_),
    .B2(_0093_),
    .A2(net81),
    .A1(net114));
 sg13g2_nor2_1 _0951_ (.A(net95),
    .B(net115),
    .Y(_0064_));
 sg13g2_nor3_1 _0952_ (.A(net93),
    .B(net85),
    .C(net78),
    .Y(_0065_));
 sg13g2_dfrbp_1 _0953_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net105),
    .D(_0011_),
    .Q_N(_0467_),
    .Q(\system_inst.neuron.v_mem[0] ));
 sg13g2_dfrbp_1 _0954_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net55),
    .D(_0012_),
    .Q_N(_0466_),
    .Q(\system_inst.neuron.v_mem[1] ));
 sg13g2_dfrbp_1 _0955_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net53),
    .D(_0013_),
    .Q_N(_0465_),
    .Q(\system_inst.neuron.v_mem[2] ));
 sg13g2_dfrbp_1 _0956_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net51),
    .D(_0014_),
    .Q_N(_0464_),
    .Q(\system_inst.neuron.v_mem[3] ));
 sg13g2_dfrbp_1 _0957_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net49),
    .D(_0015_),
    .Q_N(_0463_),
    .Q(\system_inst.neuron.v_mem[4] ));
 sg13g2_dfrbp_1 _0958_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net47),
    .D(_0016_),
    .Q_N(_0462_),
    .Q(\system_inst.neuron.v_mem[5] ));
 sg13g2_dfrbp_1 _0959_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net45),
    .D(_0017_),
    .Q_N(_0461_),
    .Q(\system_inst.neuron.v_mem[6] ));
 sg13g2_dfrbp_1 _0960_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net43),
    .D(_0018_),
    .Q_N(_0460_),
    .Q(\system_inst.neuron.v_mem[7] ));
 sg13g2_dfrbp_1 _0961_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net41),
    .D(_0019_),
    .Q_N(_0459_),
    .Q(\system_inst.neuron.v_mem[8] ));
 sg13g2_dfrbp_1 _0962_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net39),
    .D(net192),
    .Q_N(_0458_),
    .Q(\system_inst.neuron.refr_cnt[0] ));
 sg13g2_dfrbp_1 _0963_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net37),
    .D(_0021_),
    .Q_N(_0457_),
    .Q(\system_inst.neuron.refr_cnt[1] ));
 sg13g2_dfrbp_1 _0964_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net35),
    .D(_0022_),
    .Q_N(_0456_),
    .Q(\system_inst.neuron.refr_cnt[2] ));
 sg13g2_dfrbp_1 _0965_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net33),
    .D(net113),
    .Q_N(_0455_),
    .Q(\system_inst.neuron.refr_cnt[3] ));
 sg13g2_dfrbp_1 _0966_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net31),
    .D(_0024_),
    .Q_N(_0454_),
    .Q(\system_inst.neuron.leak_counter[0] ));
 sg13g2_dfrbp_1 _0967_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net29),
    .D(net120),
    .Q_N(_0453_),
    .Q(\system_inst.neuron.leak_counter[1] ));
 sg13g2_dfrbp_1 _0968_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net27),
    .D(_0026_),
    .Q_N(_0452_),
    .Q(\system_inst.neuron.leak_counter[2] ));
 sg13g2_dfrbp_1 _0969_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net25),
    .D(_0027_),
    .Q_N(_0451_),
    .Q(\system_inst.neuron.leak_counter[3] ));
 sg13g2_dfrbp_1 _0970_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net103),
    .D(net171),
    .Q_N(_0450_),
    .Q(params_ready));
 sg13g2_dfrbp_1 _0971_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net76),
    .D(_0029_),
    .Q_N(_0449_),
    .Q(\system_inst.loader.weight_a[0] ));
 sg13g2_dfrbp_1 _0972_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net74),
    .D(net181),
    .Q_N(_0448_),
    .Q(\system_inst.loader.weight_a[1] ));
 sg13g2_dfrbp_1 _0973_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net72),
    .D(_0031_),
    .Q_N(_0447_),
    .Q(\system_inst.loader.weight_a[2] ));
 sg13g2_dfrbp_1 _0974_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net70),
    .D(_0032_),
    .Q_N(_0446_),
    .Q(\system_inst.loader.weight_b[0] ));
 sg13g2_dfrbp_1 _0975_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net68),
    .D(net183),
    .Q_N(_0445_),
    .Q(\system_inst.loader.weight_b[1] ));
 sg13g2_dfrbp_1 _0976_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net66),
    .D(_0034_),
    .Q_N(_0444_),
    .Q(\system_inst.loader.weight_b[2] ));
 sg13g2_dfrbp_1 _0977_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net64),
    .D(_0035_),
    .Q_N(_0443_),
    .Q(\system_inst.leak_rate[0] ));
 sg13g2_dfrbp_1 _0978_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net62),
    .D(net151),
    .Q_N(_0442_),
    .Q(\system_inst.leak_rate[1] ));
 sg13g2_dfrbp_1 _0979_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net60),
    .D(net153),
    .Q_N(_0441_),
    .Q(\system_inst.leak_rate[2] ));
 sg13g2_dfrbp_1 _0980_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net58),
    .D(_0038_),
    .Q_N(_0440_),
    .Q(\system_inst.leak_rate[3] ));
 sg13g2_dfrbp_1 _0981_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net56),
    .D(_0039_),
    .Q_N(_0439_),
    .Q(\system_inst.leak_rate[4] ));
 sg13g2_dfrbp_1 _0982_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net52),
    .D(net126),
    .Q_N(_0438_),
    .Q(\system_inst.leak_rate[5] ));
 sg13g2_dfrbp_1 _0983_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net48),
    .D(_0041_),
    .Q_N(_0437_),
    .Q(\system_inst.leak_rate[6] ));
 sg13g2_dfrbp_1 _0984_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net44),
    .D(net128),
    .Q_N(_0436_),
    .Q(\system_inst.leak_rate[7] ));
 sg13g2_dfrbp_1 _0985_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net40),
    .D(_0043_),
    .Q_N(_0435_),
    .Q(\system_inst.loader.threshold[0] ));
 sg13g2_dfrbp_1 _0986_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net36),
    .D(net143),
    .Q_N(_0434_),
    .Q(\system_inst.loader.threshold[1] ));
 sg13g2_dfrbp_1 _0987_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net32),
    .D(net145),
    .Q_N(_0433_),
    .Q(\system_inst.loader.threshold[2] ));
 sg13g2_dfrbp_1 _0988_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net28),
    .D(net136),
    .Q_N(_0006_),
    .Q(\system_inst.loader.threshold[3] ));
 sg13g2_dfrbp_1 _0989_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net104),
    .D(net132),
    .Q_N(_0008_),
    .Q(\system_inst.loader.threshold[4] ));
 sg13g2_dfrbp_1 _0990_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net75),
    .D(_0048_),
    .Q_N(_0432_),
    .Q(\system_inst.loader.threshold[5] ));
 sg13g2_dfrbp_1 _0991_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net71),
    .D(_0049_),
    .Q_N(_0431_),
    .Q(\system_inst.loader.threshold[6] ));
 sg13g2_dfrbp_1 _0992_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net67),
    .D(_0050_),
    .Q_N(_0007_),
    .Q(\system_inst.loader.threshold[7] ));
 sg13g2_dfrbp_1 _0993_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net63),
    .D(_0051_),
    .Q_N(_0430_),
    .Q(\system_inst.leak_cycles[0] ));
 sg13g2_dfrbp_1 _0994_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net59),
    .D(net122),
    .Q_N(_0429_),
    .Q(\system_inst.leak_cycles[1] ));
 sg13g2_dfrbp_1 _0995_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net54),
    .D(net156),
    .Q_N(_0428_),
    .Q(\system_inst.leak_cycles[2] ));
 sg13g2_dfrbp_1 _0996_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net46),
    .D(_0054_),
    .Q_N(_0427_),
    .Q(\system_inst.leak_cycles[3] ));
 sg13g2_dfrbp_1 _0997_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net38),
    .D(_0055_),
    .Q_N(_0426_),
    .Q(\system_inst.loader.shift_reg[0] ));
 sg13g2_dfrbp_1 _0998_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net30),
    .D(_0056_),
    .Q_N(_0425_),
    .Q(\system_inst.loader.shift_reg[1] ));
 sg13g2_dfrbp_1 _0999_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net77),
    .D(_0057_),
    .Q_N(_0424_),
    .Q(\system_inst.loader.shift_reg[2] ));
 sg13g2_dfrbp_1 _1000_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net69),
    .D(net134),
    .Q_N(_0423_),
    .Q(\system_inst.loader.shift_reg[3] ));
 sg13g2_dfrbp_1 _1001_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net61),
    .D(_0059_),
    .Q_N(_0422_),
    .Q(\system_inst.loader.shift_reg[4] ));
 sg13g2_dfrbp_1 _1002_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net50),
    .D(_0060_),
    .Q_N(_0421_),
    .Q(\system_inst.loader.shift_reg[5] ));
 sg13g2_dfrbp_1 _1003_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net34),
    .D(_0061_),
    .Q_N(_0420_),
    .Q(\system_inst.loader.shift_reg[6] ));
 sg13g2_dfrbp_1 _1004_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net73),
    .D(_0062_),
    .Q_N(_0419_),
    .Q(\system_inst.loader.bit_count[0] ));
 sg13g2_dfrbp_1 _1005_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net57),
    .D(_0063_),
    .Q_N(_0418_),
    .Q(\system_inst.loader.bit_count[1] ));
 sg13g2_dfrbp_1 _1006_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net26),
    .D(_0064_),
    .Q_N(_0009_),
    .Q(\system_inst.loader.bit_count[2] ));
 sg13g2_dfrbp_1 _1007_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net106),
    .D(_0065_),
    .Q_N(_0468_),
    .Q(spike_out));
 sg13g2_dfrbp_1 _1008_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net107),
    .D(_0000_),
    .Q_N(_0469_),
    .Q(\system_inst.loader.current_state[0] ));
 sg13g2_dfrbp_1 _1009_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net108),
    .D(_0001_),
    .Q_N(_0470_),
    .Q(\system_inst.loader.current_state[1] ));
 sg13g2_dfrbp_1 _1010_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net109),
    .D(_0002_),
    .Q_N(_0471_),
    .Q(\system_inst.loader.current_state[2] ));
 sg13g2_dfrbp_1 _1011_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net110),
    .D(net117),
    .Q_N(_0472_),
    .Q(\system_inst.loader.current_state[4] ));
 sg13g2_dfrbp_1 _1012_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net65),
    .D(_0004_),
    .Q_N(_0010_),
    .Q(\system_inst.loader.current_state[5] ));
 sg13g2_dfrbp_1 _1013_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net42),
    .D(_0005_),
    .Q_N(_0417_),
    .Q(\system_inst.loader.current_state[6] ));
 sg13g2_tiehi _1006__26 (.L_HI(net26));
 sg13g2_tiehi _0968__27 (.L_HI(net27));
 sg13g2_tiehi _0988__28 (.L_HI(net28));
 sg13g2_tiehi _0967__29 (.L_HI(net29));
 sg13g2_tiehi _0998__30 (.L_HI(net30));
 sg13g2_tiehi _0966__31 (.L_HI(net31));
 sg13g2_tiehi _0987__32 (.L_HI(net32));
 sg13g2_tiehi _0965__33 (.L_HI(net33));
 sg13g2_tiehi _1003__34 (.L_HI(net34));
 sg13g2_tiehi _0964__35 (.L_HI(net35));
 sg13g2_tiehi _0986__36 (.L_HI(net36));
 sg13g2_tiehi _0963__37 (.L_HI(net37));
 sg13g2_tiehi _0997__38 (.L_HI(net38));
 sg13g2_tiehi _0962__39 (.L_HI(net39));
 sg13g2_tiehi _0985__40 (.L_HI(net40));
 sg13g2_tiehi _0961__41 (.L_HI(net41));
 sg13g2_tiehi _1013__42 (.L_HI(net42));
 sg13g2_tiehi _0960__43 (.L_HI(net43));
 sg13g2_tiehi _0984__44 (.L_HI(net44));
 sg13g2_tiehi _0959__45 (.L_HI(net45));
 sg13g2_tiehi _0996__46 (.L_HI(net46));
 sg13g2_tiehi _0958__47 (.L_HI(net47));
 sg13g2_tiehi _0983__48 (.L_HI(net48));
 sg13g2_tiehi _0957__49 (.L_HI(net49));
 sg13g2_tiehi _1002__50 (.L_HI(net50));
 sg13g2_tiehi _0956__51 (.L_HI(net51));
 sg13g2_tiehi _0982__52 (.L_HI(net52));
 sg13g2_tiehi _0955__53 (.L_HI(net53));
 sg13g2_tiehi _0995__54 (.L_HI(net54));
 sg13g2_tiehi _0954__55 (.L_HI(net55));
 sg13g2_tiehi _0981__56 (.L_HI(net56));
 sg13g2_tiehi _1005__57 (.L_HI(net57));
 sg13g2_tiehi _0980__58 (.L_HI(net58));
 sg13g2_tiehi _0994__59 (.L_HI(net59));
 sg13g2_tiehi _0979__60 (.L_HI(net60));
 sg13g2_tiehi _1001__61 (.L_HI(net61));
 sg13g2_tiehi _0978__62 (.L_HI(net62));
 sg13g2_tiehi _0993__63 (.L_HI(net63));
 sg13g2_tiehi _0977__64 (.L_HI(net64));
 sg13g2_tiehi _1012__65 (.L_HI(net65));
 sg13g2_tiehi _0976__66 (.L_HI(net66));
 sg13g2_tiehi _0992__67 (.L_HI(net67));
 sg13g2_tiehi _0975__68 (.L_HI(net68));
 sg13g2_tiehi _1000__69 (.L_HI(net69));
 sg13g2_tiehi _0974__70 (.L_HI(net70));
 sg13g2_tiehi _0991__71 (.L_HI(net71));
 sg13g2_tiehi _0973__72 (.L_HI(net72));
 sg13g2_tiehi _1004__73 (.L_HI(net73));
 sg13g2_tiehi _0972__74 (.L_HI(net74));
 sg13g2_tiehi _0990__75 (.L_HI(net75));
 sg13g2_tiehi _0971__76 (.L_HI(net76));
 sg13g2_tiehi _0999__77 (.L_HI(net77));
 sg13g2_tiehi _0970__78 (.L_HI(net103));
 sg13g2_tiehi _0989__79 (.L_HI(net104));
 sg13g2_tiehi _0953__80 (.L_HI(net105));
 sg13g2_tiehi _1007__81 (.L_HI(net106));
 sg13g2_tiehi _1008__82 (.L_HI(net107));
 sg13g2_tiehi _1009__83 (.L_HI(net108));
 sg13g2_tiehi _1010__84 (.L_HI(net109));
 sg13g2_tiehi _1011__85 (.L_HI(net110));
 sg13g2_tiehi tt_um_wokwi_434917577229968385_86 (.L_HI(net111));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_wokwi_434917577229968385_12 (.L_LO(net12));
 sg13g2_tielo tt_um_wokwi_434917577229968385_13 (.L_LO(net13));
 sg13g2_tielo tt_um_wokwi_434917577229968385_14 (.L_LO(net14));
 sg13g2_tielo tt_um_wokwi_434917577229968385_15 (.L_LO(net15));
 sg13g2_tielo tt_um_wokwi_434917577229968385_16 (.L_LO(net16));
 sg13g2_tielo tt_um_wokwi_434917577229968385_17 (.L_LO(net17));
 sg13g2_tielo tt_um_wokwi_434917577229968385_18 (.L_LO(net18));
 sg13g2_tielo tt_um_wokwi_434917577229968385_19 (.L_LO(net19));
 sg13g2_tielo tt_um_wokwi_434917577229968385_20 (.L_LO(net20));
 sg13g2_tielo tt_um_wokwi_434917577229968385_21 (.L_LO(net21));
 sg13g2_tielo tt_um_wokwi_434917577229968385_22 (.L_LO(net22));
 sg13g2_tielo tt_um_wokwi_434917577229968385_23 (.L_LO(net23));
 sg13g2_tielo tt_um_wokwi_434917577229968385_24 (.L_LO(net24));
 sg13g2_tiehi _0969__25 (.L_HI(net25));
 sg13g2_buf_2 _1090_ (.A(params_ready),
    .X(uio_out[0]));
 sg13g2_buf_1 _1091_ (.A(spike_out),
    .X(uo_out[0]));
 sg13g2_buf_4 fanout78 (.X(net78),
    .A(_0321_));
 sg13g2_buf_2 fanout79 (.A(net80),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_0264_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_0394_),
    .X(net81));
 sg13g2_buf_4 fanout82 (.X(net82),
    .A(_0393_));
 sg13g2_buf_2 fanout83 (.A(_0256_),
    .X(net83));
 sg13g2_buf_4 fanout84 (.X(net84),
    .A(_0256_));
 sg13g2_buf_2 fanout85 (.A(net86),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_0115_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_0107_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_0107_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_0097_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_0097_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_0092_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(net194),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(net94),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(net95),
    .X(net94));
 sg13g2_buf_4 fanout95 (.X(net95),
    .A(_0087_));
 sg13g2_buf_2 fanout96 (.A(net97),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(net98),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(rst_n),
    .X(net98));
 sg13g2_buf_4 fanout99 (.X(net99),
    .A(net102));
 sg13g2_buf_2 fanout100 (.A(net102),
    .X(net100));
 sg13g2_buf_4 fanout101 (.X(net101),
    .A(net102));
 sg13g2_buf_2 fanout102 (.A(rst_n),
    .X(net102));
 sg13g2_buf_2 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_buf_2 input10 (.A(uio_in[0]),
    .X(net10));
 sg13g2_tielo tt_um_wokwi_434917577229968385_11 (.L_LO(net11));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\system_inst.neuron.refr_cnt[3] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0023_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold3 (.A(\system_inst.loader.bit_count[2] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0416_),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold5 (.A(\system_inst.loader.current_state[4] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0003_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold7 (.A(\system_inst.neuron.leak_counter[1] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0350_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0025_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold10 (.A(\system_inst.leak_cycles[1] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0052_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold12 (.A(\system_inst.loader.current_state[0] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold13 (.A(\system_inst.loader.current_state[5] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold14 (.A(\system_inst.loader.shift_reg[4] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0040_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold16 (.A(\system_inst.loader.shift_reg[6] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0042_),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold18 (.A(\system_inst.loader.threshold[7] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold19 (.A(\system_inst.loader.threshold[5] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold20 (.A(\system_inst.loader.threshold[4] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0047_),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold22 (.A(\system_inst.loader.shift_reg[2] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0058_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold24 (.A(\system_inst.loader.threshold[3] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0046_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold26 (.A(\system_inst.loader.shift_reg[3] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold27 (.A(\system_inst.loader.bit_count[0] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold28 (.A(\system_inst.loader.current_state[6] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0101_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold30 (.A(\system_inst.loader.current_state[2] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold31 (.A(\system_inst.loader.threshold[1] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0044_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold33 (.A(\system_inst.loader.threshold[2] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0045_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold35 (.A(\system_inst.leak_rate[4] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold36 (.A(\system_inst.neuron.v_mem[2] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold37 (.A(\system_inst.loader.shift_reg[5] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0010_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold39 (.A(\system_inst.leak_rate[1] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0036_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold41 (.A(\system_inst.leak_rate[2] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0037_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold43 (.A(\system_inst.leak_rate[6] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold44 (.A(\system_inst.leak_cycles[2] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0053_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold46 (.A(\system_inst.loader.threshold[6] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold47 (.A(\system_inst.leak_cycles[0] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold48 (.A(\system_inst.neuron.v_mem[7] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold49 (.A(\system_inst.neuron.v_mem[6] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold50 (.A(\system_inst.neuron.v_mem[4] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold51 (.A(\system_inst.neuron.v_mem[3] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold52 (.A(\system_inst.loader.current_state[1] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0098_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold54 (.A(\system_inst.neuron.v_mem[5] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold55 (.A(\system_inst.leak_cycles[3] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold56 (.A(\system_inst.leak_rate[0] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold57 (.A(\system_inst.loader.shift_reg[1] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold58 (.A(\system_inst.loader.bit_count[1] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold59 (.A(params_ready),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0028_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold61 (.A(\system_inst.neuron.leak_counter[3] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0353_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold63 (.A(\system_inst.neuron.v_mem[1] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold64 (.A(\system_inst.neuron.leak_counter[2] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0352_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold66 (.A(\system_inst.leak_rate[3] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold67 (.A(\system_inst.loader.threshold[0] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold68 (.A(\system_inst.neuron.v_mem[0] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold69 (.A(\system_inst.loader.weight_a[1] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0030_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold71 (.A(\system_inst.loader.weight_b[1] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0033_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold73 (.A(\system_inst.loader.weight_a[0] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold74 (.A(\system_inst.loader.weight_b[2] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold75 (.A(\system_inst.loader.shift_reg[0] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold76 (.A(\system_inst.loader.weight_a[2] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold77 (.A(\system_inst.loader.weight_b[0] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold78 (.A(\system_inst.neuron.refr_cnt[2] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0345_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold80 (.A(\system_inst.neuron.refr_cnt[0] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0020_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold82 (.A(\system_inst.neuron.leak_counter[0] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold83 (.A(\system_inst.neuron.v_mem[8] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold84 (.A(\system_inst.neuron.refr_cnt[1] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0344_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold86 (.A(\system_inst.neuron.refr_cnt[1] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0110_),
    .X(net198));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_4 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_295 ();
 sg13g2_decap_8 FILLER_14_302 ();
 sg13g2_decap_8 FILLER_14_309 ();
 sg13g2_decap_8 FILLER_14_316 ();
 sg13g2_decap_8 FILLER_14_323 ();
 sg13g2_decap_8 FILLER_14_330 ();
 sg13g2_decap_8 FILLER_14_337 ();
 sg13g2_decap_8 FILLER_14_344 ();
 sg13g2_decap_8 FILLER_14_351 ();
 sg13g2_decap_8 FILLER_14_358 ();
 sg13g2_decap_8 FILLER_14_365 ();
 sg13g2_decap_8 FILLER_14_372 ();
 sg13g2_decap_8 FILLER_14_379 ();
 sg13g2_decap_8 FILLER_14_386 ();
 sg13g2_decap_8 FILLER_14_393 ();
 sg13g2_decap_8 FILLER_14_400 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_4 FILLER_15_196 ();
 sg13g2_fill_2 FILLER_15_200 ();
 sg13g2_decap_8 FILLER_15_206 ();
 sg13g2_fill_1 FILLER_15_213 ();
 sg13g2_decap_4 FILLER_15_240 ();
 sg13g2_fill_2 FILLER_15_244 ();
 sg13g2_fill_1 FILLER_15_272 ();
 sg13g2_decap_8 FILLER_15_306 ();
 sg13g2_decap_8 FILLER_15_313 ();
 sg13g2_decap_8 FILLER_15_320 ();
 sg13g2_decap_8 FILLER_15_327 ();
 sg13g2_decap_8 FILLER_15_334 ();
 sg13g2_decap_8 FILLER_15_341 ();
 sg13g2_decap_8 FILLER_15_348 ();
 sg13g2_decap_8 FILLER_15_355 ();
 sg13g2_decap_8 FILLER_15_362 ();
 sg13g2_decap_8 FILLER_15_369 ();
 sg13g2_decap_8 FILLER_15_376 ();
 sg13g2_decap_8 FILLER_15_383 ();
 sg13g2_decap_8 FILLER_15_390 ();
 sg13g2_decap_8 FILLER_15_397 ();
 sg13g2_decap_4 FILLER_15_404 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_4 FILLER_16_154 ();
 sg13g2_fill_2 FILLER_16_158 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_fill_2 FILLER_16_189 ();
 sg13g2_fill_2 FILLER_16_238 ();
 sg13g2_fill_1 FILLER_16_263 ();
 sg13g2_fill_2 FILLER_16_303 ();
 sg13g2_fill_1 FILLER_16_305 ();
 sg13g2_fill_1 FILLER_16_332 ();
 sg13g2_decap_8 FILLER_16_342 ();
 sg13g2_decap_8 FILLER_16_349 ();
 sg13g2_decap_8 FILLER_16_356 ();
 sg13g2_decap_8 FILLER_16_363 ();
 sg13g2_decap_8 FILLER_16_370 ();
 sg13g2_decap_8 FILLER_16_377 ();
 sg13g2_decap_8 FILLER_16_384 ();
 sg13g2_decap_8 FILLER_16_391 ();
 sg13g2_decap_8 FILLER_16_398 ();
 sg13g2_decap_4 FILLER_16_405 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_fill_1 FILLER_17_147 ();
 sg13g2_fill_1 FILLER_17_152 ();
 sg13g2_fill_1 FILLER_17_162 ();
 sg13g2_fill_1 FILLER_17_171 ();
 sg13g2_decap_4 FILLER_17_190 ();
 sg13g2_fill_1 FILLER_17_198 ();
 sg13g2_decap_8 FILLER_17_225 ();
 sg13g2_fill_2 FILLER_17_232 ();
 sg13g2_fill_1 FILLER_17_244 ();
 sg13g2_fill_1 FILLER_17_271 ();
 sg13g2_decap_8 FILLER_17_307 ();
 sg13g2_fill_2 FILLER_17_314 ();
 sg13g2_fill_1 FILLER_17_316 ();
 sg13g2_fill_1 FILLER_17_321 ();
 sg13g2_fill_1 FILLER_17_326 ();
 sg13g2_decap_8 FILLER_17_353 ();
 sg13g2_decap_8 FILLER_17_360 ();
 sg13g2_decap_8 FILLER_17_367 ();
 sg13g2_decap_8 FILLER_17_374 ();
 sg13g2_decap_8 FILLER_17_381 ();
 sg13g2_decap_8 FILLER_17_388 ();
 sg13g2_decap_8 FILLER_17_395 ();
 sg13g2_decap_8 FILLER_17_402 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_4 FILLER_18_133 ();
 sg13g2_fill_2 FILLER_18_172 ();
 sg13g2_decap_8 FILLER_18_200 ();
 sg13g2_fill_1 FILLER_18_207 ();
 sg13g2_fill_1 FILLER_18_225 ();
 sg13g2_decap_8 FILLER_18_253 ();
 sg13g2_fill_2 FILLER_18_260 ();
 sg13g2_fill_1 FILLER_18_262 ();
 sg13g2_fill_2 FILLER_18_279 ();
 sg13g2_fill_1 FILLER_18_307 ();
 sg13g2_fill_2 FILLER_18_336 ();
 sg13g2_decap_4 FILLER_18_356 ();
 sg13g2_fill_1 FILLER_18_360 ();
 sg13g2_decap_8 FILLER_18_374 ();
 sg13g2_decap_8 FILLER_18_381 ();
 sg13g2_decap_8 FILLER_18_388 ();
 sg13g2_decap_8 FILLER_18_395 ();
 sg13g2_decap_8 FILLER_18_402 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_4 FILLER_19_140 ();
 sg13g2_fill_2 FILLER_19_157 ();
 sg13g2_fill_1 FILLER_19_159 ();
 sg13g2_decap_8 FILLER_19_181 ();
 sg13g2_fill_1 FILLER_19_198 ();
 sg13g2_decap_8 FILLER_19_211 ();
 sg13g2_decap_8 FILLER_19_225 ();
 sg13g2_decap_4 FILLER_19_245 ();
 sg13g2_fill_2 FILLER_19_249 ();
 sg13g2_fill_2 FILLER_19_277 ();
 sg13g2_fill_1 FILLER_19_291 ();
 sg13g2_fill_1 FILLER_19_296 ();
 sg13g2_fill_1 FILLER_19_316 ();
 sg13g2_fill_2 FILLER_19_321 ();
 sg13g2_decap_4 FILLER_19_327 ();
 sg13g2_decap_8 FILLER_19_382 ();
 sg13g2_decap_8 FILLER_19_389 ();
 sg13g2_decap_8 FILLER_19_396 ();
 sg13g2_decap_4 FILLER_19_403 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_fill_1 FILLER_20_133 ();
 sg13g2_fill_1 FILLER_20_160 ();
 sg13g2_decap_4 FILLER_20_187 ();
 sg13g2_decap_4 FILLER_20_204 ();
 sg13g2_decap_8 FILLER_20_248 ();
 sg13g2_decap_8 FILLER_20_255 ();
 sg13g2_decap_4 FILLER_20_266 ();
 sg13g2_fill_2 FILLER_20_270 ();
 sg13g2_fill_2 FILLER_20_285 ();
 sg13g2_fill_2 FILLER_20_340 ();
 sg13g2_decap_8 FILLER_20_352 ();
 sg13g2_decap_4 FILLER_20_359 ();
 sg13g2_fill_2 FILLER_20_363 ();
 sg13g2_decap_8 FILLER_20_391 ();
 sg13g2_decap_8 FILLER_20_398 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_fill_2 FILLER_21_119 ();
 sg13g2_fill_1 FILLER_21_121 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_4 FILLER_21_133 ();
 sg13g2_fill_2 FILLER_21_137 ();
 sg13g2_decap_8 FILLER_21_144 ();
 sg13g2_decap_8 FILLER_21_151 ();
 sg13g2_fill_1 FILLER_21_158 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_fill_1 FILLER_21_180 ();
 sg13g2_fill_2 FILLER_21_195 ();
 sg13g2_fill_1 FILLER_21_197 ();
 sg13g2_fill_2 FILLER_21_220 ();
 sg13g2_fill_1 FILLER_21_267 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_fill_2 FILLER_21_301 ();
 sg13g2_fill_1 FILLER_21_303 ();
 sg13g2_decap_8 FILLER_21_307 ();
 sg13g2_decap_4 FILLER_21_314 ();
 sg13g2_fill_1 FILLER_21_332 ();
 sg13g2_fill_2 FILLER_21_342 ();
 sg13g2_fill_2 FILLER_21_365 ();
 sg13g2_decap_8 FILLER_21_388 ();
 sg13g2_decap_8 FILLER_21_395 ();
 sg13g2_decap_8 FILLER_21_402 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_4 FILLER_22_105 ();
 sg13g2_fill_2 FILLER_22_109 ();
 sg13g2_fill_2 FILLER_22_146 ();
 sg13g2_fill_1 FILLER_22_148 ();
 sg13g2_fill_1 FILLER_22_175 ();
 sg13g2_fill_2 FILLER_22_184 ();
 sg13g2_decap_8 FILLER_22_190 ();
 sg13g2_decap_4 FILLER_22_197 ();
 sg13g2_fill_2 FILLER_22_201 ();
 sg13g2_decap_8 FILLER_22_257 ();
 sg13g2_decap_8 FILLER_22_264 ();
 sg13g2_fill_2 FILLER_22_271 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_4 FILLER_22_294 ();
 sg13g2_decap_4 FILLER_22_306 ();
 sg13g2_fill_1 FILLER_22_310 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_fill_2 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_328 ();
 sg13g2_fill_2 FILLER_22_335 ();
 sg13g2_decap_8 FILLER_22_346 ();
 sg13g2_fill_2 FILLER_22_353 ();
 sg13g2_fill_1 FILLER_22_355 ();
 sg13g2_fill_1 FILLER_22_365 ();
 sg13g2_fill_2 FILLER_22_378 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_fill_2 FILLER_23_91 ();
 sg13g2_fill_2 FILLER_23_119 ();
 sg13g2_fill_1 FILLER_23_125 ();
 sg13g2_fill_1 FILLER_23_135 ();
 sg13g2_decap_8 FILLER_23_141 ();
 sg13g2_fill_2 FILLER_23_167 ();
 sg13g2_fill_1 FILLER_23_169 ();
 sg13g2_decap_4 FILLER_23_204 ();
 sg13g2_fill_1 FILLER_23_208 ();
 sg13g2_decap_4 FILLER_23_214 ();
 sg13g2_fill_2 FILLER_23_235 ();
 sg13g2_fill_1 FILLER_23_237 ();
 sg13g2_fill_2 FILLER_23_255 ();
 sg13g2_fill_1 FILLER_23_257 ();
 sg13g2_decap_4 FILLER_23_263 ();
 sg13g2_fill_2 FILLER_23_267 ();
 sg13g2_decap_4 FILLER_23_282 ();
 sg13g2_fill_1 FILLER_23_286 ();
 sg13g2_decap_4 FILLER_23_329 ();
 sg13g2_fill_2 FILLER_23_333 ();
 sg13g2_fill_2 FILLER_23_348 ();
 sg13g2_decap_4 FILLER_23_362 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_4 FILLER_24_98 ();
 sg13g2_fill_2 FILLER_24_102 ();
 sg13g2_decap_4 FILLER_24_108 ();
 sg13g2_fill_1 FILLER_24_112 ();
 sg13g2_fill_2 FILLER_24_122 ();
 sg13g2_fill_1 FILLER_24_124 ();
 sg13g2_decap_8 FILLER_24_143 ();
 sg13g2_decap_4 FILLER_24_150 ();
 sg13g2_fill_1 FILLER_24_154 ();
 sg13g2_decap_4 FILLER_24_172 ();
 sg13g2_fill_1 FILLER_24_176 ();
 sg13g2_fill_1 FILLER_24_180 ();
 sg13g2_fill_1 FILLER_24_194 ();
 sg13g2_fill_2 FILLER_24_200 ();
 sg13g2_fill_1 FILLER_24_202 ();
 sg13g2_fill_1 FILLER_24_208 ();
 sg13g2_fill_2 FILLER_24_214 ();
 sg13g2_fill_1 FILLER_24_216 ();
 sg13g2_fill_1 FILLER_24_253 ();
 sg13g2_decap_8 FILLER_24_285 ();
 sg13g2_decap_4 FILLER_24_292 ();
 sg13g2_fill_2 FILLER_24_296 ();
 sg13g2_fill_2 FILLER_24_305 ();
 sg13g2_decap_4 FILLER_24_332 ();
 sg13g2_fill_1 FILLER_24_336 ();
 sg13g2_decap_8 FILLER_24_341 ();
 sg13g2_decap_8 FILLER_24_348 ();
 sg13g2_fill_1 FILLER_24_367 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_4 FILLER_25_84 ();
 sg13g2_fill_1 FILLER_25_88 ();
 sg13g2_decap_4 FILLER_25_115 ();
 sg13g2_fill_2 FILLER_25_134 ();
 sg13g2_fill_1 FILLER_25_167 ();
 sg13g2_decap_4 FILLER_25_221 ();
 sg13g2_fill_2 FILLER_25_230 ();
 sg13g2_fill_2 FILLER_25_241 ();
 sg13g2_fill_1 FILLER_25_243 ();
 sg13g2_decap_4 FILLER_25_249 ();
 sg13g2_decap_8 FILLER_25_258 ();
 sg13g2_fill_2 FILLER_25_265 ();
 sg13g2_fill_1 FILLER_25_267 ();
 sg13g2_decap_8 FILLER_25_277 ();
 sg13g2_fill_2 FILLER_25_294 ();
 sg13g2_fill_1 FILLER_25_296 ();
 sg13g2_fill_2 FILLER_25_307 ();
 sg13g2_decap_4 FILLER_25_352 ();
 sg13g2_fill_2 FILLER_25_356 ();
 sg13g2_fill_1 FILLER_25_368 ();
 sg13g2_fill_1 FILLER_25_380 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_fill_2 FILLER_26_98 ();
 sg13g2_fill_1 FILLER_26_104 ();
 sg13g2_decap_8 FILLER_26_114 ();
 sg13g2_fill_1 FILLER_26_121 ();
 sg13g2_decap_8 FILLER_26_127 ();
 sg13g2_decap_8 FILLER_26_134 ();
 sg13g2_fill_1 FILLER_26_150 ();
 sg13g2_fill_1 FILLER_26_156 ();
 sg13g2_decap_8 FILLER_26_162 ();
 sg13g2_fill_1 FILLER_26_169 ();
 sg13g2_decap_4 FILLER_26_179 ();
 sg13g2_fill_1 FILLER_26_183 ();
 sg13g2_fill_2 FILLER_26_198 ();
 sg13g2_fill_1 FILLER_26_200 ();
 sg13g2_decap_4 FILLER_26_300 ();
 sg13g2_fill_1 FILLER_26_304 ();
 sg13g2_decap_8 FILLER_26_310 ();
 sg13g2_fill_1 FILLER_26_331 ();
 sg13g2_fill_1 FILLER_26_345 ();
 sg13g2_decap_4 FILLER_26_363 ();
 sg13g2_fill_1 FILLER_26_376 ();
 sg13g2_decap_8 FILLER_26_402 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_fill_2 FILLER_27_84 ();
 sg13g2_fill_1 FILLER_27_86 ();
 sg13g2_fill_1 FILLER_27_113 ();
 sg13g2_fill_2 FILLER_27_150 ();
 sg13g2_fill_1 FILLER_27_152 ();
 sg13g2_decap_4 FILLER_27_205 ();
 sg13g2_decap_8 FILLER_27_232 ();
 sg13g2_fill_1 FILLER_27_239 ();
 sg13g2_fill_1 FILLER_27_250 ();
 sg13g2_decap_4 FILLER_27_261 ();
 sg13g2_fill_2 FILLER_27_265 ();
 sg13g2_decap_4 FILLER_27_271 ();
 sg13g2_decap_4 FILLER_27_278 ();
 sg13g2_fill_2 FILLER_27_282 ();
 sg13g2_fill_1 FILLER_27_348 ();
 sg13g2_fill_1 FILLER_27_380 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_4 FILLER_28_91 ();
 sg13g2_fill_2 FILLER_28_95 ();
 sg13g2_decap_4 FILLER_28_114 ();
 sg13g2_decap_8 FILLER_28_123 ();
 sg13g2_decap_8 FILLER_28_134 ();
 sg13g2_decap_4 FILLER_28_141 ();
 sg13g2_fill_2 FILLER_28_145 ();
 sg13g2_fill_2 FILLER_28_161 ();
 sg13g2_fill_1 FILLER_28_163 ();
 sg13g2_fill_2 FILLER_28_168 ();
 sg13g2_decap_8 FILLER_28_174 ();
 sg13g2_decap_8 FILLER_28_181 ();
 sg13g2_fill_2 FILLER_28_188 ();
 sg13g2_decap_4 FILLER_28_194 ();
 sg13g2_fill_1 FILLER_28_198 ();
 sg13g2_decap_4 FILLER_28_244 ();
 sg13g2_fill_1 FILLER_28_248 ();
 sg13g2_fill_1 FILLER_28_275 ();
 sg13g2_fill_1 FILLER_28_285 ();
 sg13g2_decap_8 FILLER_28_291 ();
 sg13g2_decap_4 FILLER_28_310 ();
 sg13g2_fill_1 FILLER_28_314 ();
 sg13g2_fill_2 FILLER_28_328 ();
 sg13g2_fill_1 FILLER_28_330 ();
 sg13g2_fill_1 FILLER_28_340 ();
 sg13g2_decap_8 FILLER_28_350 ();
 sg13g2_decap_8 FILLER_28_357 ();
 sg13g2_fill_1 FILLER_28_364 ();
 sg13g2_decap_4 FILLER_28_369 ();
 sg13g2_fill_1 FILLER_28_373 ();
 sg13g2_decap_8 FILLER_28_379 ();
 sg13g2_decap_4 FILLER_28_403 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_4 FILLER_29_91 ();
 sg13g2_fill_1 FILLER_29_121 ();
 sg13g2_decap_4 FILLER_29_132 ();
 sg13g2_fill_1 FILLER_29_136 ();
 sg13g2_fill_2 FILLER_29_162 ();
 sg13g2_fill_1 FILLER_29_164 ();
 sg13g2_decap_4 FILLER_29_186 ();
 sg13g2_fill_2 FILLER_29_190 ();
 sg13g2_decap_4 FILLER_29_213 ();
 sg13g2_fill_1 FILLER_29_217 ();
 sg13g2_fill_1 FILLER_29_251 ();
 sg13g2_fill_2 FILLER_29_270 ();
 sg13g2_fill_2 FILLER_29_292 ();
 sg13g2_fill_1 FILLER_29_294 ();
 sg13g2_decap_4 FILLER_29_316 ();
 sg13g2_fill_2 FILLER_29_320 ();
 sg13g2_fill_1 FILLER_29_335 ();
 sg13g2_fill_2 FILLER_29_380 ();
 sg13g2_fill_1 FILLER_29_382 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_4 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_fill_2 FILLER_30_140 ();
 sg13g2_fill_1 FILLER_30_142 ();
 sg13g2_decap_8 FILLER_30_153 ();
 sg13g2_decap_8 FILLER_30_160 ();
 sg13g2_fill_2 FILLER_30_167 ();
 sg13g2_fill_1 FILLER_30_169 ();
 sg13g2_decap_8 FILLER_30_180 ();
 sg13g2_decap_4 FILLER_30_187 ();
 sg13g2_fill_1 FILLER_30_191 ();
 sg13g2_decap_8 FILLER_30_206 ();
 sg13g2_decap_8 FILLER_30_213 ();
 sg13g2_decap_8 FILLER_30_220 ();
 sg13g2_decap_4 FILLER_30_234 ();
 sg13g2_decap_8 FILLER_30_254 ();
 sg13g2_fill_2 FILLER_30_261 ();
 sg13g2_decap_8 FILLER_30_272 ();
 sg13g2_fill_2 FILLER_30_279 ();
 sg13g2_decap_8 FILLER_30_293 ();
 sg13g2_fill_2 FILLER_30_300 ();
 sg13g2_fill_2 FILLER_30_307 ();
 sg13g2_fill_1 FILLER_30_309 ();
 sg13g2_decap_8 FILLER_30_315 ();
 sg13g2_decap_8 FILLER_30_322 ();
 sg13g2_fill_1 FILLER_30_329 ();
 sg13g2_decap_8 FILLER_30_338 ();
 sg13g2_decap_4 FILLER_30_345 ();
 sg13g2_fill_2 FILLER_30_349 ();
 sg13g2_decap_4 FILLER_30_364 ();
 sg13g2_fill_2 FILLER_30_368 ();
 sg13g2_fill_2 FILLER_30_406 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_4 FILLER_31_84 ();
 sg13g2_fill_2 FILLER_31_88 ();
 sg13g2_fill_2 FILLER_31_116 ();
 sg13g2_fill_1 FILLER_31_118 ();
 sg13g2_fill_2 FILLER_31_128 ();
 sg13g2_fill_1 FILLER_31_130 ();
 sg13g2_decap_8 FILLER_31_160 ();
 sg13g2_decap_4 FILLER_31_167 ();
 sg13g2_fill_2 FILLER_31_171 ();
 sg13g2_decap_8 FILLER_31_180 ();
 sg13g2_fill_2 FILLER_31_187 ();
 sg13g2_decap_8 FILLER_31_208 ();
 sg13g2_decap_4 FILLER_31_215 ();
 sg13g2_decap_8 FILLER_31_226 ();
 sg13g2_fill_2 FILLER_31_233 ();
 sg13g2_fill_1 FILLER_31_235 ();
 sg13g2_fill_2 FILLER_31_243 ();
 sg13g2_fill_2 FILLER_31_251 ();
 sg13g2_fill_1 FILLER_31_253 ();
 sg13g2_fill_2 FILLER_31_259 ();
 sg13g2_decap_4 FILLER_31_278 ();
 sg13g2_fill_1 FILLER_31_282 ();
 sg13g2_decap_4 FILLER_31_293 ();
 sg13g2_fill_1 FILLER_31_297 ();
 sg13g2_fill_2 FILLER_31_313 ();
 sg13g2_fill_1 FILLER_31_315 ();
 sg13g2_fill_2 FILLER_31_337 ();
 sg13g2_fill_1 FILLER_31_339 ();
 sg13g2_decap_8 FILLER_31_356 ();
 sg13g2_fill_2 FILLER_31_363 ();
 sg13g2_fill_1 FILLER_31_365 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_fill_2 FILLER_32_98 ();
 sg13g2_fill_2 FILLER_32_113 ();
 sg13g2_fill_2 FILLER_32_137 ();
 sg13g2_fill_1 FILLER_32_139 ();
 sg13g2_decap_8 FILLER_32_150 ();
 sg13g2_fill_2 FILLER_32_157 ();
 sg13g2_decap_4 FILLER_32_208 ();
 sg13g2_fill_2 FILLER_32_232 ();
 sg13g2_fill_1 FILLER_32_234 ();
 sg13g2_decap_8 FILLER_32_248 ();
 sg13g2_decap_8 FILLER_32_255 ();
 sg13g2_fill_2 FILLER_32_262 ();
 sg13g2_fill_1 FILLER_32_264 ();
 sg13g2_decap_8 FILLER_32_273 ();
 sg13g2_decap_8 FILLER_32_280 ();
 sg13g2_decap_8 FILLER_32_295 ();
 sg13g2_decap_4 FILLER_32_302 ();
 sg13g2_fill_2 FILLER_32_306 ();
 sg13g2_decap_8 FILLER_32_325 ();
 sg13g2_decap_8 FILLER_32_354 ();
 sg13g2_fill_1 FILLER_32_361 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_fill_2 FILLER_33_91 ();
 sg13g2_fill_2 FILLER_33_97 ();
 sg13g2_fill_1 FILLER_33_99 ();
 sg13g2_decap_8 FILLER_33_129 ();
 sg13g2_decap_8 FILLER_33_149 ();
 sg13g2_decap_4 FILLER_33_156 ();
 sg13g2_fill_1 FILLER_33_160 ();
 sg13g2_decap_8 FILLER_33_166 ();
 sg13g2_fill_2 FILLER_33_173 ();
 sg13g2_fill_1 FILLER_33_175 ();
 sg13g2_fill_2 FILLER_33_180 ();
 sg13g2_fill_1 FILLER_33_182 ();
 sg13g2_fill_2 FILLER_33_191 ();
 sg13g2_fill_1 FILLER_33_193 ();
 sg13g2_decap_8 FILLER_33_199 ();
 sg13g2_decap_8 FILLER_33_206 ();
 sg13g2_decap_8 FILLER_33_213 ();
 sg13g2_fill_2 FILLER_33_220 ();
 sg13g2_fill_1 FILLER_33_222 ();
 sg13g2_decap_4 FILLER_33_227 ();
 sg13g2_fill_1 FILLER_33_284 ();
 sg13g2_fill_2 FILLER_33_305 ();
 sg13g2_decap_8 FILLER_33_324 ();
 sg13g2_decap_8 FILLER_33_331 ();
 sg13g2_fill_1 FILLER_33_338 ();
 sg13g2_decap_8 FILLER_33_351 ();
 sg13g2_decap_4 FILLER_33_358 ();
 sg13g2_fill_1 FILLER_33_362 ();
 sg13g2_decap_8 FILLER_33_373 ();
 sg13g2_decap_8 FILLER_33_380 ();
 sg13g2_decap_4 FILLER_33_403 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_4 FILLER_34_77 ();
 sg13g2_fill_1 FILLER_34_81 ();
 sg13g2_fill_1 FILLER_34_108 ();
 sg13g2_decap_4 FILLER_34_118 ();
 sg13g2_fill_2 FILLER_34_130 ();
 sg13g2_fill_2 FILLER_34_152 ();
 sg13g2_fill_1 FILLER_34_154 ();
 sg13g2_fill_2 FILLER_34_176 ();
 sg13g2_decap_8 FILLER_34_225 ();
 sg13g2_decap_8 FILLER_34_232 ();
 sg13g2_decap_4 FILLER_34_239 ();
 sg13g2_fill_1 FILLER_34_243 ();
 sg13g2_decap_4 FILLER_34_258 ();
 sg13g2_fill_1 FILLER_34_262 ();
 sg13g2_decap_8 FILLER_34_276 ();
 sg13g2_decap_8 FILLER_34_283 ();
 sg13g2_fill_1 FILLER_34_290 ();
 sg13g2_decap_8 FILLER_34_299 ();
 sg13g2_decap_4 FILLER_34_306 ();
 sg13g2_fill_1 FILLER_34_310 ();
 sg13g2_fill_2 FILLER_34_327 ();
 sg13g2_fill_1 FILLER_34_329 ();
 sg13g2_decap_4 FILLER_34_350 ();
 sg13g2_fill_1 FILLER_34_354 ();
 sg13g2_decap_4 FILLER_34_376 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_4 FILLER_35_98 ();
 sg13g2_fill_2 FILLER_35_116 ();
 sg13g2_fill_1 FILLER_35_122 ();
 sg13g2_decap_8 FILLER_35_128 ();
 sg13g2_decap_4 FILLER_35_135 ();
 sg13g2_fill_1 FILLER_35_139 ();
 sg13g2_decap_8 FILLER_35_148 ();
 sg13g2_decap_4 FILLER_35_155 ();
 sg13g2_fill_1 FILLER_35_159 ();
 sg13g2_decap_4 FILLER_35_165 ();
 sg13g2_fill_1 FILLER_35_169 ();
 sg13g2_decap_4 FILLER_35_176 ();
 sg13g2_fill_2 FILLER_35_180 ();
 sg13g2_decap_8 FILLER_35_194 ();
 sg13g2_decap_8 FILLER_35_201 ();
 sg13g2_decap_4 FILLER_35_208 ();
 sg13g2_fill_1 FILLER_35_230 ();
 sg13g2_fill_2 FILLER_35_236 ();
 sg13g2_decap_4 FILLER_35_243 ();
 sg13g2_decap_4 FILLER_35_284 ();
 sg13g2_fill_2 FILLER_35_288 ();
 sg13g2_fill_2 FILLER_35_303 ();
 sg13g2_fill_1 FILLER_35_305 ();
 sg13g2_fill_2 FILLER_35_314 ();
 sg13g2_decap_8 FILLER_35_328 ();
 sg13g2_fill_1 FILLER_35_335 ();
 sg13g2_decap_8 FILLER_35_344 ();
 sg13g2_fill_1 FILLER_35_351 ();
 sg13g2_decap_8 FILLER_35_356 ();
 sg13g2_fill_2 FILLER_35_371 ();
 sg13g2_fill_1 FILLER_35_373 ();
 sg13g2_decap_8 FILLER_35_379 ();
 sg13g2_decap_8 FILLER_35_386 ();
 sg13g2_fill_1 FILLER_35_393 ();
 sg13g2_decap_4 FILLER_35_403 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_fill_1 FILLER_36_110 ();
 sg13g2_decap_8 FILLER_36_120 ();
 sg13g2_decap_4 FILLER_36_127 ();
 sg13g2_fill_1 FILLER_36_131 ();
 sg13g2_decap_4 FILLER_36_147 ();
 sg13g2_decap_4 FILLER_36_159 ();
 sg13g2_fill_2 FILLER_36_163 ();
 sg13g2_fill_2 FILLER_36_172 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_fill_1 FILLER_36_196 ();
 sg13g2_fill_2 FILLER_36_201 ();
 sg13g2_fill_1 FILLER_36_203 ();
 sg13g2_decap_4 FILLER_36_210 ();
 sg13g2_fill_1 FILLER_36_214 ();
 sg13g2_fill_2 FILLER_36_219 ();
 sg13g2_fill_1 FILLER_36_221 ();
 sg13g2_decap_8 FILLER_36_234 ();
 sg13g2_decap_4 FILLER_36_241 ();
 sg13g2_fill_1 FILLER_36_245 ();
 sg13g2_decap_4 FILLER_36_256 ();
 sg13g2_fill_1 FILLER_36_260 ();
 sg13g2_decap_4 FILLER_36_283 ();
 sg13g2_fill_1 FILLER_36_287 ();
 sg13g2_decap_4 FILLER_36_295 ();
 sg13g2_fill_2 FILLER_36_299 ();
 sg13g2_decap_8 FILLER_36_315 ();
 sg13g2_fill_2 FILLER_36_322 ();
 sg13g2_fill_1 FILLER_36_324 ();
 sg13g2_decap_8 FILLER_36_330 ();
 sg13g2_decap_4 FILLER_36_337 ();
 sg13g2_fill_2 FILLER_36_341 ();
 sg13g2_fill_2 FILLER_36_347 ();
 sg13g2_fill_2 FILLER_36_363 ();
 sg13g2_fill_1 FILLER_36_365 ();
 sg13g2_fill_2 FILLER_36_381 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_4 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_99 ();
 sg13g2_decap_4 FILLER_37_106 ();
 sg13g2_decap_4 FILLER_37_115 ();
 sg13g2_fill_1 FILLER_37_119 ();
 sg13g2_fill_2 FILLER_37_132 ();
 sg13g2_fill_2 FILLER_37_148 ();
 sg13g2_fill_1 FILLER_37_158 ();
 sg13g2_decap_4 FILLER_37_186 ();
 sg13g2_fill_2 FILLER_37_190 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_fill_1 FILLER_37_222 ();
 sg13g2_decap_8 FILLER_37_236 ();
 sg13g2_fill_2 FILLER_37_304 ();
 sg13g2_fill_1 FILLER_37_306 ();
 sg13g2_fill_2 FILLER_37_320 ();
 sg13g2_fill_1 FILLER_37_322 ();
 sg13g2_fill_1 FILLER_37_342 ();
 sg13g2_decap_8 FILLER_37_375 ();
 sg13g2_fill_2 FILLER_37_382 ();
 sg13g2_fill_1 FILLER_37_384 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_fill_1 FILLER_38_100 ();
 sg13g2_fill_2 FILLER_38_139 ();
 sg13g2_fill_1 FILLER_38_141 ();
 sg13g2_decap_4 FILLER_38_176 ();
 sg13g2_fill_1 FILLER_38_180 ();
 sg13g2_decap_4 FILLER_38_207 ();
 sg13g2_fill_2 FILLER_38_211 ();
 sg13g2_decap_8 FILLER_38_239 ();
 sg13g2_fill_2 FILLER_38_246 ();
 sg13g2_fill_1 FILLER_38_248 ();
 sg13g2_decap_4 FILLER_38_275 ();
 sg13g2_fill_2 FILLER_38_279 ();
 sg13g2_decap_8 FILLER_38_285 ();
 sg13g2_decap_8 FILLER_38_292 ();
 sg13g2_decap_4 FILLER_38_299 ();
 sg13g2_fill_2 FILLER_38_303 ();
 sg13g2_fill_2 FILLER_38_327 ();
 sg13g2_fill_2 FILLER_38_334 ();
 sg13g2_fill_1 FILLER_38_349 ();
 sg13g2_fill_2 FILLER_38_365 ();
 sg13g2_fill_1 FILLER_38_367 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net111;
 assign uio_oe[1] = net11;
 assign uio_oe[2] = net12;
 assign uio_oe[3] = net13;
 assign uio_oe[4] = net14;
 assign uio_oe[5] = net15;
 assign uio_oe[6] = net16;
 assign uio_oe[7] = net17;
 assign uio_out[1] = net18;
 assign uio_out[2] = net19;
 assign uio_out[3] = net20;
 assign uio_out[4] = net21;
 assign uio_out[5] = net22;
 assign uio_out[6] = net23;
 assign uio_out[7] = net24;
endmodule
