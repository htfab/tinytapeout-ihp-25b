module tt_um_2048_vga_game (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire _4209_;
 wire _4210_;
 wire _4211_;
 wire _4212_;
 wire _4213_;
 wire _4214_;
 wire _4215_;
 wire _4216_;
 wire _4217_;
 wire _4218_;
 wire _4219_;
 wire _4220_;
 wire _4221_;
 wire _4222_;
 wire _4223_;
 wire _4224_;
 wire _4225_;
 wire _4226_;
 wire _4227_;
 wire _4228_;
 wire _4229_;
 wire _4230_;
 wire _4231_;
 wire _4232_;
 wire _4233_;
 wire _4234_;
 wire _4235_;
 wire _4236_;
 wire _4237_;
 wire _4238_;
 wire _4239_;
 wire _4240_;
 wire _4241_;
 wire _4242_;
 wire _4243_;
 wire _4244_;
 wire _4245_;
 wire _4246_;
 wire _4247_;
 wire _4248_;
 wire _4249_;
 wire _4250_;
 wire _4251_;
 wire _4252_;
 wire _4253_;
 wire _4254_;
 wire _4255_;
 wire _4256_;
 wire _4257_;
 wire _4258_;
 wire _4259_;
 wire _4260_;
 wire _4261_;
 wire _4262_;
 wire _4263_;
 wire _4264_;
 wire _4265_;
 wire _4266_;
 wire _4267_;
 wire _4268_;
 wire _4269_;
 wire _4270_;
 wire _4271_;
 wire _4272_;
 wire _4273_;
 wire _4274_;
 wire _4275_;
 wire _4276_;
 wire _4277_;
 wire _4278_;
 wire _4279_;
 wire _4280_;
 wire _4281_;
 wire _4282_;
 wire _4283_;
 wire _4284_;
 wire _4285_;
 wire _4286_;
 wire _4287_;
 wire _4288_;
 wire _4289_;
 wire _4290_;
 wire _4291_;
 wire _4292_;
 wire _4293_;
 wire _4294_;
 wire _4295_;
 wire _4296_;
 wire _4297_;
 wire _4298_;
 wire _4299_;
 wire _4300_;
 wire _4301_;
 wire _4302_;
 wire _4303_;
 wire _4304_;
 wire _4305_;
 wire _4306_;
 wire _4307_;
 wire _4308_;
 wire _4309_;
 wire _4310_;
 wire _4311_;
 wire _4312_;
 wire _4313_;
 wire _4314_;
 wire _4315_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire clknet_leaf_0_clk;
 wire \btn_down_debounce.button_sync_0 ;
 wire \btn_down_debounce.button_sync_1 ;
 wire \btn_down_debounce.debounce_counter[0] ;
 wire \btn_down_debounce.debounce_counter[10] ;
 wire \btn_down_debounce.debounce_counter[11] ;
 wire \btn_down_debounce.debounce_counter[12] ;
 wire \btn_down_debounce.debounce_counter[13] ;
 wire \btn_down_debounce.debounce_counter[14] ;
 wire \btn_down_debounce.debounce_counter[15] ;
 wire \btn_down_debounce.debounce_counter[16] ;
 wire \btn_down_debounce.debounce_counter[17] ;
 wire \btn_down_debounce.debounce_counter[1] ;
 wire \btn_down_debounce.debounce_counter[2] ;
 wire \btn_down_debounce.debounce_counter[3] ;
 wire \btn_down_debounce.debounce_counter[4] ;
 wire \btn_down_debounce.debounce_counter[5] ;
 wire \btn_down_debounce.debounce_counter[6] ;
 wire \btn_down_debounce.debounce_counter[7] ;
 wire \btn_down_debounce.debounce_counter[8] ;
 wire \btn_down_debounce.debounce_counter[9] ;
 wire \btn_down_debounce.debounced ;
 wire \btn_left_debounce.button_sync_0 ;
 wire \btn_left_debounce.button_sync_1 ;
 wire \btn_left_debounce.debounce_counter[0] ;
 wire \btn_left_debounce.debounce_counter[10] ;
 wire \btn_left_debounce.debounce_counter[11] ;
 wire \btn_left_debounce.debounce_counter[12] ;
 wire \btn_left_debounce.debounce_counter[13] ;
 wire \btn_left_debounce.debounce_counter[14] ;
 wire \btn_left_debounce.debounce_counter[15] ;
 wire \btn_left_debounce.debounce_counter[16] ;
 wire \btn_left_debounce.debounce_counter[17] ;
 wire \btn_left_debounce.debounce_counter[1] ;
 wire \btn_left_debounce.debounce_counter[2] ;
 wire \btn_left_debounce.debounce_counter[3] ;
 wire \btn_left_debounce.debounce_counter[4] ;
 wire \btn_left_debounce.debounce_counter[5] ;
 wire \btn_left_debounce.debounce_counter[6] ;
 wire \btn_left_debounce.debounce_counter[7] ;
 wire \btn_left_debounce.debounce_counter[8] ;
 wire \btn_left_debounce.debounce_counter[9] ;
 wire \btn_left_debounce.debounced ;
 wire \btn_right_debounce.button_sync_0 ;
 wire \btn_right_debounce.button_sync_1 ;
 wire \btn_right_debounce.debounce_counter[0] ;
 wire \btn_right_debounce.debounce_counter[10] ;
 wire \btn_right_debounce.debounce_counter[11] ;
 wire \btn_right_debounce.debounce_counter[12] ;
 wire \btn_right_debounce.debounce_counter[13] ;
 wire \btn_right_debounce.debounce_counter[14] ;
 wire \btn_right_debounce.debounce_counter[15] ;
 wire \btn_right_debounce.debounce_counter[16] ;
 wire \btn_right_debounce.debounce_counter[17] ;
 wire \btn_right_debounce.debounce_counter[1] ;
 wire \btn_right_debounce.debounce_counter[2] ;
 wire \btn_right_debounce.debounce_counter[3] ;
 wire \btn_right_debounce.debounce_counter[4] ;
 wire \btn_right_debounce.debounce_counter[5] ;
 wire \btn_right_debounce.debounce_counter[6] ;
 wire \btn_right_debounce.debounce_counter[7] ;
 wire \btn_right_debounce.debounce_counter[8] ;
 wire \btn_right_debounce.debounce_counter[9] ;
 wire \btn_right_debounce.debounced ;
 wire btn_select_prev;
 wire \btn_up_debounce.button_sync_0 ;
 wire \btn_up_debounce.button_sync_1 ;
 wire \btn_up_debounce.debounce_counter[0] ;
 wire \btn_up_debounce.debounce_counter[10] ;
 wire \btn_up_debounce.debounce_counter[11] ;
 wire \btn_up_debounce.debounce_counter[12] ;
 wire \btn_up_debounce.debounce_counter[13] ;
 wire \btn_up_debounce.debounce_counter[14] ;
 wire \btn_up_debounce.debounce_counter[15] ;
 wire \btn_up_debounce.debounce_counter[16] ;
 wire \btn_up_debounce.debounce_counter[17] ;
 wire \btn_up_debounce.debounce_counter[1] ;
 wire \btn_up_debounce.debounce_counter[2] ;
 wire \btn_up_debounce.debounce_counter[3] ;
 wire \btn_up_debounce.debounce_counter[4] ;
 wire \btn_up_debounce.debounce_counter[5] ;
 wire \btn_up_debounce.debounce_counter[6] ;
 wire \btn_up_debounce.debounce_counter[7] ;
 wire \btn_up_debounce.debounce_counter[8] ;
 wire \btn_up_debounce.debounce_counter[9] ;
 wire \btn_up_debounce.debounced ;
 wire debug_btn_down;
 wire debug_btn_left;
 wire debug_btn_right;
 wire debug_btn_up;
 wire \debug_controller_inst.data_out_en ;
 wire \debug_controller_inst.grid_addr[0] ;
 wire \debug_controller_inst.grid_addr[1] ;
 wire \debug_controller_inst.grid_addr[2] ;
 wire \debug_controller_inst.grid_addr[3] ;
 wire \debug_controller_inst.grid_in[0] ;
 wire \debug_controller_inst.grid_in[10] ;
 wire \debug_controller_inst.grid_in[11] ;
 wire \debug_controller_inst.grid_in[12] ;
 wire \debug_controller_inst.grid_in[13] ;
 wire \debug_controller_inst.grid_in[14] ;
 wire \debug_controller_inst.grid_in[15] ;
 wire \debug_controller_inst.grid_in[16] ;
 wire \debug_controller_inst.grid_in[17] ;
 wire \debug_controller_inst.grid_in[18] ;
 wire \debug_controller_inst.grid_in[19] ;
 wire \debug_controller_inst.grid_in[1] ;
 wire \debug_controller_inst.grid_in[20] ;
 wire \debug_controller_inst.grid_in[21] ;
 wire \debug_controller_inst.grid_in[22] ;
 wire \debug_controller_inst.grid_in[23] ;
 wire \debug_controller_inst.grid_in[24] ;
 wire \debug_controller_inst.grid_in[25] ;
 wire \debug_controller_inst.grid_in[26] ;
 wire \debug_controller_inst.grid_in[27] ;
 wire \debug_controller_inst.grid_in[28] ;
 wire \debug_controller_inst.grid_in[29] ;
 wire \debug_controller_inst.grid_in[2] ;
 wire \debug_controller_inst.grid_in[30] ;
 wire \debug_controller_inst.grid_in[31] ;
 wire \debug_controller_inst.grid_in[32] ;
 wire \debug_controller_inst.grid_in[33] ;
 wire \debug_controller_inst.grid_in[34] ;
 wire \debug_controller_inst.grid_in[35] ;
 wire \debug_controller_inst.grid_in[36] ;
 wire \debug_controller_inst.grid_in[37] ;
 wire \debug_controller_inst.grid_in[38] ;
 wire \debug_controller_inst.grid_in[39] ;
 wire \debug_controller_inst.grid_in[3] ;
 wire \debug_controller_inst.grid_in[40] ;
 wire \debug_controller_inst.grid_in[41] ;
 wire \debug_controller_inst.grid_in[42] ;
 wire \debug_controller_inst.grid_in[43] ;
 wire \debug_controller_inst.grid_in[44] ;
 wire \debug_controller_inst.grid_in[45] ;
 wire \debug_controller_inst.grid_in[46] ;
 wire \debug_controller_inst.grid_in[47] ;
 wire \debug_controller_inst.grid_in[48] ;
 wire \debug_controller_inst.grid_in[49] ;
 wire \debug_controller_inst.grid_in[4] ;
 wire \debug_controller_inst.grid_in[50] ;
 wire \debug_controller_inst.grid_in[51] ;
 wire \debug_controller_inst.grid_in[52] ;
 wire \debug_controller_inst.grid_in[53] ;
 wire \debug_controller_inst.grid_in[54] ;
 wire \debug_controller_inst.grid_in[55] ;
 wire \debug_controller_inst.grid_in[56] ;
 wire \debug_controller_inst.grid_in[57] ;
 wire \debug_controller_inst.grid_in[58] ;
 wire \debug_controller_inst.grid_in[59] ;
 wire \debug_controller_inst.grid_in[5] ;
 wire \debug_controller_inst.grid_in[60] ;
 wire \debug_controller_inst.grid_in[61] ;
 wire \debug_controller_inst.grid_in[62] ;
 wire \debug_controller_inst.grid_in[63] ;
 wire \debug_controller_inst.grid_in[6] ;
 wire \debug_controller_inst.grid_in[7] ;
 wire \debug_controller_inst.grid_in[8] ;
 wire \debug_controller_inst.grid_in[9] ;
 wire \debug_controller_inst.grid_out_addr[0] ;
 wire \debug_controller_inst.grid_out_addr[1] ;
 wire \debug_controller_inst.grid_out_addr[2] ;
 wire \debug_controller_inst.grid_out_addr[3] ;
 wire \debug_controller_inst.grid_out_data[0] ;
 wire \debug_controller_inst.grid_out_data[1] ;
 wire \debug_controller_inst.grid_out_data[2] ;
 wire \debug_controller_inst.grid_out_data[3] ;
 wire \debug_controller_inst.grid_out_valid ;
 wire \draw_game_inst.board_x[0] ;
 wire \draw_game_inst.board_x[1] ;
 wire \draw_game_inst.board_x[2] ;
 wire \draw_game_inst.board_x[3] ;
 wire \draw_game_inst.board_x[4] ;
 wire \draw_game_inst.board_x[5] ;
 wire \draw_game_inst.board_y[0] ;
 wire \draw_game_inst.board_y[1] ;
 wire \draw_game_inst.board_y[2] ;
 wire \draw_game_inst.board_y[3] ;
 wire \draw_game_inst.board_y[4] ;
 wire \draw_game_inst.board_y[5] ;
 wire \draw_game_inst.board_y[6] ;
 wire \draw_game_inst.grid[0] ;
 wire \draw_game_inst.grid[10] ;
 wire \draw_game_inst.grid[11] ;
 wire \draw_game_inst.grid[12] ;
 wire \draw_game_inst.grid[13] ;
 wire \draw_game_inst.grid[14] ;
 wire \draw_game_inst.grid[15] ;
 wire \draw_game_inst.grid[16] ;
 wire \draw_game_inst.grid[17] ;
 wire \draw_game_inst.grid[18] ;
 wire \draw_game_inst.grid[19] ;
 wire \draw_game_inst.grid[1] ;
 wire \draw_game_inst.grid[20] ;
 wire \draw_game_inst.grid[21] ;
 wire \draw_game_inst.grid[22] ;
 wire \draw_game_inst.grid[23] ;
 wire \draw_game_inst.grid[24] ;
 wire \draw_game_inst.grid[25] ;
 wire \draw_game_inst.grid[26] ;
 wire \draw_game_inst.grid[27] ;
 wire \draw_game_inst.grid[28] ;
 wire \draw_game_inst.grid[29] ;
 wire \draw_game_inst.grid[2] ;
 wire \draw_game_inst.grid[30] ;
 wire \draw_game_inst.grid[31] ;
 wire \draw_game_inst.grid[32] ;
 wire \draw_game_inst.grid[33] ;
 wire \draw_game_inst.grid[34] ;
 wire \draw_game_inst.grid[35] ;
 wire \draw_game_inst.grid[36] ;
 wire \draw_game_inst.grid[37] ;
 wire \draw_game_inst.grid[38] ;
 wire \draw_game_inst.grid[39] ;
 wire \draw_game_inst.grid[3] ;
 wire \draw_game_inst.grid[40] ;
 wire \draw_game_inst.grid[41] ;
 wire \draw_game_inst.grid[42] ;
 wire \draw_game_inst.grid[43] ;
 wire \draw_game_inst.grid[44] ;
 wire \draw_game_inst.grid[45] ;
 wire \draw_game_inst.grid[46] ;
 wire \draw_game_inst.grid[47] ;
 wire \draw_game_inst.grid[48] ;
 wire \draw_game_inst.grid[49] ;
 wire \draw_game_inst.grid[4] ;
 wire \draw_game_inst.grid[50] ;
 wire \draw_game_inst.grid[51] ;
 wire \draw_game_inst.grid[52] ;
 wire \draw_game_inst.grid[53] ;
 wire \draw_game_inst.grid[54] ;
 wire \draw_game_inst.grid[55] ;
 wire \draw_game_inst.grid[56] ;
 wire \draw_game_inst.grid[57] ;
 wire \draw_game_inst.grid[58] ;
 wire \draw_game_inst.grid[59] ;
 wire \draw_game_inst.grid[5] ;
 wire \draw_game_inst.grid[60] ;
 wire \draw_game_inst.grid[61] ;
 wire \draw_game_inst.grid[62] ;
 wire \draw_game_inst.grid[63] ;
 wire \draw_game_inst.grid[6] ;
 wire \draw_game_inst.grid[7] ;
 wire \draw_game_inst.grid[8] ;
 wire \draw_game_inst.grid[9] ;
 wire \draw_game_inst.new_tiles[0] ;
 wire \draw_game_inst.new_tiles[10] ;
 wire \draw_game_inst.new_tiles[11] ;
 wire \draw_game_inst.new_tiles[12] ;
 wire \draw_game_inst.new_tiles[13] ;
 wire \draw_game_inst.new_tiles[14] ;
 wire \draw_game_inst.new_tiles[15] ;
 wire \draw_game_inst.new_tiles[1] ;
 wire \draw_game_inst.new_tiles[2] ;
 wire \draw_game_inst.new_tiles[3] ;
 wire \draw_game_inst.new_tiles[4] ;
 wire \draw_game_inst.new_tiles[5] ;
 wire \draw_game_inst.new_tiles[6] ;
 wire \draw_game_inst.new_tiles[7] ;
 wire \draw_game_inst.new_tiles[8] ;
 wire \draw_game_inst.new_tiles[9] ;
 wire \draw_game_inst.new_tiles_counter[0] ;
 wire \draw_game_inst.new_tiles_counter[1] ;
 wire \draw_game_inst.new_tiles_counter[2] ;
 wire \draw_game_inst.x[6] ;
 wire \draw_game_inst.x[7] ;
 wire \draw_game_inst.x[8] ;
 wire \draw_game_inst.x[9] ;
 wire \draw_game_inst.y[7] ;
 wire \draw_game_inst.y[8] ;
 wire \draw_game_inst.y[9] ;
 wire \game_logic_inst.add_new_tiles[0] ;
 wire \game_logic_inst.add_new_tiles[1] ;
 wire \game_logic_inst.added_tile_index[0] ;
 wire \game_logic_inst.added_tile_index[1] ;
 wire \game_logic_inst.added_tile_index[2] ;
 wire \game_logic_inst.added_tile_index[3] ;
 wire \game_logic_inst.calculate_move ;
 wire \game_logic_inst.current_direction[1] ;
 wire \game_logic_inst.current_direction[2] ;
 wire \game_logic_inst.current_direction[3] ;
 wire \game_logic_inst.current_row_index[0] ;
 wire \game_logic_inst.current_row_index[1] ;
 wire \game_logic_inst.debug_move_reg ;
 wire \game_logic_inst.game_started ;
 wire \game_logic_inst.lfsr_shift[0] ;
 wire \game_logic_inst.lfsr_shift[1] ;
 wire \game_logic_inst.lfsr_value[0] ;
 wire \game_logic_inst.lfsr_value[10] ;
 wire \game_logic_inst.lfsr_value[11] ;
 wire \game_logic_inst.lfsr_value[12] ;
 wire \game_logic_inst.lfsr_value[13] ;
 wire \game_logic_inst.lfsr_value[14] ;
 wire \game_logic_inst.lfsr_value[15] ;
 wire \game_logic_inst.lfsr_value[1] ;
 wire \game_logic_inst.lfsr_value[2] ;
 wire \game_logic_inst.lfsr_value[3] ;
 wire \game_logic_inst.lfsr_value[4] ;
 wire \game_logic_inst.lfsr_value[5] ;
 wire \game_logic_inst.lfsr_value[6] ;
 wire \game_logic_inst.lfsr_value[7] ;
 wire \game_logic_inst.lfsr_value[8] ;
 wire \game_logic_inst.lfsr_value[9] ;
 wire \game_logic_inst.prev_any_button_pressed ;
 wire \game_logic_inst.should_transpose ;
 wire \game_logic_inst.valid_move ;
 wire \gamepad_pmod.decoder.data_reg[0] ;
 wire \gamepad_pmod.decoder.data_reg[10] ;
 wire \gamepad_pmod.decoder.data_reg[11] ;
 wire \gamepad_pmod.decoder.data_reg[1] ;
 wire \gamepad_pmod.decoder.data_reg[2] ;
 wire \gamepad_pmod.decoder.data_reg[3] ;
 wire \gamepad_pmod.decoder.data_reg[4] ;
 wire \gamepad_pmod.decoder.data_reg[5] ;
 wire \gamepad_pmod.decoder.data_reg[6] ;
 wire \gamepad_pmod.decoder.data_reg[7] ;
 wire \gamepad_pmod.decoder.data_reg[8] ;
 wire \gamepad_pmod.decoder.data_reg[9] ;
 wire \gamepad_pmod.driver.pmod_clk_prev ;
 wire \gamepad_pmod.driver.pmod_clk_sync[0] ;
 wire \gamepad_pmod.driver.pmod_clk_sync[1] ;
 wire \gamepad_pmod.driver.pmod_data_sync[0] ;
 wire \gamepad_pmod.driver.pmod_data_sync[1] ;
 wire \gamepad_pmod.driver.pmod_latch_prev ;
 wire \gamepad_pmod.driver.pmod_latch_sync[0] ;
 wire \gamepad_pmod.driver.pmod_latch_sync[1] ;
 wire \gamepad_pmod.driver.shift_reg[0] ;
 wire \gamepad_pmod.driver.shift_reg[10] ;
 wire \gamepad_pmod.driver.shift_reg[11] ;
 wire \gamepad_pmod.driver.shift_reg[1] ;
 wire \gamepad_pmod.driver.shift_reg[2] ;
 wire \gamepad_pmod.driver.shift_reg[3] ;
 wire \gamepad_pmod.driver.shift_reg[4] ;
 wire \gamepad_pmod.driver.shift_reg[5] ;
 wire \gamepad_pmod.driver.shift_reg[6] ;
 wire \gamepad_pmod.driver.shift_reg[7] ;
 wire \gamepad_pmod.driver.shift_reg[8] ;
 wire \gamepad_pmod.driver.shift_reg[9] ;
 wire hsync;
 wire \lfsr_inst.lfsr[16] ;
 wire \lfsr_inst.lfsr[17] ;
 wire \lfsr_inst.lfsr[18] ;
 wire \lfsr_inst.lfsr[19] ;
 wire \lfsr_inst.lfsr[20] ;
 wire \lfsr_inst.lfsr[21] ;
 wire \lfsr_inst.lfsr[22] ;
 wire \lfsr_inst.lfsr[23] ;
 wire \lfsr_inst.lfsr[24] ;
 wire \lfsr_inst.lfsr[25] ;
 wire \lfsr_inst.lfsr[26] ;
 wire \lfsr_inst.lfsr[27] ;
 wire \lfsr_inst.lfsr[28] ;
 wire \lfsr_inst.lfsr[29] ;
 wire \lfsr_inst.lfsr[30] ;
 wire \lfsr_inst.lfsr[31] ;
 wire \new_tiles_counter[0] ;
 wire \new_tiles_counter[4] ;
 wire retro_colors;
 wire show_welcome_screen;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire \vga_sync_gen.vsync ;
 wire vsync_prev;
 wire \welcome_screen_grid[0] ;
 wire \welcome_screen_grid[11] ;
 wire \welcome_screen_grid[12] ;
 wire \welcome_screen_grid[16] ;
 wire \welcome_screen_grid[20] ;
 wire \welcome_screen_grid[24] ;
 wire \welcome_screen_grid[28] ;
 wire \welcome_screen_grid[32] ;
 wire \welcome_screen_grid[36] ;
 wire \welcome_screen_grid[40] ;
 wire \welcome_screen_grid[44] ;
 wire \welcome_screen_grid[48] ;
 wire \welcome_screen_grid[4] ;
 wire \welcome_screen_grid[52] ;
 wire \welcome_screen_grid[56] ;
 wire \welcome_screen_grid[60] ;
 wire \welcome_screen_inst.welcome_counter[0] ;
 wire \welcome_screen_inst.welcome_counter[1] ;
 wire \welcome_screen_inst.welcome_counter[2] ;
 wire \welcome_screen_inst.welcome_counter[3] ;
 wire \welcome_screen_inst.welcome_counter[4] ;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;

 sg13g2_inv_2 _4707_ (.Y(_3929_),
    .A(\debug_controller_inst.grid_addr[3] ));
 sg13g2_inv_1 _4708_ (.Y(_3930_),
    .A(net2074));
 sg13g2_inv_2 _4709_ (.Y(_3931_),
    .A(net2077));
 sg13g2_inv_1 _4710_ (.Y(_3932_),
    .A(net2082));
 sg13g2_inv_1 _4711_ (.Y(_3933_),
    .A(net16));
 sg13g2_inv_1 _4712_ (.Y(_3934_),
    .A(net15));
 sg13g2_inv_1 _4713_ (.Y(_3935_),
    .A(net14));
 sg13g2_inv_1 _4714_ (.Y(_3936_),
    .A(net2093));
 sg13g2_inv_1 _4715_ (.Y(_3937_),
    .A(net13));
 sg13g2_inv_1 _4716_ (.Y(_3938_),
    .A(\game_logic_inst.should_transpose ));
 sg13g2_inv_1 _4717_ (.Y(_3939_),
    .A(\game_logic_inst.add_new_tiles[1] ));
 sg13g2_inv_4 _4718_ (.A(net2120),
    .Y(_3940_));
 sg13g2_inv_1 _4719_ (.Y(_3941_),
    .A(net804));
 sg13g2_inv_1 _4720_ (.Y(_3942_),
    .A(net625));
 sg13g2_inv_1 _4721_ (.Y(_3943_),
    .A(net766));
 sg13g2_inv_1 _4722_ (.Y(_3944_),
    .A(net773));
 sg13g2_inv_1 _4723_ (.Y(_3945_),
    .A(\gamepad_pmod.driver.shift_reg[8] ));
 sg13g2_inv_1 _4724_ (.Y(_3946_),
    .A(net477));
 sg13g2_inv_1 _4725_ (.Y(_3947_),
    .A(net768));
 sg13g2_inv_1 _4726_ (.Y(_3948_),
    .A(net662));
 sg13g2_inv_1 _4727_ (.Y(_3949_),
    .A(net727));
 sg13g2_inv_1 _4728_ (.Y(_3950_),
    .A(net771));
 sg13g2_inv_1 _4729_ (.Y(_3951_),
    .A(net785));
 sg13g2_inv_1 _4730_ (.Y(_3952_),
    .A(\gamepad_pmod.driver.shift_reg[1] ));
 sg13g2_inv_1 _4731_ (.Y(_3953_),
    .A(net714));
 sg13g2_inv_1 _4732_ (.Y(_3954_),
    .A(net486));
 sg13g2_inv_1 _4733_ (.Y(_3955_),
    .A(net685));
 sg13g2_inv_1 _4734_ (.Y(_3956_),
    .A(net823));
 sg13g2_inv_1 _4735_ (.Y(_3957_),
    .A(\btn_down_debounce.debounced ));
 sg13g2_inv_1 _4736_ (.Y(_3958_),
    .A(net876));
 sg13g2_inv_2 _4737_ (.Y(_3959_),
    .A(net432));
 sg13g2_inv_1 _4738_ (.Y(_3960_),
    .A(net2256));
 sg13g2_inv_1 _4739_ (.Y(_3961_),
    .A(net886));
 sg13g2_inv_1 _4740_ (.Y(_3962_),
    .A(\lfsr_inst.lfsr[31] ));
 sg13g2_inv_1 _4741_ (.Y(_3963_),
    .A(\draw_game_inst.board_x[0] ));
 sg13g2_inv_1 _4742_ (.Y(_3964_),
    .A(net497));
 sg13g2_inv_1 _4743_ (.Y(_3965_),
    .A(net550));
 sg13g2_inv_1 _4744_ (.Y(_3966_),
    .A(net469));
 sg13g2_inv_1 _4745_ (.Y(_3967_),
    .A(net465));
 sg13g2_inv_1 _4746_ (.Y(_3968_),
    .A(net683));
 sg13g2_inv_1 _4747_ (.Y(_3969_),
    .A(net648));
 sg13g2_inv_1 _4748_ (.Y(_3970_),
    .A(net705));
 sg13g2_inv_1 _4749_ (.Y(_3971_),
    .A(net677));
 sg13g2_inv_1 _4750_ (.Y(_3972_),
    .A(net703));
 sg13g2_inv_1 _4751_ (.Y(_3973_),
    .A(net758));
 sg13g2_inv_1 _4752_ (.Y(_3974_),
    .A(net467));
 sg13g2_inv_1 _4753_ (.Y(_3975_),
    .A(net531));
 sg13g2_inv_1 _4754_ (.Y(_3976_),
    .A(net8));
 sg13g2_inv_1 _4755_ (.Y(_3977_),
    .A(net2104));
 sg13g2_inv_4 _4756_ (.A(net2290),
    .Y(_3978_));
 sg13g2_inv_1 _4757_ (.Y(_3979_),
    .A(\debug_controller_inst.grid_in[20] ));
 sg13g2_inv_1 _4758_ (.Y(_3980_),
    .A(\debug_controller_inst.grid_in[52] ));
 sg13g2_inv_1 _4759_ (.Y(_3981_),
    .A(\debug_controller_inst.grid_in[21] ));
 sg13g2_inv_1 _4760_ (.Y(_3982_),
    .A(\debug_controller_inst.grid_in[53] ));
 sg13g2_inv_1 _4761_ (.Y(_3983_),
    .A(\debug_controller_inst.grid_in[22] ));
 sg13g2_inv_1 _4762_ (.Y(_3984_),
    .A(\debug_controller_inst.grid_in[54] ));
 sg13g2_inv_1 _4763_ (.Y(_3985_),
    .A(\debug_controller_inst.grid_in[23] ));
 sg13g2_inv_1 _4764_ (.Y(_3986_),
    .A(\debug_controller_inst.grid_in[55] ));
 sg13g2_inv_1 _4765_ (.Y(_3987_),
    .A(_0069_));
 sg13g2_inv_1 _4766_ (.Y(_3988_),
    .A(\btn_up_debounce.debounce_counter[13] ));
 sg13g2_inv_1 _4767_ (.Y(_3989_),
    .A(\btn_right_debounce.debounce_counter[13] ));
 sg13g2_inv_1 _4768_ (.Y(_3990_),
    .A(\btn_left_debounce.debounce_counter[14] ));
 sg13g2_inv_1 _4769_ (.Y(_3991_),
    .A(\btn_down_debounce.debounce_counter[7] ));
 sg13g2_inv_2 _4770_ (.Y(_3992_),
    .A(net896));
 sg13g2_inv_2 _4771_ (.Y(_3993_),
    .A(net2154));
 sg13g2_inv_1 _4772_ (.Y(_3994_),
    .A(net2155));
 sg13g2_inv_2 _4773_ (.Y(_3995_),
    .A(net2162));
 sg13g2_inv_1 _4774_ (.Y(_3996_),
    .A(net2175));
 sg13g2_inv_2 _4775_ (.Y(_3997_),
    .A(net2193));
 sg13g2_inv_2 _4776_ (.Y(_3998_),
    .A(net2220));
 sg13g2_inv_2 _4777_ (.Y(_3999_),
    .A(net2147));
 sg13g2_inv_1 _4778_ (.Y(_4000_),
    .A(net829));
 sg13g2_inv_1 _4779_ (.Y(_4001_),
    .A(net2136));
 sg13g2_inv_1 _4780_ (.Y(_4002_),
    .A(net2144));
 sg13g2_inv_2 _4781_ (.Y(_4003_),
    .A(net2100));
 sg13g2_inv_1 _4782_ (.Y(_4004_),
    .A(\new_tiles_counter[0] ));
 sg13g2_inv_1 _4783_ (.Y(_4005_),
    .A(\draw_game_inst.new_tiles_counter[2] ));
 sg13g2_inv_1 _4784_ (.Y(_4006_),
    .A(net689));
 sg13g2_inv_1 _4785_ (.Y(_4007_),
    .A(net499));
 sg13g2_inv_1 _4786_ (.Y(_4008_),
    .A(net843));
 sg13g2_inv_1 _4787_ (.Y(_4009_),
    .A(_0099_));
 sg13g2_inv_1 _4788_ (.Y(_4010_),
    .A(\debug_controller_inst.grid_out_valid ));
 sg13g2_inv_1 _4789_ (.Y(_4011_),
    .A(net928));
 sg13g2_inv_1 _4790_ (.Y(_4012_),
    .A(net905));
 sg13g2_inv_1 _4791_ (.Y(_4013_),
    .A(_0105_));
 sg13g2_inv_1 _4792_ (.Y(_4014_),
    .A(net981));
 sg13g2_inv_1 _4793_ (.Y(_4015_),
    .A(net900));
 sg13g2_inv_1 _4794_ (.Y(_4016_),
    .A(net1000));
 sg13g2_inv_1 _4795_ (.Y(_4017_),
    .A(net924));
 sg13g2_inv_1 _4796_ (.Y(_4018_),
    .A(net997));
 sg13g2_inv_1 _4797_ (.Y(_4019_),
    .A(net989));
 sg13g2_inv_1 _4798_ (.Y(_4020_),
    .A(net919));
 sg13g2_inv_1 _4799_ (.Y(_4021_),
    .A(net1023));
 sg13g2_inv_1 _4800_ (.Y(_4022_),
    .A(_0115_));
 sg13g2_inv_1 _4801_ (.Y(_4023_),
    .A(net1017));
 sg13g2_inv_1 _4802_ (.Y(_4024_),
    .A(net942));
 sg13g2_inv_1 _4803_ (.Y(_4025_),
    .A(net1020));
 sg13g2_inv_1 _4804_ (.Y(_4026_),
    .A(net1028));
 sg13g2_inv_1 _4805_ (.Y(_4027_),
    .A(net1035));
 sg13g2_inv_1 _4806_ (.Y(_4028_),
    .A(net1027));
 sg13g2_inv_1 _4807_ (.Y(_4029_),
    .A(net891));
 sg13g2_inv_1 _4808_ (.Y(_4030_),
    .A(_0127_));
 sg13g2_inv_1 _4809_ (.Y(_4031_),
    .A(net1001));
 sg13g2_inv_1 _4810_ (.Y(_0496_),
    .A(net1033));
 sg13g2_inv_1 _4811_ (.Y(_0497_),
    .A(net1019));
 sg13g2_inv_1 _4812_ (.Y(_0498_),
    .A(net1029));
 sg13g2_inv_1 _4813_ (.Y(_0499_),
    .A(net965));
 sg13g2_inv_1 _4814_ (.Y(_0500_),
    .A(_0151_));
 sg13g2_inv_1 _4815_ (.Y(_0501_),
    .A(_0155_));
 sg13g2_inv_1 _4816_ (.Y(_0502_),
    .A(net1036));
 sg13g2_inv_1 _4817_ (.Y(_0503_),
    .A(net1039));
 sg13g2_inv_1 _4818_ (.Y(_0504_),
    .A(net419));
 sg13g2_inv_1 _4819_ (.Y(_0505_),
    .A(net420));
 sg13g2_nand4_1 _4820_ (.B(\gamepad_pmod.decoder.data_reg[8] ),
    .C(\gamepad_pmod.decoder.data_reg[11] ),
    .A(\gamepad_pmod.decoder.data_reg[9] ),
    .Y(_0506_),
    .D(\gamepad_pmod.decoder.data_reg[10] ));
 sg13g2_nand4_1 _4821_ (.B(\gamepad_pmod.decoder.data_reg[4] ),
    .C(\gamepad_pmod.decoder.data_reg[7] ),
    .A(\gamepad_pmod.decoder.data_reg[5] ),
    .Y(_0507_),
    .D(\gamepad_pmod.decoder.data_reg[6] ));
 sg13g2_nand4_1 _4822_ (.B(\gamepad_pmod.decoder.data_reg[0] ),
    .C(\gamepad_pmod.decoder.data_reg[3] ),
    .A(\gamepad_pmod.decoder.data_reg[1] ),
    .Y(_0508_),
    .D(\gamepad_pmod.decoder.data_reg[2] ));
 sg13g2_or3_2 _4823_ (.A(_0506_),
    .B(_0507_),
    .C(_0508_),
    .X(_0509_));
 sg13g2_a21o_2 _4824_ (.A2(_0509_),
    .A1(net1034),
    .B1(\btn_down_debounce.debounced ),
    .X(_0510_));
 sg13g2_a21oi_1 _4825_ (.A1(net1002),
    .A2(_0510_),
    .Y(_0511_),
    .B1(debug_btn_down));
 sg13g2_a21o_2 _4826_ (.A2(_0509_),
    .A1(\gamepad_pmod.decoder.data_reg[7] ),
    .B1(\btn_up_debounce.debounced ),
    .X(_0512_));
 sg13g2_a21oi_2 _4827_ (.B1(debug_btn_up),
    .Y(_0513_),
    .A2(_0512_),
    .A1(net1002));
 sg13g2_a21o_2 _4828_ (.A2(_0509_),
    .A1(\gamepad_pmod.decoder.data_reg[5] ),
    .B1(\btn_left_debounce.debounced ),
    .X(_0514_));
 sg13g2_a21oi_1 _4829_ (.A1(_0165_),
    .A2(_0514_),
    .Y(_0515_),
    .B1(debug_btn_left));
 sg13g2_a21o_2 _4830_ (.A2(_0509_),
    .A1(\gamepad_pmod.decoder.data_reg[4] ),
    .B1(net685),
    .X(_0516_));
 sg13g2_a21oi_1 _4831_ (.A1(_0165_),
    .A2(_0516_),
    .Y(_0517_),
    .B1(debug_btn_right));
 sg13g2_a21o_1 _4832_ (.A2(_0516_),
    .A1(net1002),
    .B1(debug_btn_right),
    .X(_0518_));
 sg13g2_nand4_1 _4833_ (.B(_0513_),
    .C(_0515_),
    .A(_0511_),
    .Y(_0519_),
    .D(_0517_));
 sg13g2_nor2b_1 _4834_ (.A(\game_logic_inst.prev_any_button_pressed ),
    .B_N(_0519_),
    .Y(_0520_));
 sg13g2_nand2b_2 _4835_ (.Y(_0521_),
    .B(_0519_),
    .A_N(\game_logic_inst.prev_any_button_pressed ));
 sg13g2_o21ai_1 _4836_ (.B1(net2107),
    .Y(_0522_),
    .A1(net915),
    .A2(net1777));
 sg13g2_and2_1 _4837_ (.A(net2268),
    .B(_0522_),
    .X(_0523_));
 sg13g2_nor2_2 _4838_ (.A(net2257),
    .B(net915),
    .Y(_0524_));
 sg13g2_nand3_1 _4839_ (.B(net1777),
    .C(_0524_),
    .A(_0515_),
    .Y(_0525_));
 sg13g2_nor3_1 _4840_ (.A(_0511_),
    .B(_0518_),
    .C(_0525_),
    .Y(_0526_));
 sg13g2_a22oi_1 _4841_ (.Y(_0527_),
    .B1(_0526_),
    .B2(net1003),
    .A2(_0523_),
    .A1(\game_logic_inst.current_direction[3] ));
 sg13g2_inv_1 _4842_ (.Y(_0002_),
    .A(net1004));
 sg13g2_nand2_1 _4843_ (.Y(_0528_),
    .A(net955),
    .B(_0523_));
 sg13g2_o21ai_1 _4844_ (.B1(_0528_),
    .Y(_0001_),
    .A1(_0517_),
    .A2(_0525_));
 sg13g2_nor3_1 _4845_ (.A(_0513_),
    .B(_0518_),
    .C(_0525_),
    .Y(_0529_));
 sg13g2_a21o_1 _4846_ (.A2(_0523_),
    .A1(net634),
    .B1(_0529_),
    .X(_0000_));
 sg13g2_nor2_1 _4847_ (.A(\debug_controller_inst.grid_out_addr[1] ),
    .B(\debug_controller_inst.grid_out_addr[0] ),
    .Y(_0530_));
 sg13g2_nor3_2 _4848_ (.A(net2084),
    .B(\debug_controller_inst.grid_out_addr[1] ),
    .C(\debug_controller_inst.grid_out_addr[0] ),
    .Y(_0531_));
 sg13g2_nand2b_2 _4849_ (.Y(_0532_),
    .B(_0531_),
    .A_N(\debug_controller_inst.grid_out_addr[3] ));
 sg13g2_nor2_2 _4850_ (.A(_4010_),
    .B(_0532_),
    .Y(_0533_));
 sg13g2_nand2_1 _4851_ (.Y(_0534_),
    .A(net2093),
    .B(_0533_));
 sg13g2_nor2_1 _4852_ (.A(net2096),
    .B(net2099),
    .Y(_0535_));
 sg13g2_or2_1 _4853_ (.X(_0536_),
    .B(net2099),
    .A(net2096));
 sg13g2_nor2_1 _4854_ (.A(\game_logic_inst.current_direction[3] ),
    .B(\game_logic_inst.current_direction[2] ),
    .Y(_0537_));
 sg13g2_or2_1 _4855_ (.X(_0538_),
    .B(\game_logic_inst.current_direction[2] ),
    .A(\game_logic_inst.current_direction[3] ));
 sg13g2_nor2b_1 _4856_ (.A(net2096),
    .B_N(net2099),
    .Y(_0539_));
 sg13g2_nor2b_2 _4857_ (.A(net2098),
    .B_N(net2095),
    .Y(_0540_));
 sg13g2_nand2b_1 _4858_ (.Y(_0541_),
    .B(\game_logic_inst.current_row_index[1] ),
    .A_N(\game_logic_inst.current_row_index[0] ));
 sg13g2_and2_1 _4859_ (.A(net2096),
    .B(net2099),
    .X(_0542_));
 sg13g2_nand2_1 _4860_ (.Y(_0543_),
    .A(net2096),
    .B(net2099));
 sg13g2_mux4_1 _4861_ (.S0(net2098),
    .A0(\debug_controller_inst.grid_in[0] ),
    .A1(\debug_controller_inst.grid_in[16] ),
    .A2(\debug_controller_inst.grid_in[32] ),
    .A3(\debug_controller_inst.grid_in[48] ),
    .S1(net2095),
    .X(_0544_));
 sg13g2_mux4_1 _4862_ (.S0(net2097),
    .A0(\debug_controller_inst.grid_in[12] ),
    .A1(\debug_controller_inst.grid_in[28] ),
    .A2(\debug_controller_inst.grid_in[44] ),
    .A3(\debug_controller_inst.grid_in[60] ),
    .S1(net2094),
    .X(_0545_));
 sg13g2_mux2_2 _4863_ (.A0(_0544_),
    .A1(_0545_),
    .S(net2014),
    .X(_0546_));
 sg13g2_mux4_1 _4864_ (.S0(net2097),
    .A0(\debug_controller_inst.grid_in[5] ),
    .A1(\debug_controller_inst.grid_in[21] ),
    .A2(\debug_controller_inst.grid_in[37] ),
    .A3(\debug_controller_inst.grid_in[53] ),
    .S1(net2094),
    .X(_0547_));
 sg13g2_nand2_1 _4865_ (.Y(_0548_),
    .A(net2009),
    .B(_0547_));
 sg13g2_mux4_1 _4866_ (.S0(net2098),
    .A0(\debug_controller_inst.grid_in[9] ),
    .A1(\debug_controller_inst.grid_in[25] ),
    .A2(\debug_controller_inst.grid_in[41] ),
    .A3(\debug_controller_inst.grid_in[57] ),
    .S1(net2095),
    .X(_0549_));
 sg13g2_nand2_1 _4867_ (.Y(_0550_),
    .A(net2014),
    .B(_0549_));
 sg13g2_nand2_2 _4868_ (.Y(_0551_),
    .A(_0548_),
    .B(_0550_));
 sg13g2_mux4_1 _4869_ (.S0(net2097),
    .A0(\debug_controller_inst.grid_in[7] ),
    .A1(\debug_controller_inst.grid_in[23] ),
    .A2(\debug_controller_inst.grid_in[39] ),
    .A3(\debug_controller_inst.grid_in[55] ),
    .S1(net2094),
    .X(_0552_));
 sg13g2_mux4_1 _4870_ (.S0(net2097),
    .A0(\debug_controller_inst.grid_in[11] ),
    .A1(\debug_controller_inst.grid_in[27] ),
    .A2(\debug_controller_inst.grid_in[43] ),
    .A3(\debug_controller_inst.grid_in[59] ),
    .S1(net2094),
    .X(_0553_));
 sg13g2_mux2_2 _4871_ (.A0(_0552_),
    .A1(_0553_),
    .S(net2014),
    .X(_0554_));
 sg13g2_mux4_1 _4872_ (.S0(net2097),
    .A0(\debug_controller_inst.grid_in[6] ),
    .A1(\debug_controller_inst.grid_in[22] ),
    .A2(\debug_controller_inst.grid_in[38] ),
    .A3(\debug_controller_inst.grid_in[54] ),
    .S1(net2094),
    .X(_0555_));
 sg13g2_nand2_1 _4873_ (.Y(_0556_),
    .A(net2011),
    .B(_0555_));
 sg13g2_mux4_1 _4874_ (.S0(net2098),
    .A0(\debug_controller_inst.grid_in[10] ),
    .A1(\debug_controller_inst.grid_in[26] ),
    .A2(\debug_controller_inst.grid_in[42] ),
    .A3(\debug_controller_inst.grid_in[58] ),
    .S1(net2095),
    .X(_0557_));
 sg13g2_nand2_1 _4875_ (.Y(_0558_),
    .A(net2014),
    .B(_0557_));
 sg13g2_nand2_2 _4876_ (.Y(_0559_),
    .A(_0556_),
    .B(_0558_));
 sg13g2_mux4_1 _4877_ (.S0(net2099),
    .A0(\debug_controller_inst.grid_in[4] ),
    .A1(\debug_controller_inst.grid_in[20] ),
    .A2(\debug_controller_inst.grid_in[36] ),
    .A3(\debug_controller_inst.grid_in[52] ),
    .S1(net2096),
    .X(_0560_));
 sg13g2_inv_1 _4878_ (.Y(_0561_),
    .A(_0560_));
 sg13g2_mux4_1 _4879_ (.S0(net2098),
    .A0(\debug_controller_inst.grid_in[8] ),
    .A1(\debug_controller_inst.grid_in[24] ),
    .A2(\debug_controller_inst.grid_in[40] ),
    .A3(\debug_controller_inst.grid_in[56] ),
    .S1(net2095),
    .X(_0562_));
 sg13g2_nand2_1 _4880_ (.Y(_0563_),
    .A(net2014),
    .B(_0562_));
 sg13g2_o21ai_1 _4881_ (.B1(_0563_),
    .Y(_0564_),
    .A1(net2013),
    .A2(_0561_));
 sg13g2_inv_2 _4882_ (.Y(_0565_),
    .A(_0564_));
 sg13g2_nor4_2 _4883_ (.A(_0551_),
    .B(_0554_),
    .C(_0559_),
    .Y(_0566_),
    .D(_0564_));
 sg13g2_inv_2 _4884_ (.Y(_0567_),
    .A(_0566_));
 sg13g2_mux2_2 _4885_ (.A0(_0555_),
    .A1(_0557_),
    .S(net2009),
    .X(_0568_));
 sg13g2_mux2_2 _4886_ (.A0(_0552_),
    .A1(_0553_),
    .S(net2009),
    .X(_0569_));
 sg13g2_mux2_2 _4887_ (.A0(_0560_),
    .A1(_0562_),
    .S(net2009),
    .X(_0570_));
 sg13g2_mux2_2 _4888_ (.A0(_0547_),
    .A1(_0549_),
    .S(net2009),
    .X(_0571_));
 sg13g2_nor4_2 _4889_ (.A(_0568_),
    .B(_0569_),
    .C(_0570_),
    .Y(_0572_),
    .D(_0571_));
 sg13g2_mux4_1 _4890_ (.S0(net2097),
    .A0(\debug_controller_inst.grid_in[13] ),
    .A1(\debug_controller_inst.grid_in[29] ),
    .A2(\debug_controller_inst.grid_in[45] ),
    .A3(\debug_controller_inst.grid_in[61] ),
    .S1(net2094),
    .X(_0573_));
 sg13g2_mux4_1 _4891_ (.S0(net2098),
    .A0(\debug_controller_inst.grid_in[1] ),
    .A1(\debug_controller_inst.grid_in[17] ),
    .A2(\debug_controller_inst.grid_in[33] ),
    .A3(\debug_controller_inst.grid_in[49] ),
    .S1(net2095),
    .X(_0574_));
 sg13g2_mux2_2 _4892_ (.A0(_0573_),
    .A1(_0574_),
    .S(net2013),
    .X(_0575_));
 sg13g2_mux4_1 _4893_ (.S0(net2098),
    .A0(\debug_controller_inst.grid_in[2] ),
    .A1(\debug_controller_inst.grid_in[18] ),
    .A2(\debug_controller_inst.grid_in[34] ),
    .A3(\debug_controller_inst.grid_in[50] ),
    .S1(net2095),
    .X(_0576_));
 sg13g2_mux4_1 _4894_ (.S0(net2097),
    .A0(\debug_controller_inst.grid_in[14] ),
    .A1(\debug_controller_inst.grid_in[30] ),
    .A2(\debug_controller_inst.grid_in[46] ),
    .A3(\debug_controller_inst.grid_in[62] ),
    .S1(net2094),
    .X(_0577_));
 sg13g2_mux2_2 _4895_ (.A0(_0576_),
    .A1(_0577_),
    .S(net2009),
    .X(_0578_));
 sg13g2_mux2_2 _4896_ (.A0(_0544_),
    .A1(_0545_),
    .S(net2009),
    .X(_0579_));
 sg13g2_mux4_1 _4897_ (.S0(net2098),
    .A0(\debug_controller_inst.grid_in[3] ),
    .A1(\debug_controller_inst.grid_in[19] ),
    .A2(\debug_controller_inst.grid_in[35] ),
    .A3(\debug_controller_inst.grid_in[51] ),
    .S1(net2095),
    .X(_0580_));
 sg13g2_mux4_1 _4898_ (.S0(net2097),
    .A0(\debug_controller_inst.grid_in[15] ),
    .A1(\debug_controller_inst.grid_in[31] ),
    .A2(\debug_controller_inst.grid_in[47] ),
    .A3(\debug_controller_inst.grid_in[63] ),
    .S1(net2094),
    .X(_0581_));
 sg13g2_mux2_2 _4899_ (.A0(_0580_),
    .A1(_0581_),
    .S(net2009),
    .X(_0582_));
 sg13g2_nor4_2 _4900_ (.A(_0575_),
    .B(_0578_),
    .C(_0579_),
    .Y(_0583_),
    .D(_0582_));
 sg13g2_or4_2 _4901_ (.A(_0575_),
    .B(_0578_),
    .C(_0579_),
    .D(_0582_),
    .X(_0584_));
 sg13g2_and2_2 _4902_ (.A(_0572_),
    .B(_0583_),
    .X(_0585_));
 sg13g2_xnor2_1 _4903_ (.Y(_0586_),
    .A(_0569_),
    .B(_0582_));
 sg13g2_xnor2_1 _4904_ (.Y(_0587_),
    .A(_0570_),
    .B(_0579_));
 sg13g2_xnor2_1 _4905_ (.Y(_0588_),
    .A(_0568_),
    .B(_0578_));
 sg13g2_xnor2_1 _4906_ (.Y(_0589_),
    .A(_0571_),
    .B(_0575_));
 sg13g2_and4_2 _4907_ (.A(_0586_),
    .B(_0587_),
    .C(_0588_),
    .D(_0589_),
    .X(_0590_));
 sg13g2_nand4_1 _4908_ (.B(_0587_),
    .C(_0588_),
    .A(_0586_),
    .Y(_0591_),
    .D(_0589_));
 sg13g2_nand3_1 _4909_ (.B(_0584_),
    .C(_0591_),
    .A(_0568_),
    .Y(_0592_));
 sg13g2_xor2_1 _4910_ (.B(_0592_),
    .A(_0559_),
    .X(_0593_));
 sg13g2_nand3_1 _4911_ (.B(_0584_),
    .C(net1791),
    .A(_0570_),
    .Y(_0594_));
 sg13g2_xnor2_1 _4912_ (.Y(_0595_),
    .A(_0565_),
    .B(_0594_));
 sg13g2_nand3_1 _4913_ (.B(_0584_),
    .C(net1791),
    .A(_0569_),
    .Y(_0596_));
 sg13g2_xor2_1 _4914_ (.B(_0596_),
    .A(_0554_),
    .X(_0597_));
 sg13g2_nand3_1 _4915_ (.B(_0584_),
    .C(net1791),
    .A(_0571_),
    .Y(_0598_));
 sg13g2_xor2_1 _4916_ (.B(_0598_),
    .A(_0551_),
    .X(_0599_));
 sg13g2_nand4_1 _4917_ (.B(_0595_),
    .C(_0597_),
    .A(_0593_),
    .Y(_0600_),
    .D(_0599_));
 sg13g2_and2_1 _4918_ (.A(_0575_),
    .B(_0579_),
    .X(_0601_));
 sg13g2_and2_1 _4919_ (.A(_0590_),
    .B(_0601_),
    .X(_0602_));
 sg13g2_a21oi_1 _4920_ (.A1(_0590_),
    .A2(_0601_),
    .Y(_0603_),
    .B1(_0578_));
 sg13g2_nand2_1 _4921_ (.Y(_0604_),
    .A(_0578_),
    .B(_0601_));
 sg13g2_o21ai_1 _4922_ (.B1(_0584_),
    .Y(_0605_),
    .A1(net1791),
    .A2(_0604_));
 sg13g2_nand2_1 _4923_ (.Y(_0606_),
    .A(_0568_),
    .B(_0583_));
 sg13g2_o21ai_1 _4924_ (.B1(_0606_),
    .Y(_0607_),
    .A1(_0603_),
    .A2(_0605_));
 sg13g2_xnor2_1 _4925_ (.Y(_0608_),
    .A(_0559_),
    .B(_0607_));
 sg13g2_nand2b_1 _4926_ (.Y(_0609_),
    .B(net1791),
    .A_N(_0579_));
 sg13g2_a21oi_1 _4927_ (.A1(_0579_),
    .A2(_0590_),
    .Y(_0610_),
    .B1(_0583_));
 sg13g2_a22oi_1 _4928_ (.Y(_0611_),
    .B1(_0609_),
    .B2(_0610_),
    .A2(_0583_),
    .A1(_0570_));
 sg13g2_xnor2_1 _4929_ (.Y(_0612_),
    .A(_0565_),
    .B(_0611_));
 sg13g2_nand2_1 _4930_ (.Y(_0613_),
    .A(_0569_),
    .B(_0583_));
 sg13g2_o21ai_1 _4931_ (.B1(_0582_),
    .Y(_0614_),
    .A1(net1791),
    .A2(_0604_));
 sg13g2_or3_1 _4932_ (.A(_0582_),
    .B(net1791),
    .C(_0604_),
    .X(_0615_));
 sg13g2_nand3_1 _4933_ (.B(_0614_),
    .C(_0615_),
    .A(_0613_),
    .Y(_0616_));
 sg13g2_xnor2_1 _4934_ (.Y(_0617_),
    .A(_0554_),
    .B(_0616_));
 sg13g2_nand2_1 _4935_ (.Y(_0618_),
    .A(_0571_),
    .B(_0583_));
 sg13g2_a21oi_1 _4936_ (.A1(_0579_),
    .A2(_0590_),
    .Y(_0619_),
    .B1(_0575_));
 sg13g2_o21ai_1 _4937_ (.B1(_0618_),
    .Y(_0620_),
    .A1(_0602_),
    .A2(_0619_));
 sg13g2_xnor2_1 _4938_ (.Y(_0621_),
    .A(_0551_),
    .B(_0620_));
 sg13g2_and4_1 _4939_ (.A(_0608_),
    .B(_0612_),
    .C(_0617_),
    .D(_0621_),
    .X(_0622_));
 sg13g2_nand4_1 _4940_ (.B(_0612_),
    .C(_0617_),
    .A(_0608_),
    .Y(_0623_),
    .D(_0621_));
 sg13g2_nor2_2 _4941_ (.A(_0572_),
    .B(_0591_),
    .Y(_0624_));
 sg13g2_nand2b_1 _4942_ (.Y(_0625_),
    .B(_0590_),
    .A_N(_0572_));
 sg13g2_nor3_2 _4943_ (.A(_0572_),
    .B(_0583_),
    .C(_0590_),
    .Y(_0626_));
 sg13g2_inv_1 _4944_ (.Y(_0627_),
    .A(net1783));
 sg13g2_or2_1 _4945_ (.X(_0628_),
    .B(_0626_),
    .A(_0585_));
 sg13g2_a21o_1 _4946_ (.A2(_0625_),
    .A1(_0622_),
    .B1(_0628_),
    .X(_0629_));
 sg13g2_a21oi_2 _4947_ (.B1(_0585_),
    .Y(_0630_),
    .A2(_0629_),
    .A1(_0600_));
 sg13g2_nand2_1 _4948_ (.Y(_0631_),
    .A(_0567_),
    .B(_0630_));
 sg13g2_xnor2_1 _4949_ (.Y(_0632_),
    .A(_0566_),
    .B(_0630_));
 sg13g2_xnor2_1 _4950_ (.Y(_0633_),
    .A(_0567_),
    .B(_0630_));
 sg13g2_nand2b_1 _4951_ (.Y(_0634_),
    .B(_0567_),
    .A_N(_0600_));
 sg13g2_nand2_2 _4952_ (.Y(_0635_),
    .A(net1764),
    .B(net1783));
 sg13g2_nand2_1 _4953_ (.Y(_0636_),
    .A(_0631_),
    .B(_0635_));
 sg13g2_nor2_2 _4954_ (.A(_0633_),
    .B(_0635_),
    .Y(_0637_));
 sg13g2_mux2_2 _4955_ (.A0(_0580_),
    .A1(_0581_),
    .S(net2012),
    .X(_0638_));
 sg13g2_nor2b_1 _4956_ (.A(_0635_),
    .B_N(_0554_),
    .Y(_0639_));
 sg13g2_nand3_1 _4957_ (.B(net1764),
    .C(net1783),
    .A(_0554_),
    .Y(_0640_));
 sg13g2_xnor2_1 _4958_ (.Y(_0641_),
    .A(_0638_),
    .B(_0640_));
 sg13g2_nand3_1 _4959_ (.B(net1764),
    .C(net1783),
    .A(_0564_),
    .Y(_0642_));
 sg13g2_xnor2_1 _4960_ (.Y(_0643_),
    .A(_0546_),
    .B(_0642_));
 sg13g2_and2_1 _4961_ (.A(net2010),
    .B(_0576_),
    .X(_0644_));
 sg13g2_and2_1 _4962_ (.A(net2013),
    .B(_0577_),
    .X(_0645_));
 sg13g2_nor2_1 _4963_ (.A(_0644_),
    .B(_0645_),
    .Y(_0646_));
 sg13g2_or2_2 _4964_ (.X(_0647_),
    .B(_0645_),
    .A(_0644_));
 sg13g2_nor2b_1 _4965_ (.A(_0635_),
    .B_N(_0559_),
    .Y(_0648_));
 sg13g2_nand3_1 _4966_ (.B(net1764),
    .C(net1783),
    .A(_0559_),
    .Y(_0649_));
 sg13g2_xnor2_1 _4967_ (.Y(_0650_),
    .A(_0647_),
    .B(_0649_));
 sg13g2_and2_1 _4968_ (.A(net2010),
    .B(_0574_),
    .X(_0651_));
 sg13g2_a21oi_2 _4969_ (.B1(_0651_),
    .Y(_0652_),
    .A2(_0573_),
    .A1(net2012));
 sg13g2_inv_2 _4970_ (.Y(_0653_),
    .A(_0652_));
 sg13g2_nor2b_1 _4971_ (.A(_0635_),
    .B_N(_0551_),
    .Y(_0654_));
 sg13g2_nand3_1 _4972_ (.B(net1764),
    .C(net1783),
    .A(_0551_),
    .Y(_0655_));
 sg13g2_xnor2_1 _4973_ (.Y(_0656_),
    .A(_0653_),
    .B(_0655_));
 sg13g2_nor4_2 _4974_ (.A(_0641_),
    .B(_0643_),
    .C(_0650_),
    .Y(_0657_),
    .D(_0656_));
 sg13g2_nor3_2 _4975_ (.A(_0633_),
    .B(_0635_),
    .C(_0657_),
    .Y(_0658_));
 sg13g2_and2_1 _4976_ (.A(net1919),
    .B(_0658_),
    .X(_0659_));
 sg13g2_nand2_1 _4977_ (.Y(_0660_),
    .A(_0564_),
    .B(_0585_));
 sg13g2_nor4_2 _4978_ (.A(_0565_),
    .B(_0623_),
    .C(_0624_),
    .Y(_0661_),
    .D(_0626_));
 sg13g2_nand4_1 _4979_ (.B(_0622_),
    .C(_0625_),
    .A(_0567_),
    .Y(_0662_),
    .D(_0627_));
 sg13g2_a21o_1 _4980_ (.A2(_0662_),
    .A1(_0611_),
    .B1(_0661_),
    .X(_0663_));
 sg13g2_and2_1 _4981_ (.A(_0660_),
    .B(_0663_),
    .X(_0664_));
 sg13g2_nand2_1 _4982_ (.Y(_0665_),
    .A(_0660_),
    .B(_0663_));
 sg13g2_nand2_1 _4983_ (.Y(_0666_),
    .A(_0559_),
    .B(_0585_));
 sg13g2_nand2b_1 _4984_ (.Y(_0667_),
    .B(_0620_),
    .A_N(_0611_));
 sg13g2_nor4_2 _4985_ (.A(_0623_),
    .B(_0624_),
    .C(net1783),
    .Y(_0668_),
    .D(_0667_));
 sg13g2_xnor2_1 _4986_ (.Y(_0669_),
    .A(_0607_),
    .B(_0668_));
 sg13g2_nand2_1 _4987_ (.Y(_0670_),
    .A(_0666_),
    .B(_0669_));
 sg13g2_inv_1 _4988_ (.Y(_0671_),
    .A(_0670_));
 sg13g2_and3_1 _4989_ (.X(_0672_),
    .A(_0647_),
    .B(_0666_),
    .C(_0669_));
 sg13g2_a21oi_1 _4990_ (.A1(_0666_),
    .A2(_0669_),
    .Y(_0673_),
    .B1(_0647_));
 sg13g2_a21oi_1 _4991_ (.A1(net1791),
    .A2(_0623_),
    .Y(_0674_),
    .B1(_0628_));
 sg13g2_a21o_1 _4992_ (.A2(_0668_),
    .A1(_0607_),
    .B1(_0616_),
    .X(_0675_));
 sg13g2_nand3_1 _4993_ (.B(_0616_),
    .C(_0668_),
    .A(_0607_),
    .Y(_0676_));
 sg13g2_a22oi_1 _4994_ (.Y(_0677_),
    .B1(_0675_),
    .B2(_0676_),
    .A2(_0585_),
    .A1(_0554_));
 sg13g2_nand2_1 _4995_ (.Y(_0678_),
    .A(_0551_),
    .B(_0585_));
 sg13g2_inv_1 _4996_ (.Y(_0679_),
    .A(_0678_));
 sg13g2_xor2_1 _4997_ (.B(_0661_),
    .A(_0620_),
    .X(_0680_));
 sg13g2_nor2_2 _4998_ (.A(_0679_),
    .B(_0680_),
    .Y(_0681_));
 sg13g2_o21ai_1 _4999_ (.B1(_0653_),
    .Y(_0682_),
    .A1(_0679_),
    .A2(_0680_));
 sg13g2_nand3b_1 _5000_ (.B(_0652_),
    .C(_0678_),
    .Y(_0683_),
    .A_N(_0680_));
 sg13g2_a221oi_1 _5001_ (.B2(_0683_),
    .C1(_0674_),
    .B1(_0682_),
    .A1(net1919),
    .Y(_0684_),
    .A2(_0664_));
 sg13g2_xor2_1 _5002_ (.B(_0677_),
    .A(net1918),
    .X(_0685_));
 sg13g2_a21oi_1 _5003_ (.A1(_0660_),
    .A2(_0663_),
    .Y(_0686_),
    .B1(net1919));
 sg13g2_nor3_2 _5004_ (.A(_0672_),
    .B(_0673_),
    .C(_0686_),
    .Y(_0687_));
 sg13g2_and3_1 _5005_ (.X(_0688_),
    .A(_0684_),
    .B(_0685_),
    .C(_0687_));
 sg13g2_nand4_1 _5006_ (.B(_0684_),
    .C(_0685_),
    .A(_0665_),
    .Y(_0689_),
    .D(_0687_));
 sg13g2_and2_2 _5007_ (.A(_0632_),
    .B(_0635_),
    .X(_0690_));
 sg13g2_inv_1 _5008_ (.Y(_0691_),
    .A(_0690_));
 sg13g2_xnor2_1 _5009_ (.Y(_0692_),
    .A(_0665_),
    .B(_0688_));
 sg13g2_or4_2 _5010_ (.A(net1919),
    .B(_0638_),
    .C(_0647_),
    .D(_0653_),
    .X(_0693_));
 sg13g2_inv_1 _5011_ (.Y(_0694_),
    .A(_0693_));
 sg13g2_nand3_1 _5012_ (.B(_0635_),
    .C(_0693_),
    .A(_0631_),
    .Y(_0695_));
 sg13g2_inv_1 _5013_ (.Y(_0696_),
    .A(_0695_));
 sg13g2_nor3_2 _5014_ (.A(_0567_),
    .B(net1783),
    .C(_0630_),
    .Y(_0697_));
 sg13g2_a21oi_1 _5015_ (.A1(net1919),
    .A2(_0697_),
    .Y(_0698_),
    .B1(_0695_));
 sg13g2_o21ai_1 _5016_ (.B1(_0698_),
    .Y(_0699_),
    .A1(_0691_),
    .A2(_0692_));
 sg13g2_o21ai_1 _5017_ (.B1(_0699_),
    .Y(_0700_),
    .A1(_0665_),
    .A2(_0696_));
 sg13g2_nor2_1 _5018_ (.A(net2012),
    .B(_0659_),
    .Y(_0701_));
 sg13g2_a21oi_2 _5019_ (.B1(_0701_),
    .Y(_0702_),
    .A2(_0700_),
    .A1(net2012));
 sg13g2_o21ai_1 _5020_ (.B1(net2121),
    .Y(_0703_),
    .A1(_0099_),
    .A2(_0535_));
 sg13g2_a21oi_1 _5021_ (.A1(_0535_),
    .A2(_0702_),
    .Y(_0704_),
    .B1(_0703_));
 sg13g2_nor2_1 _5022_ (.A(\game_logic_inst.should_transpose ),
    .B(net1776),
    .Y(_0705_));
 sg13g2_nand2_1 _5023_ (.Y(_0706_),
    .A(_3938_),
    .B(net1775));
 sg13g2_mux4_1 _5024_ (.S0(\game_logic_inst.lfsr_shift[0] ),
    .A0(\game_logic_inst.lfsr_value[3] ),
    .A1(\game_logic_inst.lfsr_value[7] ),
    .A2(\game_logic_inst.lfsr_value[11] ),
    .A3(\game_logic_inst.lfsr_value[15] ),
    .S1(\game_logic_inst.lfsr_shift[1] ),
    .X(_0707_));
 sg13g2_inv_2 _5025_ (.Y(_0708_),
    .A(_0707_));
 sg13g2_mux2_1 _5026_ (.A0(\game_logic_inst.lfsr_value[2] ),
    .A1(\game_logic_inst.lfsr_value[6] ),
    .S(\game_logic_inst.lfsr_shift[0] ),
    .X(_0709_));
 sg13g2_nor2_1 _5027_ (.A(\game_logic_inst.lfsr_shift[1] ),
    .B(_0709_),
    .Y(_0710_));
 sg13g2_nand2_1 _5028_ (.Y(_0711_),
    .A(\game_logic_inst.lfsr_shift[0] ),
    .B(\game_logic_inst.lfsr_value[14] ));
 sg13g2_nand2b_1 _5029_ (.Y(_0712_),
    .B(\game_logic_inst.lfsr_value[10] ),
    .A_N(\game_logic_inst.lfsr_shift[0] ));
 sg13g2_nand3_1 _5030_ (.B(_0711_),
    .C(_0712_),
    .A(\game_logic_inst.lfsr_shift[1] ),
    .Y(_0713_));
 sg13g2_nand2b_2 _5031_ (.Y(_0714_),
    .B(_0713_),
    .A_N(_0710_));
 sg13g2_nor2b_2 _5032_ (.A(_0710_),
    .B_N(_0713_),
    .Y(_0715_));
 sg13g2_mux4_1 _5033_ (.S0(\game_logic_inst.lfsr_shift[0] ),
    .A0(\game_logic_inst.lfsr_value[1] ),
    .A1(\game_logic_inst.lfsr_value[5] ),
    .A2(\game_logic_inst.lfsr_value[9] ),
    .A3(\game_logic_inst.lfsr_value[13] ),
    .S1(\game_logic_inst.lfsr_shift[1] ),
    .X(_0716_));
 sg13g2_mux4_1 _5034_ (.S0(\game_logic_inst.lfsr_shift[0] ),
    .A0(\game_logic_inst.lfsr_value[0] ),
    .A1(\game_logic_inst.lfsr_value[4] ),
    .A2(\game_logic_inst.lfsr_value[8] ),
    .A3(\game_logic_inst.lfsr_value[12] ),
    .S1(\game_logic_inst.lfsr_shift[1] ),
    .X(_0717_));
 sg13g2_nand2_2 _5035_ (.Y(_0718_),
    .A(_0716_),
    .B(_0717_));
 sg13g2_nor4_1 _5036_ (.A(\debug_controller_inst.grid_in[28] ),
    .B(\debug_controller_inst.grid_in[29] ),
    .C(\debug_controller_inst.grid_in[30] ),
    .D(\debug_controller_inst.grid_in[31] ),
    .Y(_0719_));
 sg13g2_nand2b_2 _5037_ (.Y(_0720_),
    .B(_0716_),
    .A_N(_0717_));
 sg13g2_nor4_1 _5038_ (.A(\debug_controller_inst.grid_in[24] ),
    .B(\debug_controller_inst.grid_in[25] ),
    .C(\debug_controller_inst.grid_in[26] ),
    .D(\debug_controller_inst.grid_in[27] ),
    .Y(_0721_));
 sg13g2_nor2_1 _5039_ (.A(_0720_),
    .B(_0721_),
    .Y(_0722_));
 sg13g2_or2_2 _5040_ (.X(_0723_),
    .B(_0717_),
    .A(_0716_));
 sg13g2_nor4_1 _5041_ (.A(\debug_controller_inst.grid_in[16] ),
    .B(\debug_controller_inst.grid_in[17] ),
    .C(\debug_controller_inst.grid_in[18] ),
    .D(\debug_controller_inst.grid_in[19] ),
    .Y(_0724_));
 sg13g2_nand2b_2 _5042_ (.Y(_0725_),
    .B(_0717_),
    .A_N(_0716_));
 sg13g2_nor3_1 _5043_ (.A(\debug_controller_inst.grid_in[20] ),
    .B(\debug_controller_inst.grid_in[22] ),
    .C(\debug_controller_inst.grid_in[23] ),
    .Y(_0726_));
 sg13g2_a21oi_1 _5044_ (.A1(_3981_),
    .A2(_0726_),
    .Y(_0727_),
    .B1(_0725_));
 sg13g2_o21ai_1 _5045_ (.B1(_0715_),
    .Y(_0728_),
    .A1(_0723_),
    .A2(_0724_));
 sg13g2_nor3_1 _5046_ (.A(_0722_),
    .B(_0727_),
    .C(_0728_),
    .Y(_0729_));
 sg13g2_o21ai_1 _5047_ (.B1(_0729_),
    .Y(_0730_),
    .A1(_0718_),
    .A2(_0719_));
 sg13g2_nor4_1 _5048_ (.A(\debug_controller_inst.grid_in[0] ),
    .B(\debug_controller_inst.grid_in[1] ),
    .C(\debug_controller_inst.grid_in[2] ),
    .D(\debug_controller_inst.grid_in[3] ),
    .Y(_0731_));
 sg13g2_o21ai_1 _5049_ (.B1(_0714_),
    .Y(_0732_),
    .A1(_0723_),
    .A2(_0731_));
 sg13g2_nor4_1 _5050_ (.A(\debug_controller_inst.grid_in[12] ),
    .B(\debug_controller_inst.grid_in[13] ),
    .C(\debug_controller_inst.grid_in[14] ),
    .D(\debug_controller_inst.grid_in[15] ),
    .Y(_0733_));
 sg13g2_nor2_1 _5051_ (.A(_0718_),
    .B(_0733_),
    .Y(_0734_));
 sg13g2_nor4_1 _5052_ (.A(\debug_controller_inst.grid_in[4] ),
    .B(\debug_controller_inst.grid_in[5] ),
    .C(\debug_controller_inst.grid_in[6] ),
    .D(\debug_controller_inst.grid_in[7] ),
    .Y(_0735_));
 sg13g2_nor2_1 _5053_ (.A(_0725_),
    .B(_0735_),
    .Y(_0736_));
 sg13g2_nor4_1 _5054_ (.A(\debug_controller_inst.grid_in[8] ),
    .B(\debug_controller_inst.grid_in[9] ),
    .C(\debug_controller_inst.grid_in[10] ),
    .D(\debug_controller_inst.grid_in[11] ),
    .Y(_0737_));
 sg13g2_nor2_1 _5055_ (.A(_0720_),
    .B(_0737_),
    .Y(_0738_));
 sg13g2_nor4_1 _5056_ (.A(_0732_),
    .B(_0734_),
    .C(_0736_),
    .D(_0738_),
    .Y(_0739_));
 sg13g2_nor2_1 _5057_ (.A(_0707_),
    .B(_0739_),
    .Y(_0740_));
 sg13g2_nor4_1 _5058_ (.A(\debug_controller_inst.grid_in[44] ),
    .B(\debug_controller_inst.grid_in[45] ),
    .C(\debug_controller_inst.grid_in[46] ),
    .D(\debug_controller_inst.grid_in[47] ),
    .Y(_0741_));
 sg13g2_nor2_1 _5059_ (.A(_0718_),
    .B(_0741_),
    .Y(_0742_));
 sg13g2_nor4_1 _5060_ (.A(\debug_controller_inst.grid_in[36] ),
    .B(\debug_controller_inst.grid_in[37] ),
    .C(\debug_controller_inst.grid_in[38] ),
    .D(\debug_controller_inst.grid_in[39] ),
    .Y(_0743_));
 sg13g2_nor2_1 _5061_ (.A(_0725_),
    .B(_0743_),
    .Y(_0744_));
 sg13g2_nor4_1 _5062_ (.A(\debug_controller_inst.grid_in[32] ),
    .B(\debug_controller_inst.grid_in[33] ),
    .C(\debug_controller_inst.grid_in[34] ),
    .D(\debug_controller_inst.grid_in[35] ),
    .Y(_0745_));
 sg13g2_nor4_1 _5063_ (.A(\debug_controller_inst.grid_in[40] ),
    .B(\debug_controller_inst.grid_in[41] ),
    .C(\debug_controller_inst.grid_in[42] ),
    .D(\debug_controller_inst.grid_in[43] ),
    .Y(_0746_));
 sg13g2_nor2_1 _5064_ (.A(_0720_),
    .B(_0746_),
    .Y(_0747_));
 sg13g2_o21ai_1 _5065_ (.B1(_0714_),
    .Y(_0748_),
    .A1(_0723_),
    .A2(_0745_));
 sg13g2_nor4_1 _5066_ (.A(_0742_),
    .B(_0744_),
    .C(_0747_),
    .D(_0748_),
    .Y(_0749_));
 sg13g2_nor4_1 _5067_ (.A(\debug_controller_inst.grid_in[48] ),
    .B(\debug_controller_inst.grid_in[49] ),
    .C(\debug_controller_inst.grid_in[50] ),
    .D(\debug_controller_inst.grid_in[51] ),
    .Y(_0750_));
 sg13g2_nor2_1 _5068_ (.A(_0723_),
    .B(_0750_),
    .Y(_0751_));
 sg13g2_nor4_1 _5069_ (.A(\debug_controller_inst.grid_in[56] ),
    .B(\debug_controller_inst.grid_in[57] ),
    .C(\debug_controller_inst.grid_in[58] ),
    .D(\debug_controller_inst.grid_in[59] ),
    .Y(_0752_));
 sg13g2_nor2_1 _5070_ (.A(_0720_),
    .B(_0752_),
    .Y(_0753_));
 sg13g2_nor4_1 _5071_ (.A(\debug_controller_inst.grid_in[52] ),
    .B(\debug_controller_inst.grid_in[53] ),
    .C(\debug_controller_inst.grid_in[54] ),
    .D(\debug_controller_inst.grid_in[55] ),
    .Y(_0754_));
 sg13g2_nor4_1 _5072_ (.A(\debug_controller_inst.grid_in[60] ),
    .B(\debug_controller_inst.grid_in[61] ),
    .C(\debug_controller_inst.grid_in[62] ),
    .D(\debug_controller_inst.grid_in[63] ),
    .Y(_0755_));
 sg13g2_nor2_1 _5073_ (.A(_0718_),
    .B(_0755_),
    .Y(_0756_));
 sg13g2_o21ai_1 _5074_ (.B1(_0715_),
    .Y(_0757_),
    .A1(_0725_),
    .A2(_0754_));
 sg13g2_nor4_1 _5075_ (.A(_0751_),
    .B(_0753_),
    .C(_0756_),
    .D(_0757_),
    .Y(_0758_));
 sg13g2_nor3_2 _5076_ (.A(_0708_),
    .B(_0749_),
    .C(_0758_),
    .Y(_0759_));
 sg13g2_nor2_2 _5077_ (.A(\game_logic_inst.add_new_tiles[1] ),
    .B(\game_logic_inst.add_new_tiles[0] ),
    .Y(_0760_));
 sg13g2_a21oi_2 _5078_ (.B1(_0759_),
    .Y(_0761_),
    .A2(_0740_),
    .A1(_0730_));
 sg13g2_nand2b_1 _5079_ (.Y(_0762_),
    .B(_0761_),
    .A_N(_0760_));
 sg13g2_inv_1 _5080_ (.Y(_0763_),
    .A(_0762_));
 sg13g2_nor2_1 _5081_ (.A(_0707_),
    .B(_0762_),
    .Y(_0764_));
 sg13g2_nor2_1 _5082_ (.A(_0715_),
    .B(_0723_),
    .Y(_0765_));
 sg13g2_and2_1 _5083_ (.A(_0764_),
    .B(_0765_),
    .X(_0766_));
 sg13g2_nor3_1 _5084_ (.A(net2121),
    .B(_4009_),
    .C(_0766_),
    .Y(_0767_));
 sg13g2_nor3_1 _5085_ (.A(_0704_),
    .B(net1759),
    .C(_0767_),
    .Y(_0768_));
 sg13g2_o21ai_1 _5086_ (.B1(net2106),
    .Y(_0769_),
    .A1(net959),
    .A2(net1763));
 sg13g2_o21ai_1 _5087_ (.B1(net2275),
    .Y(_0770_),
    .A1(_4010_),
    .A2(_0532_));
 sg13g2_a21oi_1 _5088_ (.A1(net2057),
    .A2(net959),
    .Y(_0771_),
    .B1(_0770_));
 sg13g2_o21ai_1 _5089_ (.B1(_0771_),
    .Y(_0772_),
    .A1(_0768_),
    .A2(_0769_));
 sg13g2_nand2_1 _5090_ (.Y(_0003_),
    .A(_0534_),
    .B(_0772_));
 sg13g2_nand2_1 _5091_ (.Y(_0773_),
    .A(net2090),
    .B(_0533_));
 sg13g2_nor2_1 _5092_ (.A(_3940_),
    .B(net1761),
    .Y(_0774_));
 sg13g2_nand2_1 _5093_ (.Y(_0775_),
    .A(net2120),
    .B(net1762));
 sg13g2_or3_1 _5094_ (.A(_0100_),
    .B(net1759),
    .C(_0766_),
    .X(_0776_));
 sg13g2_and2_1 _5095_ (.A(_0653_),
    .B(_0658_),
    .X(_0777_));
 sg13g2_nand2_1 _5096_ (.Y(_0778_),
    .A(_0681_),
    .B(_0689_));
 sg13g2_nor2_1 _5097_ (.A(_0664_),
    .B(_0681_),
    .Y(_0779_));
 sg13g2_nand4_1 _5098_ (.B(_0685_),
    .C(_0687_),
    .A(_0684_),
    .Y(_0780_),
    .D(_0779_));
 sg13g2_a21o_1 _5099_ (.A2(_0780_),
    .A1(_0690_),
    .B1(_0695_),
    .X(_0781_));
 sg13g2_a22oi_1 _5100_ (.Y(_0782_),
    .B1(_0778_),
    .B2(_0781_),
    .A2(_0697_),
    .A1(_0653_));
 sg13g2_a21oi_2 _5101_ (.B1(_0782_),
    .Y(_0783_),
    .A2(_0695_),
    .A1(_0681_));
 sg13g2_a22oi_1 _5102_ (.Y(_0784_),
    .B1(_0783_),
    .B2(net2012),
    .A2(_0658_),
    .A1(_0651_));
 sg13g2_mux2_1 _5103_ (.A0(_0777_),
    .A1(_0783_),
    .S(net2015),
    .X(_0785_));
 sg13g2_nor2_1 _5104_ (.A(_0100_),
    .B(net2020),
    .Y(_0786_));
 sg13g2_a21oi_1 _5105_ (.A1(net2020),
    .A2(_0785_),
    .Y(_0787_),
    .B1(_0786_));
 sg13g2_a22oi_1 _5106_ (.Y(_0788_),
    .B1(_0787_),
    .B2(net2121),
    .A2(_0776_),
    .A1(net1734));
 sg13g2_o21ai_1 _5107_ (.B1(net2113),
    .Y(_0789_),
    .A1(net936),
    .A2(net1763));
 sg13g2_a21oi_1 _5108_ (.A1(net2057),
    .A2(net936),
    .Y(_0790_),
    .B1(_0770_));
 sg13g2_o21ai_1 _5109_ (.B1(_0790_),
    .Y(_0791_),
    .A1(_0788_),
    .A2(_0789_));
 sg13g2_nand2_1 _5110_ (.Y(_0014_),
    .A(_0773_),
    .B(net937));
 sg13g2_nor3_1 _5111_ (.A(net928),
    .B(net1759),
    .C(_0766_),
    .Y(_0792_));
 sg13g2_nand2_1 _5112_ (.Y(_0793_),
    .A(_0647_),
    .B(_0697_));
 sg13g2_a21o_1 _5113_ (.A2(_0793_),
    .A1(_0780_),
    .B1(_0695_),
    .X(_0794_));
 sg13g2_nand2b_1 _5114_ (.Y(_0795_),
    .B(_0670_),
    .A_N(_0780_));
 sg13g2_o21ai_1 _5115_ (.B1(_0690_),
    .Y(_0796_),
    .A1(_0671_),
    .A2(_0780_));
 sg13g2_and2_1 _5116_ (.A(_0696_),
    .B(_0796_),
    .X(_0797_));
 sg13g2_a22oi_1 _5117_ (.Y(_0798_),
    .B1(_0797_),
    .B2(_0793_),
    .A2(_0794_),
    .A1(_0671_));
 sg13g2_nand2_1 _5118_ (.Y(_0799_),
    .A(net2013),
    .B(_0798_));
 sg13g2_a22oi_1 _5119_ (.Y(_0800_),
    .B1(_0798_),
    .B2(net2012),
    .A2(_0658_),
    .A1(_0644_));
 sg13g2_a21oi_1 _5120_ (.A1(_4011_),
    .A2(net2018),
    .Y(_0801_),
    .B1(_3940_));
 sg13g2_o21ai_1 _5121_ (.B1(_0801_),
    .Y(_0802_),
    .A1(net2018),
    .A2(_0800_));
 sg13g2_o21ai_1 _5122_ (.B1(_0802_),
    .Y(_0803_),
    .A1(net1739),
    .A2(_0792_));
 sg13g2_a21oi_1 _5123_ (.A1(_4011_),
    .A2(net1759),
    .Y(_0804_),
    .B1(net2057));
 sg13g2_a221oi_1 _5124_ (.B2(_0804_),
    .C1(_0770_),
    .B1(_0803_),
    .A1(net2057),
    .Y(_0805_),
    .A2(net928));
 sg13g2_a21o_1 _5125_ (.A2(_0533_),
    .A1(net2088),
    .B1(_0805_),
    .X(_0025_));
 sg13g2_nor3_1 _5126_ (.A(net905),
    .B(net1759),
    .C(_0766_),
    .Y(_0806_));
 sg13g2_a21oi_1 _5127_ (.A1(_0696_),
    .A2(_0796_),
    .Y(_0807_),
    .B1(_0677_));
 sg13g2_nand2_1 _5128_ (.Y(_0808_),
    .A(net1918),
    .B(_0697_));
 sg13g2_nand2_1 _5129_ (.Y(_0809_),
    .A(_0677_),
    .B(_0690_));
 sg13g2_o21ai_1 _5130_ (.B1(_0808_),
    .Y(_0810_),
    .A1(_0795_),
    .A2(_0809_));
 sg13g2_o21ai_1 _5131_ (.B1(net2012),
    .Y(_0811_),
    .A1(_0807_),
    .A2(_0810_));
 sg13g2_nand3_1 _5132_ (.B(net1918),
    .C(_0658_),
    .A(net2011),
    .Y(_0812_));
 sg13g2_and2_2 _5133_ (.A(_0811_),
    .B(_0812_),
    .X(_0813_));
 sg13g2_a21oi_1 _5134_ (.A1(_4012_),
    .A2(net2018),
    .Y(_0814_),
    .B1(_3940_));
 sg13g2_o21ai_1 _5135_ (.B1(_0814_),
    .Y(_0815_),
    .A1(net2018),
    .A2(_0813_));
 sg13g2_o21ai_1 _5136_ (.B1(_0815_),
    .Y(_0816_),
    .A1(net1739),
    .A2(_0806_));
 sg13g2_a21oi_1 _5137_ (.A1(_4012_),
    .A2(net1759),
    .Y(_0817_),
    .B1(net2057));
 sg13g2_a221oi_1 _5138_ (.B2(_0817_),
    .C1(_0770_),
    .B1(_0816_),
    .A1(net2057),
    .Y(_0818_),
    .A2(net905));
 sg13g2_a21o_1 _5139_ (.A2(_0533_),
    .A1(net2086),
    .B1(_0818_),
    .X(_0036_));
 sg13g2_xnor2_1 _5140_ (.Y(_0819_),
    .A(\debug_controller_inst.grid_out_addr[3] ),
    .B(_0531_));
 sg13g2_nand2_2 _5141_ (.Y(_0820_),
    .A(\debug_controller_inst.grid_out_valid ),
    .B(_0819_));
 sg13g2_nand2b_2 _5142_ (.Y(_0821_),
    .B(\debug_controller_inst.grid_out_addr[0] ),
    .A_N(\debug_controller_inst.grid_out_addr[1] ));
 sg13g2_nor3_2 _5143_ (.A(net2084),
    .B(_0820_),
    .C(_0821_),
    .Y(_0822_));
 sg13g2_nor3_1 _5144_ (.A(_0561_),
    .B(_0566_),
    .C(net1764),
    .Y(_0823_));
 sg13g2_a21o_1 _5145_ (.A2(_0634_),
    .A1(_0594_),
    .B1(_0823_),
    .X(_0824_));
 sg13g2_o21ai_1 _5146_ (.B1(_0824_),
    .Y(_0825_),
    .A1(_0565_),
    .A2(_0629_));
 sg13g2_nand2b_1 _5147_ (.Y(_0826_),
    .B(_0570_),
    .A_N(_0598_));
 sg13g2_nor3_1 _5148_ (.A(_0566_),
    .B(net1764),
    .C(_0826_),
    .Y(_0827_));
 sg13g2_nor4_1 _5149_ (.A(_0566_),
    .B(_0592_),
    .C(net1764),
    .D(_0826_),
    .Y(_0828_));
 sg13g2_xnor2_1 _5150_ (.Y(_0829_),
    .A(_0592_),
    .B(_0827_));
 sg13g2_a221oi_1 _5151_ (.B2(_0625_),
    .C1(_0628_),
    .B1(_0622_),
    .A1(_0556_),
    .Y(_0830_),
    .A2(_0558_));
 sg13g2_nor2_1 _5152_ (.A(_0829_),
    .B(_0830_),
    .Y(_0831_));
 sg13g2_o21ai_1 _5153_ (.B1(_0646_),
    .Y(_0832_),
    .A1(_0829_),
    .A2(_0830_));
 sg13g2_or3_1 _5154_ (.A(_0646_),
    .B(_0829_),
    .C(_0830_),
    .X(_0833_));
 sg13g2_nor2b_1 _5155_ (.A(_0628_),
    .B_N(_0554_),
    .Y(_0834_));
 sg13g2_o21ai_1 _5156_ (.B1(_0834_),
    .Y(_0835_),
    .A1(_0623_),
    .A2(_0624_));
 sg13g2_mux2_1 _5157_ (.A0(_0596_),
    .A1(_0569_),
    .S(_0828_),
    .X(_0836_));
 sg13g2_and2_1 _5158_ (.A(_0835_),
    .B(_0836_),
    .X(_0837_));
 sg13g2_nand3_1 _5159_ (.B(_0835_),
    .C(_0836_),
    .A(net1918),
    .Y(_0838_));
 sg13g2_a21o_1 _5160_ (.A2(_0836_),
    .A1(_0835_),
    .B1(net1918),
    .X(_0839_));
 sg13g2_a221oi_1 _5161_ (.B2(_0625_),
    .C1(_0628_),
    .B1(_0622_),
    .A1(_0548_),
    .Y(_0840_),
    .A2(_0550_));
 sg13g2_xnor2_1 _5162_ (.Y(_0841_),
    .A(_0598_),
    .B(_0823_));
 sg13g2_nor2_2 _5163_ (.A(_0840_),
    .B(_0841_),
    .Y(_0842_));
 sg13g2_or3_1 _5164_ (.A(_0652_),
    .B(_0840_),
    .C(_0841_),
    .X(_0843_));
 sg13g2_o21ai_1 _5165_ (.B1(_0652_),
    .Y(_0844_),
    .A1(_0840_),
    .A2(_0841_));
 sg13g2_xnor2_1 _5166_ (.Y(_0845_),
    .A(net1919),
    .B(_0825_));
 sg13g2_and3_1 _5167_ (.X(_0846_),
    .A(_0634_),
    .B(_0843_),
    .C(_0844_));
 sg13g2_and4_1 _5168_ (.A(_0832_),
    .B(_0833_),
    .C(_0838_),
    .D(_0839_),
    .X(_0847_));
 sg13g2_and3_1 _5169_ (.X(_0848_),
    .A(_0845_),
    .B(_0846_),
    .C(_0847_));
 sg13g2_a21oi_2 _5170_ (.B1(_0632_),
    .Y(_0849_),
    .A2(_0627_),
    .A1(_0566_));
 sg13g2_nor2b_2 _5171_ (.A(_0848_),
    .B_N(_0849_),
    .Y(_0850_));
 sg13g2_nor2b_1 _5172_ (.A(_0642_),
    .B_N(_0657_),
    .Y(_0851_));
 sg13g2_xnor2_1 _5173_ (.Y(_0852_),
    .A(_0642_),
    .B(_0657_));
 sg13g2_a22oi_1 _5174_ (.Y(_0853_),
    .B1(_0852_),
    .B2(_0637_),
    .A2(_0850_),
    .A1(net1919));
 sg13g2_nor3_1 _5175_ (.A(_0637_),
    .B(_0694_),
    .C(_0697_),
    .Y(_0854_));
 sg13g2_o21ai_1 _5176_ (.B1(_0693_),
    .Y(_0855_),
    .A1(_0690_),
    .A2(_0849_));
 sg13g2_nand4_1 _5177_ (.B(_0685_),
    .C(_0687_),
    .A(_0684_),
    .Y(_0856_),
    .D(_0690_));
 sg13g2_nand3b_1 _5178_ (.B(_0854_),
    .C(_0856_),
    .Y(_0857_),
    .A_N(_0850_));
 sg13g2_nor2_1 _5179_ (.A(_0688_),
    .B(_0691_),
    .Y(_0858_));
 sg13g2_nand2_1 _5180_ (.Y(_0859_),
    .A(_0848_),
    .B(_0849_));
 sg13g2_nor2_1 _5181_ (.A(_0825_),
    .B(_0859_),
    .Y(_0860_));
 sg13g2_a221oi_1 _5182_ (.B2(net1919),
    .C1(_0860_),
    .B1(_0858_),
    .A1(_0825_),
    .Y(_0861_),
    .A2(_0857_));
 sg13g2_mux2_2 _5183_ (.A0(_0853_),
    .A1(_0861_),
    .S(net2015),
    .X(_0862_));
 sg13g2_nor2_1 _5184_ (.A(_0103_),
    .B(net2020),
    .Y(_0863_));
 sg13g2_o21ai_1 _5185_ (.B1(net1737),
    .Y(_0864_),
    .A1(net2016),
    .A2(_0862_));
 sg13g2_nor2_1 _5186_ (.A(_3938_),
    .B(net1776),
    .Y(_0865_));
 sg13g2_nor2_2 _5187_ (.A(_0715_),
    .B(_0725_),
    .Y(_0866_));
 sg13g2_nor3_2 _5188_ (.A(net1776),
    .B(_0707_),
    .C(_0762_),
    .Y(_0867_));
 sg13g2_nor2_2 _5189_ (.A(\game_logic_inst.should_transpose ),
    .B(net2120),
    .Y(_0868_));
 sg13g2_nand2_2 _5190_ (.Y(_0869_),
    .A(_3938_),
    .B(_3940_));
 sg13g2_nand2_1 _5191_ (.Y(_0870_),
    .A(net1775),
    .B(net1917));
 sg13g2_nand2_1 _5192_ (.Y(_0871_),
    .A(_0103_),
    .B(net1745));
 sg13g2_a21oi_1 _5193_ (.A1(_0866_),
    .A2(net1728),
    .Y(_0872_),
    .B1(_0871_));
 sg13g2_a21oi_1 _5194_ (.A1(net914),
    .A2(net1750),
    .Y(_0873_),
    .B1(_0872_));
 sg13g2_o21ai_1 _5195_ (.B1(_0873_),
    .Y(_0874_),
    .A1(_0863_),
    .A2(_0864_));
 sg13g2_nand2_1 _5196_ (.Y(_0875_),
    .A(net2104),
    .B(_0874_));
 sg13g2_nand2b_2 _5197_ (.Y(_0876_),
    .B(net2269),
    .A_N(_0822_));
 sg13g2_a21oi_1 _5198_ (.A1(net2053),
    .A2(net935),
    .Y(_0877_),
    .B1(_0876_));
 sg13g2_a22oi_1 _5199_ (.Y(_0878_),
    .B1(_0875_),
    .B2(_0877_),
    .A2(_0822_),
    .A1(net2092));
 sg13g2_inv_1 _5200_ (.Y(_0047_),
    .A(_0878_));
 sg13g2_nand2_2 _5201_ (.Y(_0879_),
    .A(_0551_),
    .B(_0851_));
 sg13g2_nand2_1 _5202_ (.Y(_0880_),
    .A(_0637_),
    .B(_0879_));
 sg13g2_nand4_1 _5203_ (.B(_0693_),
    .C(_0859_),
    .A(_0636_),
    .Y(_0881_),
    .D(_0880_));
 sg13g2_and3_1 _5204_ (.X(_0882_),
    .A(_0637_),
    .B(_0851_),
    .C(_0879_));
 sg13g2_a221oi_1 _5205_ (.B2(_0654_),
    .C1(_0882_),
    .B1(_0881_),
    .A1(_0653_),
    .Y(_0883_),
    .A2(_0850_));
 sg13g2_nand2_1 _5206_ (.Y(_0884_),
    .A(_0842_),
    .B(_0855_));
 sg13g2_nor3_1 _5207_ (.A(_0652_),
    .B(_0688_),
    .C(_0691_),
    .Y(_0885_));
 sg13g2_nand4_1 _5208_ (.B(_0845_),
    .C(_0846_),
    .A(_0825_),
    .Y(_0886_),
    .D(_0847_));
 sg13g2_o21ai_1 _5209_ (.B1(_0849_),
    .Y(_0887_),
    .A1(_0842_),
    .A2(_0886_));
 sg13g2_a22oi_1 _5210_ (.Y(_0888_),
    .B1(_0887_),
    .B2(_0854_),
    .A2(_0886_),
    .A1(_0842_));
 sg13g2_o21ai_1 _5211_ (.B1(_0884_),
    .Y(_0889_),
    .A1(_0885_),
    .A2(_0888_));
 sg13g2_mux2_2 _5212_ (.A0(_0883_),
    .A1(_0889_),
    .S(net2015),
    .X(_0890_));
 sg13g2_a21oi_1 _5213_ (.A1(_4013_),
    .A2(net2016),
    .Y(_0891_),
    .B1(net1733));
 sg13g2_o21ai_1 _5214_ (.B1(_0891_),
    .Y(_0892_),
    .A1(net2016),
    .A2(_0890_));
 sg13g2_a22oi_1 _5215_ (.Y(_0893_),
    .B1(net1744),
    .B2(net907),
    .A2(net1750),
    .A1(_0106_));
 sg13g2_nand3_1 _5216_ (.B(net1728),
    .C(_0868_),
    .A(_0866_),
    .Y(_0894_));
 sg13g2_nor2_2 _5217_ (.A(net1776),
    .B(net1917),
    .Y(_0895_));
 sg13g2_nand3_1 _5218_ (.B(_0893_),
    .C(_0894_),
    .A(_0892_),
    .Y(_0896_));
 sg13g2_nand2_1 _5219_ (.Y(_0897_),
    .A(net2104),
    .B(_0896_));
 sg13g2_a21oi_1 _5220_ (.A1(net2053),
    .A2(net907),
    .Y(_0898_),
    .B1(_0876_));
 sg13g2_a22oi_1 _5221_ (.Y(_0899_),
    .B1(_0897_),
    .B2(_0898_),
    .A2(_0822_),
    .A1(net2090));
 sg13g2_inv_1 _5222_ (.Y(_0058_),
    .A(net908));
 sg13g2_o21ai_1 _5223_ (.B1(_0637_),
    .Y(_0900_),
    .A1(_0649_),
    .A2(_0879_));
 sg13g2_nor2_1 _5224_ (.A(_0879_),
    .B(_0900_),
    .Y(_0901_));
 sg13g2_a221oi_1 _5225_ (.B2(_0648_),
    .C1(_0901_),
    .B1(_0881_),
    .A1(_0647_),
    .Y(_0902_),
    .A2(_0850_));
 sg13g2_or3_1 _5226_ (.A(_0831_),
    .B(_0842_),
    .C(_0886_),
    .X(_0903_));
 sg13g2_and2_1 _5227_ (.A(_0849_),
    .B(_0903_),
    .X(_0904_));
 sg13g2_o21ai_1 _5228_ (.B1(_0831_),
    .Y(_0905_),
    .A1(_0842_),
    .A2(_0886_));
 sg13g2_a221oi_1 _5229_ (.B2(_0905_),
    .C1(_0855_),
    .B1(_0904_),
    .A1(_0647_),
    .Y(_0906_),
    .A2(_0858_));
 sg13g2_a21o_1 _5230_ (.A2(_0855_),
    .A1(_0831_),
    .B1(_0906_),
    .X(_0907_));
 sg13g2_mux2_2 _5231_ (.A0(_0902_),
    .A1(_0907_),
    .S(net2015),
    .X(_0908_));
 sg13g2_o21ai_1 _5232_ (.B1(net1737),
    .Y(_0909_),
    .A1(net2017),
    .A2(_0908_));
 sg13g2_a21oi_1 _5233_ (.A1(_4015_),
    .A2(net2016),
    .Y(_0910_),
    .B1(_0909_));
 sg13g2_a22oi_1 _5234_ (.Y(_0911_),
    .B1(net1744),
    .B2(net900),
    .A2(net1750),
    .A1(_0108_));
 sg13g2_nand2_1 _5235_ (.Y(_0912_),
    .A(_0894_),
    .B(_0911_));
 sg13g2_o21ai_1 _5236_ (.B1(net2106),
    .Y(_0913_),
    .A1(_0910_),
    .A2(_0912_));
 sg13g2_a21oi_1 _5237_ (.A1(net2054),
    .A2(net900),
    .Y(_0914_),
    .B1(_0876_));
 sg13g2_a22oi_1 _5238_ (.Y(_0915_),
    .B1(_0913_),
    .B2(_0914_),
    .A2(_0822_),
    .A1(net2088));
 sg13g2_inv_1 _5239_ (.Y(_0063_),
    .A(net901));
 sg13g2_nand4_1 _5240_ (.B(_0693_),
    .C(_0859_),
    .A(_0636_),
    .Y(_0916_),
    .D(_0900_));
 sg13g2_nor3_1 _5241_ (.A(_0554_),
    .B(_0649_),
    .C(_0879_),
    .Y(_0917_));
 sg13g2_a221oi_1 _5242_ (.B2(_0639_),
    .C1(_0917_),
    .B1(_0916_),
    .A1(net1918),
    .Y(_0918_),
    .A2(_0850_));
 sg13g2_a221oi_1 _5243_ (.B2(_0903_),
    .C1(_0855_),
    .B1(_0849_),
    .A1(_0688_),
    .Y(_0919_),
    .A2(_0690_));
 sg13g2_nor2_1 _5244_ (.A(_0837_),
    .B(_0919_),
    .Y(_0920_));
 sg13g2_nand2_1 _5245_ (.Y(_0921_),
    .A(_0837_),
    .B(_0849_));
 sg13g2_nor2_1 _5246_ (.A(_0903_),
    .B(_0921_),
    .Y(_0922_));
 sg13g2_a21oi_1 _5247_ (.A1(net1918),
    .A2(_0858_),
    .Y(_0923_),
    .B1(_0922_));
 sg13g2_nor2b_1 _5248_ (.A(_0920_),
    .B_N(_0923_),
    .Y(_0924_));
 sg13g2_mux2_2 _5249_ (.A0(_0918_),
    .A1(_0924_),
    .S(net2015),
    .X(_0925_));
 sg13g2_o21ai_1 _5250_ (.B1(net1737),
    .Y(_0926_),
    .A1(net2016),
    .A2(_0925_));
 sg13g2_a21oi_1 _5251_ (.A1(_4017_),
    .A2(net2016),
    .Y(_0927_),
    .B1(_0926_));
 sg13g2_a22oi_1 _5252_ (.Y(_0928_),
    .B1(net1744),
    .B2(net924),
    .A2(net1750),
    .A1(net1047));
 sg13g2_nand2_1 _5253_ (.Y(_0929_),
    .A(_0894_),
    .B(_0928_));
 sg13g2_o21ai_1 _5254_ (.B1(net2104),
    .Y(_0930_),
    .A1(_0927_),
    .A2(_0929_));
 sg13g2_a21oi_1 _5255_ (.A1(net2053),
    .A2(net924),
    .Y(_0931_),
    .B1(_0876_));
 sg13g2_a22oi_1 _5256_ (.Y(_0932_),
    .B1(_0930_),
    .B2(_0931_),
    .A2(_0822_),
    .A1(net2086));
 sg13g2_inv_1 _5257_ (.Y(_0064_),
    .A(_0932_));
 sg13g2_nand2_1 _5258_ (.Y(_0933_),
    .A(net2093),
    .B(_0532_));
 sg13g2_nor2b_1 _5259_ (.A(\debug_controller_inst.grid_out_addr[0] ),
    .B_N(\debug_controller_inst.grid_out_addr[1] ),
    .Y(_0934_));
 sg13g2_nor2b_2 _5260_ (.A(net2085),
    .B_N(_0934_),
    .Y(_0935_));
 sg13g2_nand3_1 _5261_ (.B(_0819_),
    .C(_0935_),
    .A(\debug_controller_inst.grid_out_valid ),
    .Y(_0936_));
 sg13g2_mux2_2 _5262_ (.A0(_0853_),
    .A1(_0861_),
    .S(net2011),
    .X(_0937_));
 sg13g2_nor2_1 _5263_ (.A(_0111_),
    .B(net2020),
    .Y(_0938_));
 sg13g2_o21ai_1 _5264_ (.B1(net1739),
    .Y(_0939_),
    .A1(net2018),
    .A2(_0937_));
 sg13g2_nor2_1 _5265_ (.A(_0715_),
    .B(_0720_),
    .Y(_0940_));
 sg13g2_nand2_1 _5266_ (.Y(_0941_),
    .A(_0111_),
    .B(net1748));
 sg13g2_a21oi_1 _5267_ (.A1(_0867_),
    .A2(_0940_),
    .Y(_0942_),
    .B1(_0941_));
 sg13g2_a21oi_1 _5268_ (.A1(_0112_),
    .A2(net1756),
    .Y(_0943_),
    .B1(_0942_));
 sg13g2_o21ai_1 _5269_ (.B1(_0943_),
    .Y(_0944_),
    .A1(_0938_),
    .A2(_0939_));
 sg13g2_nand2_1 _5270_ (.Y(_0945_),
    .A(net2113),
    .B(_0944_));
 sg13g2_nand2_1 _5271_ (.Y(_0946_),
    .A(net2058),
    .B(net902));
 sg13g2_and2_1 _5272_ (.A(net2275),
    .B(_0936_),
    .X(_0947_));
 sg13g2_nand3_1 _5273_ (.B(_0946_),
    .C(_0947_),
    .A(_0945_),
    .Y(_0948_));
 sg13g2_o21ai_1 _5274_ (.B1(net903),
    .Y(_0065_),
    .A1(_0933_),
    .A2(_0936_));
 sg13g2_nand2_2 _5275_ (.Y(_0949_),
    .A(net2091),
    .B(_0532_));
 sg13g2_mux2_2 _5276_ (.A0(_0883_),
    .A1(_0889_),
    .S(net2011),
    .X(_0950_));
 sg13g2_o21ai_1 _5277_ (.B1(net1739),
    .Y(_0951_),
    .A1(net2019),
    .A2(_0950_));
 sg13g2_a21oi_1 _5278_ (.A1(_4020_),
    .A2(net2019),
    .Y(_0952_),
    .B1(_0951_));
 sg13g2_a22oi_1 _5279_ (.Y(_0953_),
    .B1(net1748),
    .B2(net919),
    .A2(net1756),
    .A1(_0114_));
 sg13g2_nand3_1 _5280_ (.B(_0868_),
    .C(_0940_),
    .A(net1728),
    .Y(_0954_));
 sg13g2_nand2_1 _5281_ (.Y(_0955_),
    .A(_0953_),
    .B(_0954_));
 sg13g2_o21ai_1 _5282_ (.B1(net2111),
    .Y(_0956_),
    .A1(_0952_),
    .A2(_0955_));
 sg13g2_nand2_1 _5283_ (.Y(_0957_),
    .A(net2058),
    .B(net919));
 sg13g2_nand3_1 _5284_ (.B(_0956_),
    .C(_0957_),
    .A(_0947_),
    .Y(_0958_));
 sg13g2_o21ai_1 _5285_ (.B1(net920),
    .Y(_0066_),
    .A1(_0936_),
    .A2(_0949_));
 sg13g2_nand2_2 _5286_ (.Y(_0959_),
    .A(net2089),
    .B(_0532_));
 sg13g2_mux2_2 _5287_ (.A0(_0902_),
    .A1(_0907_),
    .S(net2011),
    .X(_0960_));
 sg13g2_o21ai_1 _5288_ (.B1(net1739),
    .Y(_0961_),
    .A1(net2019),
    .A2(_0960_));
 sg13g2_a21oi_1 _5289_ (.A1(_4022_),
    .A2(net2018),
    .Y(_0962_),
    .B1(_0961_));
 sg13g2_a22oi_1 _5290_ (.Y(_0963_),
    .B1(net1748),
    .B2(net967),
    .A2(net1756),
    .A1(_0116_));
 sg13g2_nand2_1 _5291_ (.Y(_0964_),
    .A(_0954_),
    .B(_0963_));
 sg13g2_o21ai_1 _5292_ (.B1(net2111),
    .Y(_0965_),
    .A1(_0962_),
    .A2(_0964_));
 sg13g2_nand2_1 _5293_ (.Y(_0966_),
    .A(net2058),
    .B(net967));
 sg13g2_nand3_1 _5294_ (.B(_0965_),
    .C(_0966_),
    .A(_0947_),
    .Y(_0967_));
 sg13g2_o21ai_1 _5295_ (.B1(net968),
    .Y(_0004_),
    .A1(_0936_),
    .A2(_0959_));
 sg13g2_nand2_2 _5296_ (.Y(_0968_),
    .A(net2087),
    .B(_0532_));
 sg13g2_mux2_2 _5297_ (.A0(_0918_),
    .A1(_0924_),
    .S(net2011),
    .X(_0969_));
 sg13g2_o21ai_1 _5298_ (.B1(net1739),
    .Y(_0970_),
    .A1(net2018),
    .A2(_0969_));
 sg13g2_a21oi_1 _5299_ (.A1(_4024_),
    .A2(net2018),
    .Y(_0971_),
    .B1(_0970_));
 sg13g2_a22oi_1 _5300_ (.Y(_0972_),
    .B1(net1748),
    .B2(net942),
    .A2(net1756),
    .A1(_0118_));
 sg13g2_nand2_1 _5301_ (.Y(_0973_),
    .A(_0954_),
    .B(_0972_));
 sg13g2_o21ai_1 _5302_ (.B1(net2112),
    .Y(_0974_),
    .A1(_0971_),
    .A2(_0973_));
 sg13g2_nand2_1 _5303_ (.Y(_0975_),
    .A(net2057),
    .B(net942));
 sg13g2_nand3_1 _5304_ (.B(_0974_),
    .C(_0975_),
    .A(_0947_),
    .Y(_0976_));
 sg13g2_o21ai_1 _5305_ (.B1(net943),
    .Y(_0005_),
    .A1(_0936_),
    .A2(_0968_));
 sg13g2_nand2_2 _5306_ (.Y(_0977_),
    .A(\debug_controller_inst.grid_out_addr[1] ),
    .B(\debug_controller_inst.grid_out_addr[0] ));
 sg13g2_nor3_2 _5307_ (.A(net2084),
    .B(_0820_),
    .C(_0977_),
    .Y(_0978_));
 sg13g2_nor2_1 _5308_ (.A(net2010),
    .B(_0659_),
    .Y(_0979_));
 sg13g2_a21o_2 _5309_ (.A2(_0700_),
    .A1(net2010),
    .B1(_0979_),
    .X(_0980_));
 sg13g2_nor2_1 _5310_ (.A(net1028),
    .B(net2020),
    .Y(_0981_));
 sg13g2_o21ai_1 _5311_ (.B1(net1738),
    .Y(_0982_),
    .A1(net2016),
    .A2(_0980_));
 sg13g2_nor2_2 _5312_ (.A(_0715_),
    .B(_0718_),
    .Y(_0983_));
 sg13g2_a21oi_1 _5313_ (.A1(net1728),
    .A2(_0983_),
    .Y(_0984_),
    .B1(_4026_));
 sg13g2_a22oi_1 _5314_ (.Y(_0985_),
    .B1(net1744),
    .B2(_0984_),
    .A2(net1751),
    .A1(net881));
 sg13g2_o21ai_1 _5315_ (.B1(_0985_),
    .Y(_0986_),
    .A1(_0981_),
    .A2(_0982_));
 sg13g2_nor2_2 _5316_ (.A(net2258),
    .B(_0978_),
    .Y(_0987_));
 sg13g2_o21ai_1 _5317_ (.B1(_0987_),
    .Y(_0988_),
    .A1(net2105),
    .A2(_4026_));
 sg13g2_a21oi_1 _5318_ (.A1(net2105),
    .A2(_0986_),
    .Y(_0989_),
    .B1(_0988_));
 sg13g2_a21o_1 _5319_ (.A2(_0978_),
    .A1(net2092),
    .B1(_0989_),
    .X(_0006_));
 sg13g2_mux2_2 _5320_ (.A0(_0777_),
    .A1(_0783_),
    .S(net2011),
    .X(_0990_));
 sg13g2_a21oi_1 _5321_ (.A1(net2020),
    .A2(_0990_),
    .Y(_0991_),
    .B1(net1733));
 sg13g2_o21ai_1 _5322_ (.B1(_0991_),
    .Y(_0992_),
    .A1(net1035),
    .A2(net2020));
 sg13g2_nand3_1 _5323_ (.B(_0868_),
    .C(_0983_),
    .A(net1728),
    .Y(_0993_));
 sg13g2_a22oi_1 _5324_ (.Y(_0994_),
    .B1(net1744),
    .B2(net1035),
    .A2(net1751),
    .A1(net878));
 sg13g2_nand3_1 _5325_ (.B(_0993_),
    .C(_0994_),
    .A(_0992_),
    .Y(_0995_));
 sg13g2_o21ai_1 _5326_ (.B1(_0987_),
    .Y(_0996_),
    .A1(net2105),
    .A2(_4027_));
 sg13g2_a21oi_1 _5327_ (.A1(net2105),
    .A2(_0995_),
    .Y(_0997_),
    .B1(_0996_));
 sg13g2_a21o_1 _5328_ (.A2(_0978_),
    .A1(net2090),
    .B1(_0997_),
    .X(_0007_));
 sg13g2_nand2_1 _5329_ (.Y(_0998_),
    .A(net2010),
    .B(_0798_));
 sg13g2_a22oi_1 _5330_ (.Y(_0999_),
    .B1(_0798_),
    .B2(net2010),
    .A2(_0658_),
    .A1(_0645_));
 sg13g2_nand2_1 _5331_ (.Y(_1000_),
    .A(_4028_),
    .B(net2017));
 sg13g2_o21ai_1 _5332_ (.B1(_1000_),
    .Y(_1001_),
    .A1(net2017),
    .A2(_0999_));
 sg13g2_nand2_1 _5333_ (.Y(_1002_),
    .A(_4028_),
    .B(_0993_));
 sg13g2_a22oi_1 _5334_ (.Y(_1003_),
    .B1(net1745),
    .B2(_1002_),
    .A2(net1751),
    .A1(net869));
 sg13g2_o21ai_1 _5335_ (.B1(_1003_),
    .Y(_1004_),
    .A1(net1733),
    .A2(_1001_));
 sg13g2_o21ai_1 _5336_ (.B1(_0987_),
    .Y(_1005_),
    .A1(net2105),
    .A2(_4028_));
 sg13g2_a21oi_1 _5337_ (.A1(net2105),
    .A2(_1004_),
    .Y(_1006_),
    .B1(_1005_));
 sg13g2_a21o_1 _5338_ (.A2(_0978_),
    .A1(net2088),
    .B1(_1006_),
    .X(_0008_));
 sg13g2_o21ai_1 _5339_ (.B1(net2010),
    .Y(_1007_),
    .A1(_0807_),
    .A2(_0810_));
 sg13g2_nand3_1 _5340_ (.B(net1918),
    .C(_0658_),
    .A(net2012),
    .Y(_1008_));
 sg13g2_and2_2 _5341_ (.A(_1007_),
    .B(_1008_),
    .X(_1009_));
 sg13g2_o21ai_1 _5342_ (.B1(net1738),
    .Y(_1010_),
    .A1(net2017),
    .A2(_1009_));
 sg13g2_a21o_1 _5343_ (.A2(net2017),
    .A1(_4029_),
    .B1(_1010_),
    .X(_1011_));
 sg13g2_a22oi_1 _5344_ (.Y(_1012_),
    .B1(net1745),
    .B2(net891),
    .A2(net1751),
    .A1(_0126_));
 sg13g2_nand3_1 _5345_ (.B(_1011_),
    .C(_1012_),
    .A(_0993_),
    .Y(_1013_));
 sg13g2_o21ai_1 _5346_ (.B1(_0987_),
    .Y(_1014_),
    .A1(net2106),
    .A2(_4029_));
 sg13g2_a21oi_1 _5347_ (.A1(net2106),
    .A2(_1013_),
    .Y(_1015_),
    .B1(_1014_));
 sg13g2_a21o_1 _5348_ (.A2(_0978_),
    .A1(net2086),
    .B1(_1015_),
    .X(_0009_));
 sg13g2_nand2_2 _5349_ (.Y(_1016_),
    .A(net2084),
    .B(_0530_));
 sg13g2_nor2_2 _5350_ (.A(_0820_),
    .B(_1016_),
    .Y(_1017_));
 sg13g2_nor2_2 _5351_ (.A(_0098_),
    .B(net2020),
    .Y(_1018_));
 sg13g2_nand2b_2 _5352_ (.Y(_1019_),
    .B(net2016),
    .A_N(_0098_));
 sg13g2_and3_1 _5353_ (.X(_1020_),
    .A(net1998),
    .B(_0702_),
    .C(_1018_));
 sg13g2_o21ai_1 _5354_ (.B1(net1737),
    .Y(_1021_),
    .A1(_0104_),
    .A2(net2006));
 sg13g2_nor2_2 _5355_ (.A(_0714_),
    .B(_0723_),
    .Y(_1022_));
 sg13g2_nand2_1 _5356_ (.Y(_1023_),
    .A(net1728),
    .B(_1022_));
 sg13g2_nand3_1 _5357_ (.B(net1745),
    .C(_1023_),
    .A(_0104_),
    .Y(_1024_));
 sg13g2_o21ai_1 _5358_ (.B1(_1024_),
    .Y(_1025_),
    .A1(_1020_),
    .A2(_1021_));
 sg13g2_a21oi_1 _5359_ (.A1(_0103_),
    .A2(net1750),
    .Y(_1026_),
    .B1(_1025_));
 sg13g2_nor2_2 _5360_ (.A(net2258),
    .B(_1017_),
    .Y(_1027_));
 sg13g2_o21ai_1 _5361_ (.B1(_1027_),
    .Y(_1028_),
    .A1(net2053),
    .A2(_1026_));
 sg13g2_a21oi_1 _5362_ (.A1(net2053),
    .A2(net914),
    .Y(_1029_),
    .B1(_1028_));
 sg13g2_a21o_1 _5363_ (.A2(_1017_),
    .A1(net2092),
    .B1(_1029_),
    .X(_0010_));
 sg13g2_nand2_1 _5364_ (.Y(_1030_),
    .A(net2090),
    .B(_1017_));
 sg13g2_nor2_2 _5365_ (.A(_0784_),
    .B(_1019_),
    .Y(_1031_));
 sg13g2_o21ai_1 _5366_ (.B1(net1737),
    .Y(_1032_),
    .A1(_0106_),
    .A2(net2006));
 sg13g2_a21oi_1 _5367_ (.A1(net1998),
    .A2(_1031_),
    .Y(_1033_),
    .B1(_1032_));
 sg13g2_nand3_1 _5368_ (.B(_0868_),
    .C(_1022_),
    .A(net1728),
    .Y(_1034_));
 sg13g2_a221oi_1 _5369_ (.B2(net981),
    .C1(_1033_),
    .B1(net1744),
    .A1(net907),
    .Y(_1035_),
    .A2(net1750));
 sg13g2_a21oi_1 _5370_ (.A1(_1034_),
    .A2(_1035_),
    .Y(_1036_),
    .B1(net2053));
 sg13g2_o21ai_1 _5371_ (.B1(_1027_),
    .Y(_1037_),
    .A1(net2104),
    .A2(_4014_));
 sg13g2_o21ai_1 _5372_ (.B1(_1030_),
    .Y(_0011_),
    .A1(_1036_),
    .A2(_1037_));
 sg13g2_nand2_1 _5373_ (.Y(_1038_),
    .A(net2088),
    .B(_1017_));
 sg13g2_nor2_1 _5374_ (.A(_0800_),
    .B(net1914),
    .Y(_1039_));
 sg13g2_o21ai_1 _5375_ (.B1(net1738),
    .Y(_1040_),
    .A1(_0108_),
    .A2(net2006));
 sg13g2_a21oi_1 _5376_ (.A1(net1998),
    .A2(_1039_),
    .Y(_1041_),
    .B1(_1040_));
 sg13g2_a221oi_1 _5377_ (.B2(net1000),
    .C1(_1041_),
    .B1(net1744),
    .A1(net900),
    .Y(_1042_),
    .A2(net1750));
 sg13g2_a21oi_1 _5378_ (.A1(_1034_),
    .A2(_1042_),
    .Y(_1043_),
    .B1(net2054));
 sg13g2_o21ai_1 _5379_ (.B1(_1027_),
    .Y(_1044_),
    .A1(net2106),
    .A2(_4016_));
 sg13g2_o21ai_1 _5380_ (.B1(_1038_),
    .Y(_0012_),
    .A1(_1043_),
    .A2(_1044_));
 sg13g2_nand2_1 _5381_ (.Y(_1045_),
    .A(net2086),
    .B(_1017_));
 sg13g2_nor2_1 _5382_ (.A(_0813_),
    .B(net1914),
    .Y(_1046_));
 sg13g2_o21ai_1 _5383_ (.B1(net1737),
    .Y(_1047_),
    .A1(net1048),
    .A2(net2006));
 sg13g2_a21oi_1 _5384_ (.A1(net1998),
    .A2(_1046_),
    .Y(_1048_),
    .B1(_1047_));
 sg13g2_a221oi_1 _5385_ (.B2(net997),
    .C1(_1048_),
    .B1(net1744),
    .A1(net924),
    .Y(_1049_),
    .A2(net1750));
 sg13g2_a21oi_1 _5386_ (.A1(_1034_),
    .A2(_1049_),
    .Y(_1050_),
    .B1(net2053));
 sg13g2_o21ai_1 _5387_ (.B1(_1027_),
    .Y(_1051_),
    .A1(net2104),
    .A2(_4018_));
 sg13g2_o21ai_1 _5388_ (.B1(_1045_),
    .Y(_0013_),
    .A1(_1050_),
    .A2(_1051_));
 sg13g2_nand3b_1 _5389_ (.B(\debug_controller_inst.grid_out_addr[0] ),
    .C(net2084),
    .Y(_1052_),
    .A_N(\debug_controller_inst.grid_out_addr[1] ));
 sg13g2_nor2_2 _5390_ (.A(_0820_),
    .B(_1052_),
    .Y(_1053_));
 sg13g2_nor2_2 _5391_ (.A(_0862_),
    .B(net1915),
    .Y(_1054_));
 sg13g2_o21ai_1 _5392_ (.B1(net2118),
    .Y(_1055_),
    .A1(_0127_),
    .A2(net2007));
 sg13g2_a21oi_1 _5393_ (.A1(net1997),
    .A2(_1054_),
    .Y(_1056_),
    .B1(_1055_));
 sg13g2_nor2_1 _5394_ (.A(_0714_),
    .B(_0725_),
    .Y(_1057_));
 sg13g2_and2_2 _5395_ (.A(_0764_),
    .B(_1057_),
    .X(_1058_));
 sg13g2_nor3_1 _5396_ (.A(net2118),
    .B(_4030_),
    .C(_1058_),
    .Y(_1059_));
 sg13g2_nor3_1 _5397_ (.A(net1758),
    .B(_1056_),
    .C(_1059_),
    .Y(_1060_));
 sg13g2_o21ai_1 _5398_ (.B1(net2108),
    .Y(_1061_),
    .A1(_0127_),
    .A2(net1762));
 sg13g2_nor2_2 _5399_ (.A(net2258),
    .B(_1053_),
    .Y(_1062_));
 sg13g2_o21ai_1 _5400_ (.B1(_1062_),
    .Y(_1063_),
    .A1(_1060_),
    .A2(_1061_));
 sg13g2_a21oi_1 _5401_ (.A1(net2055),
    .A2(net957),
    .Y(_1064_),
    .B1(_1063_));
 sg13g2_a21o_1 _5402_ (.A2(_1053_),
    .A1(net2092),
    .B1(_1064_),
    .X(_0015_));
 sg13g2_or3_1 _5403_ (.A(_0128_),
    .B(net1758),
    .C(_1058_),
    .X(_1065_));
 sg13g2_nor2_1 _5404_ (.A(_0890_),
    .B(net1914),
    .Y(_1066_));
 sg13g2_nor2_1 _5405_ (.A(_0128_),
    .B(net2007),
    .Y(_1067_));
 sg13g2_a21oi_1 _5406_ (.A1(net1997),
    .A2(_1066_),
    .Y(_1068_),
    .B1(_1067_));
 sg13g2_a22oi_1 _5407_ (.Y(_1069_),
    .B1(_1068_),
    .B2(net2118),
    .A2(_1065_),
    .A1(net1736));
 sg13g2_o21ai_1 _5408_ (.B1(net2107),
    .Y(_1070_),
    .A1(_0128_),
    .A2(net1762));
 sg13g2_o21ai_1 _5409_ (.B1(_1062_),
    .Y(_1071_),
    .A1(_1069_),
    .A2(_1070_));
 sg13g2_a21oi_1 _5410_ (.A1(net2055),
    .A2(net966),
    .Y(_1072_),
    .B1(_1071_));
 sg13g2_a21o_1 _5411_ (.A2(_1053_),
    .A1(net2090),
    .B1(_1072_),
    .X(_0016_));
 sg13g2_or3_1 _5412_ (.A(_0129_),
    .B(net1758),
    .C(_1058_),
    .X(_1073_));
 sg13g2_nor2_2 _5413_ (.A(_0908_),
    .B(net1915),
    .Y(_1074_));
 sg13g2_nor2_1 _5414_ (.A(_0129_),
    .B(net2007),
    .Y(_1075_));
 sg13g2_a21oi_1 _5415_ (.A1(net1997),
    .A2(_1074_),
    .Y(_1076_),
    .B1(_1075_));
 sg13g2_a22oi_1 _5416_ (.Y(_1077_),
    .B1(_1076_),
    .B2(net2118),
    .A2(_1073_),
    .A1(net1736));
 sg13g2_o21ai_1 _5417_ (.B1(net2108),
    .Y(_1078_),
    .A1(_0129_),
    .A2(net1762));
 sg13g2_o21ai_1 _5418_ (.B1(_1062_),
    .Y(_1079_),
    .A1(_1077_),
    .A2(_1078_));
 sg13g2_a21oi_1 _5419_ (.A1(net2055),
    .A2(net948),
    .Y(_1080_),
    .B1(_1079_));
 sg13g2_a21o_1 _5420_ (.A2(_1053_),
    .A1(net2088),
    .B1(_1080_),
    .X(_0017_));
 sg13g2_or3_1 _5421_ (.A(_0130_),
    .B(net1758),
    .C(_1058_),
    .X(_1081_));
 sg13g2_nor2_1 _5422_ (.A(_0925_),
    .B(net1914),
    .Y(_1082_));
 sg13g2_nor2_1 _5423_ (.A(_0130_),
    .B(net2006),
    .Y(_1083_));
 sg13g2_a21oi_1 _5424_ (.A1(net1997),
    .A2(_1082_),
    .Y(_1084_),
    .B1(_1083_));
 sg13g2_a22oi_1 _5425_ (.Y(_1085_),
    .B1(_1084_),
    .B2(net2118),
    .A2(_1081_),
    .A1(net1736));
 sg13g2_o21ai_1 _5426_ (.B1(net2107),
    .Y(_1086_),
    .A1(_0130_),
    .A2(net1762));
 sg13g2_o21ai_1 _5427_ (.B1(_1062_),
    .Y(_1087_),
    .A1(_1085_),
    .A2(_1086_));
 sg13g2_a21oi_1 _5428_ (.A1(net2055),
    .A2(net911),
    .Y(_1088_),
    .B1(_1087_));
 sg13g2_a21o_1 _5429_ (.A2(_1053_),
    .A1(net2087),
    .B1(net912),
    .X(_0018_));
 sg13g2_nor2_1 _5430_ (.A(_0937_),
    .B(_1019_),
    .Y(_1089_));
 sg13g2_o21ai_1 _5431_ (.B1(net1740),
    .Y(_1090_),
    .A1(_0131_),
    .A2(net2008));
 sg13g2_a21oi_1 _5432_ (.A1(net1999),
    .A2(_1089_),
    .Y(_1091_),
    .B1(_1090_));
 sg13g2_nor2_1 _5433_ (.A(_0714_),
    .B(_0720_),
    .Y(_1092_));
 sg13g2_nand2_1 _5434_ (.Y(_1093_),
    .A(_0867_),
    .B(_1092_));
 sg13g2_and2_1 _5435_ (.A(_0131_),
    .B(_1093_),
    .X(_1094_));
 sg13g2_a221oi_1 _5436_ (.B2(_1094_),
    .C1(_1091_),
    .B1(net1749),
    .A1(_0132_),
    .Y(_1095_),
    .A2(net1755));
 sg13g2_nand4_1 _5437_ (.B(\debug_controller_inst.grid_out_valid ),
    .C(_0819_),
    .A(net2085),
    .Y(_1096_),
    .D(_0934_));
 sg13g2_and2_1 _5438_ (.A(net2275),
    .B(_1096_),
    .X(_1097_));
 sg13g2_o21ai_1 _5439_ (.B1(_1097_),
    .Y(_1098_),
    .A1(net2059),
    .A2(_1095_));
 sg13g2_a21o_1 _5440_ (.A2(net963),
    .A1(net2059),
    .B1(_1098_),
    .X(_1099_));
 sg13g2_o21ai_1 _5441_ (.B1(_1099_),
    .Y(_0019_),
    .A1(_3936_),
    .A2(_1096_));
 sg13g2_nor2_1 _5442_ (.A(_0950_),
    .B(net1915),
    .Y(_1100_));
 sg13g2_nand2_1 _5443_ (.Y(_1101_),
    .A(net1999),
    .B(_1100_));
 sg13g2_o21ai_1 _5444_ (.B1(_1101_),
    .Y(_1102_),
    .A1(_0133_),
    .A2(net2008));
 sg13g2_nor2_1 _5445_ (.A(_0869_),
    .B(_1093_),
    .Y(_1103_));
 sg13g2_a22oi_1 _5446_ (.Y(_1104_),
    .B1(net1749),
    .B2(net930),
    .A2(net1755),
    .A1(_0134_));
 sg13g2_o21ai_1 _5447_ (.B1(_1104_),
    .Y(_1105_),
    .A1(net1735),
    .A2(_1102_));
 sg13g2_o21ai_1 _5448_ (.B1(net2116),
    .Y(_1106_),
    .A1(_1103_),
    .A2(_1105_));
 sg13g2_nand2_1 _5449_ (.Y(_1107_),
    .A(net2060),
    .B(net930));
 sg13g2_nand3_1 _5450_ (.B(_1106_),
    .C(_1107_),
    .A(_1097_),
    .Y(_1108_));
 sg13g2_o21ai_1 _5451_ (.B1(net931),
    .Y(_0020_),
    .A1(_0949_),
    .A2(_1096_));
 sg13g2_nor2_1 _5452_ (.A(_0960_),
    .B(net1915),
    .Y(_1109_));
 sg13g2_nor3_1 _5453_ (.A(net2001),
    .B(_0960_),
    .C(net1915),
    .Y(_1110_));
 sg13g2_o21ai_1 _5454_ (.B1(net1740),
    .Y(_1111_),
    .A1(_0135_),
    .A2(net2008));
 sg13g2_a22oi_1 _5455_ (.Y(_1112_),
    .B1(net1747),
    .B2(_0135_),
    .A2(net1755),
    .A1(_0136_));
 sg13g2_o21ai_1 _5456_ (.B1(_1112_),
    .Y(_1113_),
    .A1(_1110_),
    .A2(_1111_));
 sg13g2_o21ai_1 _5457_ (.B1(net2116),
    .Y(_1114_),
    .A1(_1103_),
    .A2(_1113_));
 sg13g2_nand2_1 _5458_ (.Y(_1115_),
    .A(net2060),
    .B(net977));
 sg13g2_nand3_1 _5459_ (.B(_1114_),
    .C(_1115_),
    .A(_1097_),
    .Y(_1116_));
 sg13g2_o21ai_1 _5460_ (.B1(net978),
    .Y(_0021_),
    .A1(_0959_),
    .A2(_1096_));
 sg13g2_nor2_1 _5461_ (.A(_0969_),
    .B(net1915),
    .Y(_1117_));
 sg13g2_nor3_1 _5462_ (.A(net2001),
    .B(_0969_),
    .C(net1915),
    .Y(_1118_));
 sg13g2_o21ai_1 _5463_ (.B1(net1740),
    .Y(_1119_),
    .A1(_0137_),
    .A2(net2008));
 sg13g2_a22oi_1 _5464_ (.Y(_1120_),
    .B1(net1747),
    .B2(_0137_),
    .A2(net1755),
    .A1(_0138_));
 sg13g2_o21ai_1 _5465_ (.B1(_1120_),
    .Y(_1121_),
    .A1(_1118_),
    .A2(_1119_));
 sg13g2_o21ai_1 _5466_ (.B1(net2115),
    .Y(_1122_),
    .A1(_1103_),
    .A2(_1121_));
 sg13g2_nand2_1 _5467_ (.Y(_1123_),
    .A(net2059),
    .B(net985));
 sg13g2_nand3_1 _5468_ (.B(_1122_),
    .C(_1123_),
    .A(_1097_),
    .Y(_1124_));
 sg13g2_o21ai_1 _5469_ (.B1(net986),
    .Y(_0022_),
    .A1(_0968_),
    .A2(_1096_));
 sg13g2_nand3_1 _5470_ (.B(\debug_controller_inst.grid_out_addr[1] ),
    .C(\debug_controller_inst.grid_out_addr[0] ),
    .A(net2084),
    .Y(_1125_));
 sg13g2_nor2_2 _5471_ (.A(_0820_),
    .B(_1125_),
    .Y(_1126_));
 sg13g2_nor3_1 _5472_ (.A(net2000),
    .B(_0980_),
    .C(net1914),
    .Y(_1127_));
 sg13g2_o21ai_1 _5473_ (.B1(net1741),
    .Y(_1128_),
    .A1(_0139_),
    .A2(net2006));
 sg13g2_nor2_1 _5474_ (.A(_0714_),
    .B(_0718_),
    .Y(_1129_));
 sg13g2_nand2_2 _5475_ (.Y(_1130_),
    .A(net1728),
    .B(_1129_));
 sg13g2_and2_1 _5476_ (.A(_0139_),
    .B(net1746),
    .X(_1131_));
 sg13g2_a22oi_1 _5477_ (.Y(_1132_),
    .B1(_1130_),
    .B2(_1131_),
    .A2(net1752),
    .A1(net1046));
 sg13g2_o21ai_1 _5478_ (.B1(_1132_),
    .Y(_1133_),
    .A1(_1127_),
    .A2(_1128_));
 sg13g2_nand2_1 _5479_ (.Y(_1134_),
    .A(net2109),
    .B(_1133_));
 sg13g2_o21ai_1 _5480_ (.B1(net2274),
    .Y(_1135_),
    .A1(_0820_),
    .A2(_1125_));
 sg13g2_a21oi_1 _5481_ (.A1(net2056),
    .A2(net939),
    .Y(_1136_),
    .B1(_1135_));
 sg13g2_a22oi_1 _5482_ (.Y(_1137_),
    .B1(_1134_),
    .B2(_1136_),
    .A2(_1126_),
    .A1(net2092));
 sg13g2_inv_1 _5483_ (.Y(_0023_),
    .A(_1137_));
 sg13g2_nand3_1 _5484_ (.B(_0990_),
    .C(_1018_),
    .A(net1998),
    .Y(_1138_));
 sg13g2_o21ai_1 _5485_ (.B1(_1138_),
    .Y(_1139_),
    .A1(_0141_),
    .A2(net2006));
 sg13g2_nor2_1 _5486_ (.A(net1917),
    .B(_1130_),
    .Y(_1140_));
 sg13g2_a221oi_1 _5487_ (.B2(_0141_),
    .C1(_1140_),
    .B1(net1746),
    .A1(net898),
    .Y(_1141_),
    .A2(net1752));
 sg13g2_o21ai_1 _5488_ (.B1(_1141_),
    .Y(_1142_),
    .A1(net1733),
    .A2(_1139_));
 sg13g2_nand2_1 _5489_ (.Y(_1143_),
    .A(net2056),
    .B(net973));
 sg13g2_a21oi_1 _5490_ (.A1(net2109),
    .A2(_1142_),
    .Y(_1144_),
    .B1(_1135_));
 sg13g2_a22oi_1 _5491_ (.Y(_1145_),
    .B1(_1143_),
    .B2(_1144_),
    .A2(_1126_),
    .A1(net2090));
 sg13g2_inv_1 _5492_ (.Y(_0024_),
    .A(_1145_));
 sg13g2_nor2_1 _5493_ (.A(_0999_),
    .B(net1914),
    .Y(_1146_));
 sg13g2_o21ai_1 _5494_ (.B1(net1738),
    .Y(_1147_),
    .A1(_0143_),
    .A2(net2007));
 sg13g2_a21oi_1 _5495_ (.A1(net1999),
    .A2(_1146_),
    .Y(_1148_),
    .B1(_1147_));
 sg13g2_a22oi_1 _5496_ (.Y(_1149_),
    .B1(net1746),
    .B2(_0143_),
    .A2(net1752),
    .A1(_0144_));
 sg13g2_o21ai_1 _5497_ (.B1(_1149_),
    .Y(_1150_),
    .A1(net1917),
    .A2(_1130_));
 sg13g2_o21ai_1 _5498_ (.B1(net2108),
    .Y(_1151_),
    .A1(_1148_),
    .A2(_1150_));
 sg13g2_a21oi_1 _5499_ (.A1(net2056),
    .A2(net949),
    .Y(_1152_),
    .B1(_1135_));
 sg13g2_a22oi_1 _5500_ (.Y(_1153_),
    .B1(_1151_),
    .B2(_1152_),
    .A2(_1126_),
    .A1(net2088));
 sg13g2_inv_1 _5501_ (.Y(_0026_),
    .A(net950));
 sg13g2_nor2_1 _5502_ (.A(_1009_),
    .B(net1914),
    .Y(_1154_));
 sg13g2_o21ai_1 _5503_ (.B1(net1738),
    .Y(_1155_),
    .A1(_0145_),
    .A2(net2006));
 sg13g2_a21oi_1 _5504_ (.A1(net1997),
    .A2(_1154_),
    .Y(_1156_),
    .B1(_1155_));
 sg13g2_a22oi_1 _5505_ (.Y(_1157_),
    .B1(net1746),
    .B2(net953),
    .A2(net1752),
    .A1(_0146_));
 sg13g2_o21ai_1 _5506_ (.B1(_1157_),
    .Y(_1158_),
    .A1(net1917),
    .A2(_1130_));
 sg13g2_o21ai_1 _5507_ (.B1(net2109),
    .Y(_1159_),
    .A1(_1156_),
    .A2(_1158_));
 sg13g2_a21oi_1 _5508_ (.A1(net2056),
    .A2(net953),
    .Y(_1160_),
    .B1(_1135_));
 sg13g2_a22oi_1 _5509_ (.Y(_1161_),
    .B1(_1159_),
    .B2(_1160_),
    .A2(_1126_),
    .A1(net2086));
 sg13g2_inv_1 _5510_ (.Y(_0027_),
    .A(net954));
 sg13g2_and3_2 _5511_ (.X(_1162_),
    .A(net895),
    .B(\debug_controller_inst.grid_out_valid ),
    .C(_0531_));
 sg13g2_nand2_1 _5512_ (.Y(_1163_),
    .A(net2093),
    .B(_1162_));
 sg13g2_o21ai_1 _5513_ (.B1(net1739),
    .Y(_1164_),
    .A1(net989),
    .A2(net2005));
 sg13g2_a21oi_1 _5514_ (.A1(net2005),
    .A2(_0702_),
    .Y(_1165_),
    .B1(_1164_));
 sg13g2_nor3_2 _5515_ (.A(_0708_),
    .B(_0759_),
    .C(_0760_),
    .Y(_1166_));
 sg13g2_nand3_1 _5516_ (.B(_0765_),
    .C(_1166_),
    .A(_0521_),
    .Y(_1167_));
 sg13g2_a21oi_1 _5517_ (.A1(_0521_),
    .A2(net1916),
    .Y(_1168_),
    .B1(_4019_));
 sg13g2_a221oi_1 _5518_ (.B2(_1168_),
    .C1(_1165_),
    .B1(_1167_),
    .A1(net902),
    .Y(_1169_),
    .A2(net1756));
 sg13g2_nor2_1 _5519_ (.A(net2058),
    .B(_1169_),
    .Y(_1170_));
 sg13g2_nor2_2 _5520_ (.A(net2260),
    .B(_1162_),
    .Y(_1171_));
 sg13g2_o21ai_1 _5521_ (.B1(_1171_),
    .Y(_1172_),
    .A1(net2112),
    .A2(_4019_));
 sg13g2_o21ai_1 _5522_ (.B1(_1163_),
    .Y(_0028_),
    .A1(_1170_),
    .A2(_1172_));
 sg13g2_o21ai_1 _5523_ (.B1(net1739),
    .Y(_1173_),
    .A1(_0114_),
    .A2(net2005));
 sg13g2_a21o_1 _5524_ (.A2(_0785_),
    .A1(net2005),
    .B1(_1173_),
    .X(_1174_));
 sg13g2_or2_1 _5525_ (.X(_1175_),
    .B(_1167_),
    .A(net1916));
 sg13g2_a22oi_1 _5526_ (.Y(_1176_),
    .B1(net1748),
    .B2(net1023),
    .A2(net1756),
    .A1(_0113_));
 sg13g2_nand3_1 _5527_ (.B(_1175_),
    .C(_1176_),
    .A(_1174_),
    .Y(_1177_));
 sg13g2_o21ai_1 _5528_ (.B1(_1171_),
    .Y(_1178_),
    .A1(net2111),
    .A2(_4021_));
 sg13g2_a21oi_1 _5529_ (.A1(net2111),
    .A2(_1177_),
    .Y(_1179_),
    .B1(_1178_));
 sg13g2_a21o_1 _5530_ (.A2(_1162_),
    .A1(net2091),
    .B1(net1024),
    .X(_0029_));
 sg13g2_a21oi_1 _5531_ (.A1(_4023_),
    .A2(net2004),
    .Y(_1180_),
    .B1(net1734));
 sg13g2_o21ai_1 _5532_ (.B1(_1180_),
    .Y(_1181_),
    .A1(net2004),
    .A2(_0800_));
 sg13g2_a22oi_1 _5533_ (.Y(_1182_),
    .B1(net1748),
    .B2(net1017),
    .A2(net1756),
    .A1(_0115_));
 sg13g2_nand3_1 _5534_ (.B(_1181_),
    .C(_1182_),
    .A(_1175_),
    .Y(_1183_));
 sg13g2_o21ai_1 _5535_ (.B1(_1171_),
    .Y(_1184_),
    .A1(net2111),
    .A2(_4023_));
 sg13g2_a21oi_1 _5536_ (.A1(net2111),
    .A2(_1183_),
    .Y(_1185_),
    .B1(_1184_));
 sg13g2_a21o_1 _5537_ (.A2(_1162_),
    .A1(net2089),
    .B1(net1018),
    .X(_0030_));
 sg13g2_a21oi_1 _5538_ (.A1(_4025_),
    .A2(net2004),
    .Y(_1186_),
    .B1(net1734));
 sg13g2_o21ai_1 _5539_ (.B1(_1186_),
    .Y(_1187_),
    .A1(net2004),
    .A2(_0813_));
 sg13g2_a22oi_1 _5540_ (.Y(_1188_),
    .B1(net1748),
    .B2(net1020),
    .A2(net1756),
    .A1(_0117_));
 sg13g2_nand3_1 _5541_ (.B(_1187_),
    .C(_1188_),
    .A(_1175_),
    .Y(_1189_));
 sg13g2_o21ai_1 _5542_ (.B1(_1171_),
    .Y(_1190_),
    .A1(net2111),
    .A2(_4025_));
 sg13g2_a21oi_1 _5543_ (.A1(net2111),
    .A2(_1189_),
    .Y(_1191_),
    .B1(_1190_));
 sg13g2_a21o_1 _5544_ (.A2(_1162_),
    .A1(net2087),
    .B1(net1021),
    .X(_0031_));
 sg13g2_nand2b_2 _5545_ (.Y(_1192_),
    .B(\debug_controller_inst.grid_out_valid ),
    .A_N(_0819_));
 sg13g2_inv_1 _5546_ (.Y(_1193_),
    .A(_1192_));
 sg13g2_nor3_2 _5547_ (.A(net2084),
    .B(_0821_),
    .C(_1192_),
    .Y(_1194_));
 sg13g2_nor2_1 _5548_ (.A(net2003),
    .B(_0862_),
    .Y(_1195_));
 sg13g2_o21ai_1 _5549_ (.B1(net1740),
    .Y(_1196_),
    .A1(_0132_),
    .A2(_0540_));
 sg13g2_nand3_1 _5550_ (.B(_0866_),
    .C(_1166_),
    .A(net1775),
    .Y(_1197_));
 sg13g2_a21oi_1 _5551_ (.A1(net1775),
    .A2(net1916),
    .Y(_1198_),
    .B1(_4031_));
 sg13g2_a22oi_1 _5552_ (.Y(_1199_),
    .B1(_1197_),
    .B2(_1198_),
    .A2(net1755),
    .A1(_0131_));
 sg13g2_o21ai_1 _5553_ (.B1(_1199_),
    .Y(_1200_),
    .A1(_1195_),
    .A2(_1196_));
 sg13g2_nor2_2 _5554_ (.A(net2260),
    .B(_1194_),
    .Y(_1201_));
 sg13g2_o21ai_1 _5555_ (.B1(_1201_),
    .Y(_1202_),
    .A1(net2115),
    .A2(_4031_));
 sg13g2_a21oi_1 _5556_ (.A1(net2115),
    .A2(_1200_),
    .Y(_1203_),
    .B1(_1202_));
 sg13g2_a21o_1 _5557_ (.A2(_1194_),
    .A1(net2093),
    .B1(_1203_),
    .X(_0032_));
 sg13g2_a21oi_1 _5558_ (.A1(_0496_),
    .A2(net2002),
    .Y(_1204_),
    .B1(net1735));
 sg13g2_o21ai_1 _5559_ (.B1(_1204_),
    .Y(_1205_),
    .A1(net2003),
    .A2(_0890_));
 sg13g2_or2_1 _5560_ (.X(_1206_),
    .B(_1197_),
    .A(net1916));
 sg13g2_a22oi_1 _5561_ (.Y(_1207_),
    .B1(net1747),
    .B2(net1033),
    .A2(net1755),
    .A1(_0133_));
 sg13g2_nand3_1 _5562_ (.B(_1206_),
    .C(_1207_),
    .A(_1205_),
    .Y(_1208_));
 sg13g2_o21ai_1 _5563_ (.B1(_1201_),
    .Y(_1209_),
    .A1(net2115),
    .A2(_0496_));
 sg13g2_a21oi_1 _5564_ (.A1(net2116),
    .A2(_1208_),
    .Y(_1210_),
    .B1(_1209_));
 sg13g2_a21o_1 _5565_ (.A2(_1194_),
    .A1(net2091),
    .B1(_1210_),
    .X(_0033_));
 sg13g2_a21oi_1 _5566_ (.A1(_0497_),
    .A2(net2002),
    .Y(_1211_),
    .B1(net1735));
 sg13g2_o21ai_1 _5567_ (.B1(_1211_),
    .Y(_1212_),
    .A1(net2003),
    .A2(_0908_));
 sg13g2_a22oi_1 _5568_ (.Y(_1213_),
    .B1(net1747),
    .B2(net1019),
    .A2(net1755),
    .A1(_0135_));
 sg13g2_nand3_1 _5569_ (.B(_1212_),
    .C(_1213_),
    .A(_1206_),
    .Y(_1214_));
 sg13g2_o21ai_1 _5570_ (.B1(_1201_),
    .Y(_1215_),
    .A1(net2115),
    .A2(_0497_));
 sg13g2_a21oi_1 _5571_ (.A1(net2115),
    .A2(_1214_),
    .Y(_1216_),
    .B1(_1215_));
 sg13g2_a21o_1 _5572_ (.A2(_1194_),
    .A1(net2089),
    .B1(_1216_),
    .X(_0034_));
 sg13g2_a21oi_1 _5573_ (.A1(_0498_),
    .A2(net2002),
    .Y(_1217_),
    .B1(net1735));
 sg13g2_o21ai_1 _5574_ (.B1(_1217_),
    .Y(_1218_),
    .A1(net2003),
    .A2(_0925_));
 sg13g2_a22oi_1 _5575_ (.Y(_1219_),
    .B1(net1747),
    .B2(net1029),
    .A2(net1755),
    .A1(_0137_));
 sg13g2_nand3_1 _5576_ (.B(_1218_),
    .C(_1219_),
    .A(_1206_),
    .Y(_1220_));
 sg13g2_o21ai_1 _5577_ (.B1(_1201_),
    .Y(_1221_),
    .A1(net2115),
    .A2(_0498_));
 sg13g2_a21oi_1 _5578_ (.A1(net2115),
    .A2(_1220_),
    .Y(_1222_),
    .B1(_1221_));
 sg13g2_a21o_1 _5579_ (.A2(_1194_),
    .A1(net2087),
    .B1(_1222_),
    .X(_0035_));
 sg13g2_nand2_2 _5580_ (.Y(_1223_),
    .A(_0935_),
    .B(_1193_));
 sg13g2_or2_1 _5581_ (.X(_1224_),
    .B(_1223_),
    .A(_0933_));
 sg13g2_a21oi_1 _5582_ (.A1(_0499_),
    .A2(net2004),
    .Y(_1225_),
    .B1(_3940_));
 sg13g2_o21ai_1 _5583_ (.B1(_1225_),
    .Y(_1226_),
    .A1(net2004),
    .A2(_0937_));
 sg13g2_and2_1 _5584_ (.A(_0940_),
    .B(_1166_),
    .X(_1227_));
 sg13g2_nor3_1 _5585_ (.A(net2121),
    .B(_0499_),
    .C(_1227_),
    .Y(_1228_));
 sg13g2_nor2_1 _5586_ (.A(net1760),
    .B(_1228_),
    .Y(_1229_));
 sg13g2_a221oi_1 _5587_ (.B2(_1229_),
    .C1(net2057),
    .B1(_1226_),
    .A1(_0499_),
    .Y(_1230_),
    .A2(net1760));
 sg13g2_a21oi_2 _5588_ (.B1(net2260),
    .Y(_1231_),
    .A2(_1193_),
    .A1(_0935_));
 sg13g2_o21ai_1 _5589_ (.B1(_1231_),
    .Y(_1232_),
    .A1(net2113),
    .A2(_0499_));
 sg13g2_o21ai_1 _5590_ (.B1(_1224_),
    .Y(_0037_),
    .A1(_1230_),
    .A2(_1232_));
 sg13g2_or3_1 _5591_ (.A(_0148_),
    .B(net1760),
    .C(_1227_),
    .X(_1233_));
 sg13g2_mux2_1 _5592_ (.A0(_0148_),
    .A1(_0950_),
    .S(net2005),
    .X(_1234_));
 sg13g2_a22oi_1 _5593_ (.Y(_1235_),
    .B1(_1234_),
    .B2(net2121),
    .A2(_1233_),
    .A1(net1734));
 sg13g2_o21ai_1 _5594_ (.B1(net2112),
    .Y(_1236_),
    .A1(net933),
    .A2(net1763));
 sg13g2_o21ai_1 _5595_ (.B1(_1231_),
    .Y(_1237_),
    .A1(_1235_),
    .A2(_1236_));
 sg13g2_a21o_1 _5596_ (.A2(net933),
    .A1(net2058),
    .B1(_1237_),
    .X(_1238_));
 sg13g2_o21ai_1 _5597_ (.B1(_1238_),
    .Y(_0038_),
    .A1(_0949_),
    .A2(_1223_));
 sg13g2_or3_1 _5598_ (.A(_0149_),
    .B(net1759),
    .C(_1227_),
    .X(_1239_));
 sg13g2_mux2_1 _5599_ (.A0(_0149_),
    .A1(_0960_),
    .S(net2005),
    .X(_1240_));
 sg13g2_a22oi_1 _5600_ (.Y(_1241_),
    .B1(_1240_),
    .B2(net2121),
    .A2(_1239_),
    .A1(net1734));
 sg13g2_o21ai_1 _5601_ (.B1(net2112),
    .Y(_1242_),
    .A1(net917),
    .A2(net1763));
 sg13g2_o21ai_1 _5602_ (.B1(_1231_),
    .Y(_1243_),
    .A1(_1241_),
    .A2(_1242_));
 sg13g2_a21o_1 _5603_ (.A2(net917),
    .A1(net2058),
    .B1(_1243_),
    .X(_1244_));
 sg13g2_o21ai_1 _5604_ (.B1(_1244_),
    .Y(_0039_),
    .A1(_0959_),
    .A2(_1223_));
 sg13g2_or3_1 _5605_ (.A(_0150_),
    .B(net1759),
    .C(_1227_),
    .X(_1245_));
 sg13g2_mux2_1 _5606_ (.A0(_0150_),
    .A1(_0969_),
    .S(net2005),
    .X(_1246_));
 sg13g2_a22oi_1 _5607_ (.Y(_1247_),
    .B1(_1246_),
    .B2(net2121),
    .A2(_1245_),
    .A1(net1734));
 sg13g2_o21ai_1 _5608_ (.B1(net2113),
    .Y(_1248_),
    .A1(net922),
    .A2(net1763));
 sg13g2_o21ai_1 _5609_ (.B1(_1231_),
    .Y(_1249_),
    .A1(_1247_),
    .A2(_1248_));
 sg13g2_a21o_1 _5610_ (.A2(net922),
    .A1(net2058),
    .B1(_1249_),
    .X(_1250_));
 sg13g2_o21ai_1 _5611_ (.B1(_1250_),
    .Y(_0040_),
    .A1(_0968_),
    .A2(_1223_));
 sg13g2_nor3_2 _5612_ (.A(net2084),
    .B(_0977_),
    .C(_1192_),
    .Y(_1251_));
 sg13g2_nor2_1 _5613_ (.A(net2002),
    .B(_0980_),
    .Y(_1252_));
 sg13g2_o21ai_1 _5614_ (.B1(net1740),
    .Y(_1253_),
    .A1(_0151_),
    .A2(_0540_));
 sg13g2_nand3_1 _5615_ (.B(_0983_),
    .C(_1166_),
    .A(net1775),
    .Y(_1254_));
 sg13g2_a21oi_1 _5616_ (.A1(net1775),
    .A2(net1916),
    .Y(_1255_),
    .B1(_0500_));
 sg13g2_a22oi_1 _5617_ (.Y(_1256_),
    .B1(_1254_),
    .B2(_1255_),
    .A2(net1754),
    .A1(_0152_));
 sg13g2_o21ai_1 _5618_ (.B1(_1256_),
    .Y(_1257_),
    .A1(_1252_),
    .A2(_1253_));
 sg13g2_nor2_2 _5619_ (.A(net2260),
    .B(_1251_),
    .Y(_1258_));
 sg13g2_o21ai_1 _5620_ (.B1(_1258_),
    .Y(_1259_),
    .A1(net2117),
    .A2(_0500_));
 sg13g2_a21oi_1 _5621_ (.A1(net2114),
    .A2(_1257_),
    .Y(_1260_),
    .B1(_1259_));
 sg13g2_a21o_1 _5622_ (.A2(_1251_),
    .A1(net2093),
    .B1(_1260_),
    .X(_0041_));
 sg13g2_nand2_1 _5623_ (.Y(_1261_),
    .A(net2091),
    .B(_1251_));
 sg13g2_o21ai_1 _5624_ (.B1(net1740),
    .Y(_1262_),
    .A1(_0153_),
    .A2(_0540_));
 sg13g2_a21oi_1 _5625_ (.A1(net2005),
    .A2(_0990_),
    .Y(_1263_),
    .B1(_1262_));
 sg13g2_or2_1 _5626_ (.X(_1264_),
    .B(_1254_),
    .A(net1916));
 sg13g2_a22oi_1 _5627_ (.Y(_1265_),
    .B1(net1747),
    .B2(_0153_),
    .A2(net1754),
    .A1(_0154_));
 sg13g2_nand2_1 _5628_ (.Y(_1266_),
    .A(_1264_),
    .B(_1265_));
 sg13g2_o21ai_1 _5629_ (.B1(net2117),
    .Y(_1267_),
    .A1(_1263_),
    .A2(_1266_));
 sg13g2_nand2_1 _5630_ (.Y(_1268_),
    .A(net2059),
    .B(_0153_));
 sg13g2_nand3_1 _5631_ (.B(_1267_),
    .C(_1268_),
    .A(_1258_),
    .Y(_1269_));
 sg13g2_nand2_1 _5632_ (.Y(_0042_),
    .A(_1261_),
    .B(_1269_));
 sg13g2_a21oi_1 _5633_ (.A1(_0501_),
    .A2(net2002),
    .Y(_1270_),
    .B1(net1734));
 sg13g2_o21ai_1 _5634_ (.B1(_1270_),
    .Y(_1271_),
    .A1(net2002),
    .A2(_0999_));
 sg13g2_a22oi_1 _5635_ (.Y(_1272_),
    .B1(net1747),
    .B2(_0155_),
    .A2(net1754),
    .A1(net909));
 sg13g2_nand3_1 _5636_ (.B(_1271_),
    .C(_1272_),
    .A(_1264_),
    .Y(_1273_));
 sg13g2_o21ai_1 _5637_ (.B1(_1258_),
    .Y(_1274_),
    .A1(net2117),
    .A2(_0501_));
 sg13g2_a21oi_1 _5638_ (.A1(net2114),
    .A2(_1273_),
    .Y(_1275_),
    .B1(_1274_));
 sg13g2_a21o_1 _5639_ (.A2(_1251_),
    .A1(net2089),
    .B1(_1275_),
    .X(_0043_));
 sg13g2_a21oi_1 _5640_ (.A1(_0502_),
    .A2(net2002),
    .Y(_1276_),
    .B1(net1734));
 sg13g2_o21ai_1 _5641_ (.B1(_1276_),
    .Y(_1277_),
    .A1(net2002),
    .A2(_1009_));
 sg13g2_a22oi_1 _5642_ (.Y(_1278_),
    .B1(net1747),
    .B2(net1036),
    .A2(net1754),
    .A1(_0158_));
 sg13g2_nand3_1 _5643_ (.B(_1277_),
    .C(_1278_),
    .A(_1264_),
    .Y(_1279_));
 sg13g2_o21ai_1 _5644_ (.B1(_1258_),
    .Y(_1280_),
    .A1(net2114),
    .A2(_0502_));
 sg13g2_a21oi_1 _5645_ (.A1(net2114),
    .A2(_1279_),
    .Y(_1281_),
    .B1(_1280_));
 sg13g2_a21o_1 _5646_ (.A2(_1251_),
    .A1(net2086),
    .B1(_1281_),
    .X(_0044_));
 sg13g2_nand2_1 _5647_ (.Y(_1282_),
    .A(net2001),
    .B(net1740));
 sg13g2_a21oi_1 _5648_ (.A1(_0702_),
    .A2(_1018_),
    .Y(_1283_),
    .B1(net1726));
 sg13g2_a21oi_2 _5649_ (.B1(net1776),
    .Y(_1284_),
    .A2(net1738),
    .A1(net1998));
 sg13g2_and2_1 _5650_ (.A(_1022_),
    .B(_1166_),
    .X(_1285_));
 sg13g2_nand2_1 _5651_ (.Y(_1286_),
    .A(net1916),
    .B(_1284_));
 sg13g2_o21ai_1 _5652_ (.B1(_1284_),
    .Y(_1287_),
    .A1(net1917),
    .A2(_1285_));
 sg13g2_a221oi_1 _5653_ (.B2(net881),
    .C1(_1283_),
    .B1(_1287_),
    .A1(_0119_),
    .Y(_1288_),
    .A2(net1751));
 sg13g2_nand2b_1 _5654_ (.Y(_1289_),
    .B(net2105),
    .A_N(_1288_));
 sg13g2_nor2_2 _5655_ (.A(_1016_),
    .B(_1192_),
    .Y(_1290_));
 sg13g2_o21ai_1 _5656_ (.B1(net2269),
    .Y(_1291_),
    .A1(_1016_),
    .A2(_1192_));
 sg13g2_a21oi_1 _5657_ (.A1(net2054),
    .A2(net881),
    .Y(_1292_),
    .B1(_1291_));
 sg13g2_a22oi_1 _5658_ (.Y(_1293_),
    .B1(_1292_),
    .B2(_1289_),
    .A2(_1290_),
    .A1(net2092));
 sg13g2_inv_1 _5659_ (.Y(_0045_),
    .A(net882));
 sg13g2_and2_1 _5660_ (.A(_0895_),
    .B(_1285_),
    .X(_1294_));
 sg13g2_a221oi_1 _5661_ (.B2(net878),
    .C1(_1294_),
    .B1(net1725),
    .A1(net1045),
    .Y(_1295_),
    .A2(net1753));
 sg13g2_o21ai_1 _5662_ (.B1(_1295_),
    .Y(_1296_),
    .A1(_1031_),
    .A2(net1726));
 sg13g2_nand2_1 _5663_ (.Y(_1297_),
    .A(net2054),
    .B(net878));
 sg13g2_a21oi_1 _5664_ (.A1(net2106),
    .A2(_1296_),
    .Y(_1298_),
    .B1(_1291_));
 sg13g2_a22oi_1 _5665_ (.Y(_1299_),
    .B1(_1297_),
    .B2(_1298_),
    .A2(_1290_),
    .A1(net2090));
 sg13g2_inv_1 _5666_ (.Y(_0046_),
    .A(_1299_));
 sg13g2_a221oi_1 _5667_ (.B2(net869),
    .C1(_1294_),
    .B1(net1725),
    .A1(_0123_),
    .Y(_1300_),
    .A2(net1751));
 sg13g2_o21ai_1 _5668_ (.B1(_1300_),
    .Y(_1301_),
    .A1(_1039_),
    .A2(net1726));
 sg13g2_nand2_1 _5669_ (.Y(_1302_),
    .A(net2054),
    .B(net869));
 sg13g2_a21oi_1 _5670_ (.A1(net2106),
    .A2(_1301_),
    .Y(_1303_),
    .B1(_1291_));
 sg13g2_a22oi_1 _5671_ (.Y(_1304_),
    .B1(_1302_),
    .B2(_1303_),
    .A2(_1290_),
    .A1(net2088));
 sg13g2_inv_1 _5672_ (.Y(_0048_),
    .A(net870));
 sg13g2_a22oi_1 _5673_ (.Y(_1305_),
    .B1(net1725),
    .B2(_0126_),
    .A2(net1751),
    .A1(net891));
 sg13g2_o21ai_1 _5674_ (.B1(net892),
    .Y(_1306_),
    .A1(_1046_),
    .A2(net1726));
 sg13g2_o21ai_1 _5675_ (.B1(net2105),
    .Y(_1307_),
    .A1(_1294_),
    .A2(_1306_));
 sg13g2_a21oi_1 _5676_ (.A1(net2054),
    .A2(_0126_),
    .Y(_1308_),
    .B1(_1291_));
 sg13g2_a22oi_1 _5677_ (.Y(_1309_),
    .B1(_1307_),
    .B2(_1308_),
    .A2(_1290_),
    .A1(net2086));
 sg13g2_inv_1 _5678_ (.Y(_0049_),
    .A(net893));
 sg13g2_nor2_2 _5679_ (.A(_1052_),
    .B(_1192_),
    .Y(_1310_));
 sg13g2_nand2_1 _5680_ (.Y(_1311_),
    .A(net2092),
    .B(_1310_));
 sg13g2_and2_1 _5681_ (.A(_1057_),
    .B(_1166_),
    .X(_1312_));
 sg13g2_o21ai_1 _5682_ (.B1(_1284_),
    .Y(_1313_),
    .A1(net1917),
    .A2(_1312_));
 sg13g2_a22oi_1 _5683_ (.Y(_1314_),
    .B1(_1313_),
    .B2(net980),
    .A2(net1752),
    .A1(_0139_));
 sg13g2_o21ai_1 _5684_ (.B1(_1314_),
    .Y(_1315_),
    .A1(_1054_),
    .A2(net1726));
 sg13g2_o21ai_1 _5685_ (.B1(net2274),
    .Y(_1316_),
    .A1(_1052_),
    .A2(_1192_));
 sg13g2_mux2_1 _5686_ (.A0(net980),
    .A1(_1315_),
    .S(net2109),
    .X(_1317_));
 sg13g2_o21ai_1 _5687_ (.B1(_1311_),
    .Y(_0050_),
    .A1(_1316_),
    .A2(_1317_));
 sg13g2_nand2_1 _5688_ (.Y(_1318_),
    .A(net2091),
    .B(_1310_));
 sg13g2_and2_1 _5689_ (.A(_0895_),
    .B(_1312_),
    .X(_1319_));
 sg13g2_a221oi_1 _5690_ (.B2(net898),
    .C1(_1319_),
    .B1(net1725),
    .A1(_0141_),
    .Y(_1320_),
    .A2(net1753));
 sg13g2_o21ai_1 _5691_ (.B1(_1320_),
    .Y(_1321_),
    .A1(_1066_),
    .A2(net1726));
 sg13g2_mux2_1 _5692_ (.A0(net898),
    .A1(_1321_),
    .S(net2108),
    .X(_1322_));
 sg13g2_o21ai_1 _5693_ (.B1(_1318_),
    .Y(_0051_),
    .A1(_1316_),
    .A2(_1322_));
 sg13g2_nand2_1 _5694_ (.Y(_1323_),
    .A(net2089),
    .B(_1310_));
 sg13g2_a221oi_1 _5695_ (.B2(net970),
    .C1(_1319_),
    .B1(net1725),
    .A1(_0143_),
    .Y(_1324_),
    .A2(net1752));
 sg13g2_o21ai_1 _5696_ (.B1(_1324_),
    .Y(_1325_),
    .A1(_1074_),
    .A2(net1726));
 sg13g2_mux2_1 _5697_ (.A0(net970),
    .A1(_1325_),
    .S(net2108),
    .X(_1326_));
 sg13g2_o21ai_1 _5698_ (.B1(_1323_),
    .Y(_0052_),
    .A1(_1316_),
    .A2(net971));
 sg13g2_a221oi_1 _5699_ (.B2(net946),
    .C1(_1319_),
    .B1(net1725),
    .A1(_0145_),
    .Y(_1327_),
    .A2(net1753));
 sg13g2_o21ai_1 _5700_ (.B1(_1327_),
    .Y(_1328_),
    .A1(_1082_),
    .A2(net1726));
 sg13g2_nand2_1 _5701_ (.Y(_1329_),
    .A(net2056),
    .B(net946));
 sg13g2_a21oi_1 _5702_ (.A1(net2108),
    .A2(_1328_),
    .Y(_1330_),
    .B1(_1316_));
 sg13g2_a22oi_1 _5703_ (.Y(_1331_),
    .B1(_1329_),
    .B2(_1330_),
    .A2(_1310_),
    .A1(net2087));
 sg13g2_inv_1 _5704_ (.Y(_0053_),
    .A(net947));
 sg13g2_and2_1 _5705_ (.A(_1092_),
    .B(_1166_),
    .X(_1332_));
 sg13g2_o21ai_1 _5706_ (.B1(_1284_),
    .Y(_1333_),
    .A1(net1916),
    .A2(_1332_));
 sg13g2_a22oi_1 _5707_ (.Y(_1334_),
    .B1(_1333_),
    .B2(net1016),
    .A2(net1754),
    .A1(_0151_));
 sg13g2_o21ai_1 _5708_ (.B1(_1334_),
    .Y(_1335_),
    .A1(_1089_),
    .A2(net1727));
 sg13g2_nand3_1 _5709_ (.B(_0934_),
    .C(_1193_),
    .A(net2085),
    .Y(_1336_));
 sg13g2_and2_1 _5710_ (.A(net2275),
    .B(_1336_),
    .X(_1337_));
 sg13g2_nor2b_1 _5711_ (.A(net2114),
    .B_N(net1016),
    .Y(_1338_));
 sg13g2_a21oi_1 _5712_ (.A1(net2114),
    .A2(_1335_),
    .Y(_1339_),
    .B1(_1338_));
 sg13g2_nand2_1 _5713_ (.Y(_1340_),
    .A(_1337_),
    .B(_1339_));
 sg13g2_o21ai_1 _5714_ (.B1(_1340_),
    .Y(_0054_),
    .A1(_0933_),
    .A2(_1336_));
 sg13g2_and2_1 _5715_ (.A(_0895_),
    .B(_1332_),
    .X(_1341_));
 sg13g2_a221oi_1 _5716_ (.B2(net1008),
    .C1(_1341_),
    .B1(_1286_),
    .A1(_0153_),
    .Y(_1342_),
    .A2(net1754));
 sg13g2_o21ai_1 _5717_ (.B1(_1342_),
    .Y(_1343_),
    .A1(_1100_),
    .A2(net1727));
 sg13g2_nor2b_1 _5718_ (.A(net2116),
    .B_N(net1008),
    .Y(_1344_));
 sg13g2_a21oi_1 _5719_ (.A1(net2116),
    .A2(_1343_),
    .Y(_1345_),
    .B1(_1344_));
 sg13g2_nand2_1 _5720_ (.Y(_1346_),
    .A(_1337_),
    .B(_1345_));
 sg13g2_o21ai_1 _5721_ (.B1(_1346_),
    .Y(_0055_),
    .A1(_0949_),
    .A2(_1336_));
 sg13g2_a22oi_1 _5722_ (.Y(_1347_),
    .B1(net1725),
    .B2(net909),
    .A2(net1754),
    .A1(_0155_));
 sg13g2_o21ai_1 _5723_ (.B1(_1347_),
    .Y(_1348_),
    .A1(_1109_),
    .A2(net1727));
 sg13g2_o21ai_1 _5724_ (.B1(net2114),
    .Y(_1349_),
    .A1(_1341_),
    .A2(_1348_));
 sg13g2_nand2_1 _5725_ (.Y(_1350_),
    .A(net2059),
    .B(net909));
 sg13g2_nand3_1 _5726_ (.B(_1349_),
    .C(_1350_),
    .A(_1337_),
    .Y(_1351_));
 sg13g2_o21ai_1 _5727_ (.B1(_1351_),
    .Y(_0056_),
    .A1(_0959_),
    .A2(_1336_));
 sg13g2_a22oi_1 _5728_ (.Y(_1352_),
    .B1(net1725),
    .B2(_0158_),
    .A2(net1754),
    .A1(_0157_));
 sg13g2_o21ai_1 _5729_ (.B1(_1352_),
    .Y(_1353_),
    .A1(_1117_),
    .A2(net1727));
 sg13g2_o21ai_1 _5730_ (.B1(net2114),
    .Y(_1354_),
    .A1(_1341_),
    .A2(_1353_));
 sg13g2_nand2_1 _5731_ (.Y(_1355_),
    .A(net2059),
    .B(net974));
 sg13g2_nand3_1 _5732_ (.B(_1354_),
    .C(_1355_),
    .A(_1337_),
    .Y(_1356_));
 sg13g2_o21ai_1 _5733_ (.B1(net975),
    .Y(_0057_),
    .A1(_0968_),
    .A2(_1336_));
 sg13g2_nor2_2 _5734_ (.A(_1125_),
    .B(_1192_),
    .Y(_1357_));
 sg13g2_nor3_1 _5735_ (.A(net1997),
    .B(_0980_),
    .C(net1914),
    .Y(_1358_));
 sg13g2_o21ai_1 _5736_ (.B1(net2118),
    .Y(_1359_),
    .A1(_0159_),
    .A2(net2000));
 sg13g2_and2_1 _5737_ (.A(_1129_),
    .B(_1166_),
    .X(_1360_));
 sg13g2_nor3_1 _5738_ (.A(net2118),
    .B(_0503_),
    .C(_1360_),
    .Y(_1361_));
 sg13g2_nor2_1 _5739_ (.A(net1761),
    .B(_1361_),
    .Y(_1362_));
 sg13g2_o21ai_1 _5740_ (.B1(_1362_),
    .Y(_1363_),
    .A1(_1358_),
    .A2(_1359_));
 sg13g2_a21oi_1 _5741_ (.A1(_0503_),
    .A2(net1758),
    .Y(_1364_),
    .B1(net2055));
 sg13g2_nor2_2 _5742_ (.A(net2258),
    .B(_1357_),
    .Y(_1365_));
 sg13g2_o21ai_1 _5743_ (.B1(_1365_),
    .Y(_1366_),
    .A1(net2108),
    .A2(_0503_));
 sg13g2_a21oi_1 _5744_ (.A1(_1363_),
    .A2(_1364_),
    .Y(_1367_),
    .B1(_1366_));
 sg13g2_a21o_1 _5745_ (.A2(_1357_),
    .A1(net2092),
    .B1(_1367_),
    .X(_0059_));
 sg13g2_or3_1 _5746_ (.A(_0160_),
    .B(net1758),
    .C(_1360_),
    .X(_1368_));
 sg13g2_nand3_1 _5747_ (.B(_0990_),
    .C(_1018_),
    .A(net2001),
    .Y(_1369_));
 sg13g2_o21ai_1 _5748_ (.B1(net2118),
    .Y(_1370_),
    .A1(_0160_),
    .A2(net2000));
 sg13g2_inv_1 _5749_ (.Y(_1371_),
    .A(_1370_));
 sg13g2_a22oi_1 _5750_ (.Y(_1372_),
    .B1(_1369_),
    .B2(_1371_),
    .A2(_1368_),
    .A1(net1733));
 sg13g2_o21ai_1 _5751_ (.B1(net2107),
    .Y(_1373_),
    .A1(_0160_),
    .A2(net1762));
 sg13g2_o21ai_1 _5752_ (.B1(_1365_),
    .Y(_1374_),
    .A1(_1372_),
    .A2(_1373_));
 sg13g2_a21oi_1 _5753_ (.A1(net2055),
    .A2(net961),
    .Y(_1375_),
    .B1(_1374_));
 sg13g2_a21o_1 _5754_ (.A2(_1357_),
    .A1(net2090),
    .B1(_1375_),
    .X(_0060_));
 sg13g2_or3_1 _5755_ (.A(_0161_),
    .B(net1758),
    .C(_1360_),
    .X(_1376_));
 sg13g2_nor2_1 _5756_ (.A(_0161_),
    .B(net2000),
    .Y(_1377_));
 sg13g2_a21oi_1 _5757_ (.A1(net2000),
    .A2(_1146_),
    .Y(_1378_),
    .B1(_1377_));
 sg13g2_a22oi_1 _5758_ (.Y(_1379_),
    .B1(_1378_),
    .B2(net2119),
    .A2(_1376_),
    .A1(net1733));
 sg13g2_o21ai_1 _5759_ (.B1(net2107),
    .Y(_1380_),
    .A1(_0161_),
    .A2(net1762));
 sg13g2_o21ai_1 _5760_ (.B1(_1365_),
    .Y(_1381_),
    .A1(_1379_),
    .A2(_1380_));
 sg13g2_a21oi_1 _5761_ (.A1(net2055),
    .A2(net958),
    .Y(_1382_),
    .B1(_1381_));
 sg13g2_a21o_1 _5762_ (.A2(_1357_),
    .A1(net2088),
    .B1(_1382_),
    .X(_0061_));
 sg13g2_or3_1 _5763_ (.A(_0162_),
    .B(net1758),
    .C(_1360_),
    .X(_1383_));
 sg13g2_nor2_1 _5764_ (.A(_0162_),
    .B(net2000),
    .Y(_1384_));
 sg13g2_a21oi_1 _5765_ (.A1(net2000),
    .A2(_1154_),
    .Y(_1385_),
    .B1(_1384_));
 sg13g2_a22oi_1 _5766_ (.Y(_1386_),
    .B1(_1385_),
    .B2(net2119),
    .A2(_1383_),
    .A1(net1733));
 sg13g2_o21ai_1 _5767_ (.B1(net2107),
    .Y(_1387_),
    .A1(_0162_),
    .A2(net1762));
 sg13g2_o21ai_1 _5768_ (.B1(_1365_),
    .Y(_1388_),
    .A1(_1386_),
    .A2(_1387_));
 sg13g2_a21oi_1 _5769_ (.A1(net2056),
    .A2(net925),
    .Y(_1389_),
    .B1(_1388_));
 sg13g2_a21o_1 _5770_ (.A2(_1357_),
    .A1(net2086),
    .B1(net926),
    .X(_0062_));
 sg13g2_nor2_1 _5771_ (.A(net2196),
    .B(net2036),
    .Y(_1390_));
 sg13g2_nor2_2 _5772_ (.A(net2050),
    .B(net2193),
    .Y(_1391_));
 sg13g2_nand2_2 _5773_ (.Y(_1392_),
    .A(net2175),
    .B(net2043));
 sg13g2_nor2_2 _5774_ (.A(net2029),
    .B(net1902),
    .Y(_1393_));
 sg13g2_nand2_1 _5775_ (.Y(_1394_),
    .A(net2212),
    .B(net1911));
 sg13g2_nor2_2 _5776_ (.A(net2051),
    .B(net2162),
    .Y(_1395_));
 sg13g2_nand2_1 _5777_ (.Y(_1396_),
    .A(net2157),
    .B(_3995_));
 sg13g2_nor2b_1 _5778_ (.A(net896),
    .B_N(net883),
    .Y(_1397_));
 sg13g2_and2_2 _5779_ (.A(net2152),
    .B(\draw_game_inst.board_y[6] ),
    .X(_1398_));
 sg13g2_nand4_1 _5780_ (.B(net1899),
    .C(_1397_),
    .A(_1393_),
    .Y(_0068_),
    .D(_1398_));
 sg13g2_nor2_1 _5781_ (.A(net2136),
    .B(net2140),
    .Y(_1399_));
 sg13g2_nand2_2 _5782_ (.Y(_1400_),
    .A(net2024),
    .B(net2022));
 sg13g2_nor2_2 _5783_ (.A(net2026),
    .B(net2023),
    .Y(_1401_));
 sg13g2_nand2_2 _5784_ (.Y(_1402_),
    .A(net2135),
    .B(net2144));
 sg13g2_nand3b_1 _5785_ (.B(net2125),
    .C(net945),
    .Y(_1403_),
    .A_N(net1007));
 sg13g2_a21oi_1 _5786_ (.A1(net2129),
    .A2(_1401_),
    .Y(_1404_),
    .B1(_1403_));
 sg13g2_o21ai_1 _5787_ (.B1(_1404_),
    .Y(_0067_),
    .A1(net2129),
    .A2(net1892));
 sg13g2_and2_1 _5788_ (.A(net2277),
    .B(net596),
    .X(_0176_));
 sg13g2_nand3_1 _5789_ (.B(net2157),
    .C(_1398_),
    .A(\draw_game_inst.y[8] ),
    .Y(_1405_));
 sg13g2_o21ai_1 _5790_ (.B1(net1040),
    .Y(_1406_),
    .A1(net2122),
    .A2(net2123));
 sg13g2_nand2_1 _5791_ (.Y(_1407_),
    .A(net2290),
    .B(_3992_));
 sg13g2_nand4_1 _5792_ (.B(_3992_),
    .C(_1405_),
    .A(net2290),
    .Y(_1408_),
    .D(_1406_));
 sg13g2_nor2b_2 _5793_ (.A(\draw_game_inst.board_y[6] ),
    .B_N(net2152),
    .Y(_1409_));
 sg13g2_nor2_1 _5794_ (.A(net2175),
    .B(net2193),
    .Y(_1410_));
 sg13g2_nand2_1 _5795_ (.Y(_1411_),
    .A(net2050),
    .B(net2043));
 sg13g2_nor2_1 _5796_ (.A(net2248),
    .B(net2221),
    .Y(_1412_));
 sg13g2_or2_1 _5797_ (.X(_1413_),
    .B(net2204),
    .A(net2231));
 sg13g2_nor3_1 _5798_ (.A(net2157),
    .B(net2162),
    .C(net1981),
    .Y(_1414_));
 sg13g2_and2_1 _5799_ (.A(net1992),
    .B(_1414_),
    .X(_1415_));
 sg13g2_or2_1 _5800_ (.X(_1416_),
    .B(\draw_game_inst.y[8] ),
    .A(net1042));
 sg13g2_nor2_1 _5801_ (.A(\draw_game_inst.y[8] ),
    .B(_0088_),
    .Y(_1417_));
 sg13g2_a221oi_1 _5802_ (.B2(_0088_),
    .C1(_1417_),
    .B1(_1416_),
    .A1(_1409_),
    .Y(_1418_),
    .A2(_1415_));
 sg13g2_and2_1 _5803_ (.A(net2123),
    .B(net2128),
    .X(_1419_));
 sg13g2_or2_1 _5804_ (.X(_1420_),
    .B(net1979),
    .A(net2122));
 sg13g2_a21oi_1 _5805_ (.A1(net2122),
    .A2(net1979),
    .Y(_1421_),
    .B1(net1040));
 sg13g2_nand3_1 _5806_ (.B(_1420_),
    .C(_1421_),
    .A(_3992_),
    .Y(_1422_));
 sg13g2_and3_1 _5807_ (.X(_1423_),
    .A(_1397_),
    .B(_1409_),
    .C(_1415_));
 sg13g2_nor3_2 _5808_ (.A(_1418_),
    .B(_1422_),
    .C(_1423_),
    .Y(_1424_));
 sg13g2_inv_1 _5809_ (.Y(_1425_),
    .A(_1424_));
 sg13g2_nor2_2 _5810_ (.A(net2123),
    .B(net2128),
    .Y(_1426_));
 sg13g2_nor2_2 _5811_ (.A(net1980),
    .B(net1978),
    .Y(_1427_));
 sg13g2_mux2_1 _5812_ (.A0(\draw_game_inst.grid[47] ),
    .A1(\draw_game_inst.grid[43] ),
    .S(net2127),
    .X(_1428_));
 sg13g2_a21oi_1 _5813_ (.A1(\draw_game_inst.grid[39] ),
    .A2(net1978),
    .Y(_1429_),
    .B1(net2154));
 sg13g2_a22oi_1 _5814_ (.Y(_1430_),
    .B1(_1427_),
    .B2(_1428_),
    .A2(net1980),
    .A1(\draw_game_inst.grid[35] ));
 sg13g2_mux2_1 _5815_ (.A0(\draw_game_inst.grid[63] ),
    .A1(\draw_game_inst.grid[59] ),
    .S(net2127),
    .X(_1431_));
 sg13g2_a21oi_1 _5816_ (.A1(\draw_game_inst.grid[55] ),
    .A2(net1978),
    .Y(_1432_),
    .B1(_3993_));
 sg13g2_a22oi_1 _5817_ (.Y(_1433_),
    .B1(_1427_),
    .B2(_1431_),
    .A2(net1980),
    .A1(\draw_game_inst.grid[51] ));
 sg13g2_a221oi_1 _5818_ (.B2(_1433_),
    .C1(net2153),
    .B1(_1432_),
    .A1(_1429_),
    .Y(_1434_),
    .A2(_1430_));
 sg13g2_mux4_1 _5819_ (.S0(net2126),
    .A0(\draw_game_inst.grid[7] ),
    .A1(\draw_game_inst.grid[11] ),
    .A2(\draw_game_inst.grid[15] ),
    .A3(\draw_game_inst.grid[3] ),
    .S1(net2124),
    .X(_1435_));
 sg13g2_mux4_1 _5820_ (.S0(net2126),
    .A0(\draw_game_inst.grid[23] ),
    .A1(\draw_game_inst.grid[27] ),
    .A2(\draw_game_inst.grid[31] ),
    .A3(\draw_game_inst.grid[19] ),
    .S1(net2124),
    .X(_1436_));
 sg13g2_a22oi_1 _5821_ (.Y(_1437_),
    .B1(_1436_),
    .B2(_1398_),
    .A2(_1435_),
    .A1(_1409_));
 sg13g2_nand2b_2 _5822_ (.Y(_1438_),
    .B(_1437_),
    .A_N(_1434_));
 sg13g2_mux2_1 _5823_ (.A0(\draw_game_inst.grid[61] ),
    .A1(\draw_game_inst.grid[57] ),
    .S(net2126),
    .X(_1439_));
 sg13g2_nand2_1 _5824_ (.Y(_1440_),
    .A(\draw_game_inst.grid[53] ),
    .B(net1978));
 sg13g2_a221oi_1 _5825_ (.B2(_1439_),
    .C1(_3993_),
    .B1(_1427_),
    .A1(\draw_game_inst.grid[49] ),
    .Y(_1441_),
    .A2(net1980));
 sg13g2_mux2_1 _5826_ (.A0(\draw_game_inst.grid[45] ),
    .A1(\draw_game_inst.grid[41] ),
    .S(net2127),
    .X(_1442_));
 sg13g2_a21oi_1 _5827_ (.A1(\draw_game_inst.grid[37] ),
    .A2(net1978),
    .Y(_1443_),
    .B1(net2154));
 sg13g2_a22oi_1 _5828_ (.Y(_1444_),
    .B1(_1427_),
    .B2(_1442_),
    .A2(net1980),
    .A1(\draw_game_inst.grid[33] ));
 sg13g2_a221oi_1 _5829_ (.B2(_1444_),
    .C1(net2153),
    .B1(_1443_),
    .A1(_1440_),
    .Y(_1445_),
    .A2(_1441_));
 sg13g2_mux4_1 _5830_ (.S0(net2126),
    .A0(\draw_game_inst.grid[5] ),
    .A1(\draw_game_inst.grid[9] ),
    .A2(\draw_game_inst.grid[13] ),
    .A3(\draw_game_inst.grid[1] ),
    .S1(net2124),
    .X(_1446_));
 sg13g2_mux4_1 _5831_ (.S0(net2126),
    .A0(\draw_game_inst.grid[21] ),
    .A1(\draw_game_inst.grid[25] ),
    .A2(\draw_game_inst.grid[29] ),
    .A3(\draw_game_inst.grid[17] ),
    .S1(net2124),
    .X(_1447_));
 sg13g2_a22oi_1 _5832_ (.Y(_1448_),
    .B1(_1447_),
    .B2(_1398_),
    .A2(_1446_),
    .A1(_1409_));
 sg13g2_nand2b_1 _5833_ (.Y(_1449_),
    .B(_1448_),
    .A_N(_1445_));
 sg13g2_inv_2 _5834_ (.Y(_1450_),
    .A(_1449_));
 sg13g2_mux2_1 _5835_ (.A0(\draw_game_inst.grid[62] ),
    .A1(\draw_game_inst.grid[58] ),
    .S(net2128),
    .X(_1451_));
 sg13g2_nand2_1 _5836_ (.Y(_1452_),
    .A(\draw_game_inst.grid[54] ),
    .B(net1978));
 sg13g2_a221oi_1 _5837_ (.B2(_1451_),
    .C1(_3993_),
    .B1(_1427_),
    .A1(\draw_game_inst.grid[50] ),
    .Y(_1453_),
    .A2(net1979));
 sg13g2_mux2_1 _5838_ (.A0(\draw_game_inst.grid[46] ),
    .A1(\draw_game_inst.grid[42] ),
    .S(net2128),
    .X(_1454_));
 sg13g2_a21oi_1 _5839_ (.A1(\draw_game_inst.grid[38] ),
    .A2(_1426_),
    .Y(_1455_),
    .B1(net2154));
 sg13g2_a22oi_1 _5840_ (.Y(_1456_),
    .B1(_1427_),
    .B2(_1454_),
    .A2(net1979),
    .A1(\draw_game_inst.grid[34] ));
 sg13g2_a221oi_1 _5841_ (.B2(_1456_),
    .C1(net2152),
    .B1(_1455_),
    .A1(_1452_),
    .Y(_1457_),
    .A2(_1453_));
 sg13g2_mux4_1 _5842_ (.S0(net2128),
    .A0(\draw_game_inst.grid[6] ),
    .A1(\draw_game_inst.grid[10] ),
    .A2(\draw_game_inst.grid[14] ),
    .A3(\draw_game_inst.grid[2] ),
    .S1(net2123),
    .X(_1458_));
 sg13g2_mux4_1 _5843_ (.S0(net2128),
    .A0(\draw_game_inst.grid[22] ),
    .A1(\draw_game_inst.grid[26] ),
    .A2(\draw_game_inst.grid[30] ),
    .A3(\draw_game_inst.grid[18] ),
    .S1(net2123),
    .X(_1459_));
 sg13g2_a22oi_1 _5844_ (.Y(_1460_),
    .B1(_1459_),
    .B2(_1398_),
    .A2(_1458_),
    .A1(_1409_));
 sg13g2_nand2b_2 _5845_ (.Y(_1461_),
    .B(_1460_),
    .A_N(_1457_));
 sg13g2_nor2b_2 _5846_ (.A(_1461_),
    .B_N(_1438_),
    .Y(_1462_));
 sg13g2_inv_1 _5847_ (.Y(_1463_),
    .A(_1462_));
 sg13g2_nand2b_2 _5848_ (.Y(_1464_),
    .B(_1461_),
    .A_N(_1438_));
 sg13g2_o21ai_1 _5849_ (.B1(_1464_),
    .Y(_1465_),
    .A1(_1438_),
    .A2(_1450_));
 sg13g2_nor2_1 _5850_ (.A(_1462_),
    .B(_1465_),
    .Y(_1466_));
 sg13g2_mux4_1 _5851_ (.S0(net2126),
    .A0(\draw_game_inst.grid[20] ),
    .A1(\draw_game_inst.grid[24] ),
    .A2(\draw_game_inst.grid[28] ),
    .A3(\draw_game_inst.grid[16] ),
    .S1(net2124),
    .X(_1467_));
 sg13g2_mux4_1 _5852_ (.S0(net2126),
    .A0(\draw_game_inst.grid[52] ),
    .A1(\draw_game_inst.grid[56] ),
    .A2(\draw_game_inst.grid[60] ),
    .A3(\draw_game_inst.grid[48] ),
    .S1(net2124),
    .X(_1468_));
 sg13g2_mux4_1 _5853_ (.S0(net2126),
    .A0(\draw_game_inst.grid[4] ),
    .A1(\draw_game_inst.grid[8] ),
    .A2(\draw_game_inst.grid[12] ),
    .A3(\draw_game_inst.grid[0] ),
    .S1(net2124),
    .X(_1469_));
 sg13g2_mux4_1 _5854_ (.S0(net2127),
    .A0(\draw_game_inst.grid[36] ),
    .A1(\draw_game_inst.grid[40] ),
    .A2(\draw_game_inst.grid[44] ),
    .A3(\draw_game_inst.grid[32] ),
    .S1(net2124),
    .X(_1470_));
 sg13g2_nand2_1 _5855_ (.Y(_1471_),
    .A(_3993_),
    .B(_1470_));
 sg13g2_nand2_1 _5856_ (.Y(_1472_),
    .A(net2154),
    .B(_1468_));
 sg13g2_a21oi_1 _5857_ (.A1(_1471_),
    .A2(_1472_),
    .Y(_1473_),
    .B1(net2153));
 sg13g2_a221oi_1 _5858_ (.B2(_1409_),
    .C1(_1473_),
    .B1(_1469_),
    .A1(_1398_),
    .Y(_1474_),
    .A2(_1467_));
 sg13g2_or2_1 _5859_ (.X(_1475_),
    .B(_1474_),
    .A(_1449_));
 sg13g2_nor2_2 _5860_ (.A(_1438_),
    .B(_1461_),
    .Y(_1476_));
 sg13g2_inv_1 _5861_ (.Y(_1477_),
    .A(_1476_));
 sg13g2_o21ai_1 _5862_ (.B1(net1731),
    .Y(_1478_),
    .A1(_1475_),
    .A2(_1477_));
 sg13g2_nor2_2 _5863_ (.A(_1464_),
    .B(_1475_),
    .Y(_1479_));
 sg13g2_nor2_2 _5864_ (.A(net2172),
    .B(net2205),
    .Y(_1480_));
 sg13g2_nand2_2 _5865_ (.Y(_1481_),
    .A(net2049),
    .B(net2035));
 sg13g2_nor2_1 _5866_ (.A(net2212),
    .B(net1889),
    .Y(_1482_));
 sg13g2_nand2_2 _5867_ (.Y(_1483_),
    .A(net2033),
    .B(net1993));
 sg13g2_nor2_2 _5868_ (.A(net2028),
    .B(net2144),
    .Y(_1484_));
 sg13g2_nand2_2 _5869_ (.Y(_1485_),
    .A(net2150),
    .B(net2021));
 sg13g2_nor2b_1 _5870_ (.A(net2150),
    .B_N(net2136),
    .Y(_1486_));
 sg13g2_nand2_1 _5871_ (.Y(_1487_),
    .A(net2028),
    .B(net2136));
 sg13g2_nor2_1 _5872_ (.A(net2149),
    .B(net2021),
    .Y(_1488_));
 sg13g2_nand2_1 _5873_ (.Y(_1489_),
    .A(_3999_),
    .B(net2141));
 sg13g2_nor2_2 _5874_ (.A(net2149),
    .B(net1996),
    .Y(_1490_));
 sg13g2_nand2_2 _5875_ (.Y(_1491_),
    .A(net2027),
    .B(_1400_));
 sg13g2_nor2_1 _5876_ (.A(net1886),
    .B(net1881),
    .Y(_1492_));
 sg13g2_nand2_1 _5877_ (.Y(_1493_),
    .A(_1485_),
    .B(net1879));
 sg13g2_nor2_1 _5878_ (.A(net2027),
    .B(net2022),
    .Y(_1494_));
 sg13g2_nand2_1 _5879_ (.Y(_1495_),
    .A(net2147),
    .B(net2144));
 sg13g2_nor2_2 _5880_ (.A(net2204),
    .B(net1876),
    .Y(_1496_));
 sg13g2_nor2_2 _5881_ (.A(net2147),
    .B(net2135),
    .Y(_1497_));
 sg13g2_nor2_1 _5882_ (.A(net2149),
    .B(net2141),
    .Y(_1498_));
 sg13g2_nand2_2 _5883_ (.Y(_1499_),
    .A(_3999_),
    .B(net2021));
 sg13g2_nand2_2 _5884_ (.Y(_1500_),
    .A(net2023),
    .B(net1973));
 sg13g2_o21ai_1 _5885_ (.B1(net1813),
    .Y(_1501_),
    .A1(net1976),
    .A2(net1807));
 sg13g2_nand3_1 _5886_ (.B(net2163),
    .C(_1501_),
    .A(net2158),
    .Y(_1502_));
 sg13g2_nand2_1 _5887_ (.Y(_1503_),
    .A(net1743),
    .B(_1502_));
 sg13g2_and2_1 _5888_ (.A(net2246),
    .B(net2220),
    .X(_1504_));
 sg13g2_nand2_2 _5889_ (.Y(_1505_),
    .A(net2246),
    .B(net2220));
 sg13g2_nor2_2 _5890_ (.A(net2139),
    .B(net2023),
    .Y(_1506_));
 sg13g2_nand2b_2 _5891_ (.Y(_1507_),
    .B(net2144),
    .A_N(net2135));
 sg13g2_nor2_1 _5892_ (.A(net2148),
    .B(net1958),
    .Y(_1508_));
 sg13g2_nand2_2 _5893_ (.Y(_1509_),
    .A(net2028),
    .B(_1506_));
 sg13g2_nor2_1 _5894_ (.A(net2132),
    .B(net1878),
    .Y(_1510_));
 sg13g2_nand2b_1 _5895_ (.Y(_1511_),
    .B(net1881),
    .A_N(net2132));
 sg13g2_nor2_2 _5896_ (.A(net1875),
    .B(net1806),
    .Y(_1512_));
 sg13g2_nand2_2 _5897_ (.Y(_1513_),
    .A(_1509_),
    .B(net1805));
 sg13g2_nand2_2 _5898_ (.Y(_1514_),
    .A(net2219),
    .B(net1878));
 sg13g2_nand2_2 _5899_ (.Y(_1515_),
    .A(net2214),
    .B(net2138));
 sg13g2_nand2_2 _5900_ (.Y(_1516_),
    .A(net2217),
    .B(_1509_));
 sg13g2_nor2_2 _5901_ (.A(net2032),
    .B(net1806),
    .Y(_1517_));
 sg13g2_o21ai_1 _5902_ (.B1(net1964),
    .Y(_1518_),
    .A1(net2033),
    .A2(_1513_));
 sg13g2_nand2b_2 _5903_ (.Y(_1519_),
    .B(net1879),
    .A_N(net2244));
 sg13g2_nor2b_1 _5904_ (.A(net2205),
    .B_N(net2231),
    .Y(_1520_));
 sg13g2_nand2_2 _5905_ (.Y(_1521_),
    .A(net2236),
    .B(net2031));
 sg13g2_nor2b_2 _5906_ (.A(net1875),
    .B_N(net2248),
    .Y(_1522_));
 sg13g2_nor2_1 _5907_ (.A(net1875),
    .B(_1521_),
    .Y(_1523_));
 sg13g2_a21oi_2 _5908_ (.B1(_1523_),
    .Y(_1524_),
    .A2(net1879),
    .A1(net1988));
 sg13g2_nor2_2 _5909_ (.A(_1510_),
    .B(_1524_),
    .Y(_1525_));
 sg13g2_nor3_1 _5910_ (.A(net2193),
    .B(_1518_),
    .C(_1525_),
    .Y(_1526_));
 sg13g2_nand2_2 _5911_ (.Y(_1527_),
    .A(net2193),
    .B(net1983));
 sg13g2_inv_1 _5912_ (.Y(_1528_),
    .A(_1527_));
 sg13g2_nor2b_1 _5913_ (.A(net2136),
    .B_N(net2149),
    .Y(_1529_));
 sg13g2_nand2_2 _5914_ (.Y(_1530_),
    .A(net2150),
    .B(net2024));
 sg13g2_nor2_1 _5915_ (.A(net2134),
    .B(net1974),
    .Y(_1531_));
 sg13g2_nand2_1 _5916_ (.Y(_1532_),
    .A(net2140),
    .B(net1952));
 sg13g2_nor2_2 _5917_ (.A(net2211),
    .B(net1870),
    .Y(_1533_));
 sg13g2_nor2_2 _5918_ (.A(net2024),
    .B(net2140),
    .Y(_1534_));
 sg13g2_nand2b_1 _5919_ (.Y(_1535_),
    .B(net2135),
    .A_N(net2144));
 sg13g2_nor2_2 _5920_ (.A(_1506_),
    .B(net1868),
    .Y(_1536_));
 sg13g2_nand2_2 _5921_ (.Y(_1537_),
    .A(net1958),
    .B(net1951));
 sg13g2_nor2_2 _5922_ (.A(net2027),
    .B(_1536_),
    .Y(_1538_));
 sg13g2_nand2_1 _5923_ (.Y(_1539_),
    .A(net2151),
    .B(_1537_));
 sg13g2_nand2_1 _5924_ (.Y(_1540_),
    .A(net2211),
    .B(_1538_));
 sg13g2_a21oi_1 _5925_ (.A1(net2211),
    .A2(_1538_),
    .Y(_1541_),
    .B1(_1533_));
 sg13g2_o21ai_1 _5926_ (.B1(net2048),
    .Y(_1542_),
    .A1(_1527_),
    .A2(_1541_));
 sg13g2_nor2_1 _5927_ (.A(net1959),
    .B(net1869),
    .Y(_1543_));
 sg13g2_nand2_2 _5928_ (.Y(_1544_),
    .A(net1965),
    .B(net1871));
 sg13g2_nor2_1 _5929_ (.A(net1902),
    .B(net1960),
    .Y(_1545_));
 sg13g2_nand2_2 _5930_ (.Y(_1546_),
    .A(net1910),
    .B(net1968));
 sg13g2_nand2_1 _5931_ (.Y(_1547_),
    .A(net1911),
    .B(net1803));
 sg13g2_nand2_1 _5932_ (.Y(_1548_),
    .A(_1546_),
    .B(_1547_));
 sg13g2_nor2_2 _5933_ (.A(net1976),
    .B(net1952),
    .Y(_1549_));
 sg13g2_nand2_2 _5934_ (.Y(_1550_),
    .A(net1883),
    .B(_1530_));
 sg13g2_nor2_2 _5935_ (.A(net2147),
    .B(net1950),
    .Y(_1551_));
 sg13g2_nand2_1 _5936_ (.Y(_1552_),
    .A(net2021),
    .B(net1976));
 sg13g2_nor2_2 _5937_ (.A(net2140),
    .B(_1530_),
    .Y(_1553_));
 sg13g2_nand2_2 _5938_ (.Y(_1554_),
    .A(net2021),
    .B(net1952));
 sg13g2_nor2_2 _5939_ (.A(net2141),
    .B(_1549_),
    .Y(_1555_));
 sg13g2_nand2_2 _5940_ (.Y(_1556_),
    .A(net2022),
    .B(_1550_));
 sg13g2_nand2_1 _5941_ (.Y(_1557_),
    .A(net2230),
    .B(net1950));
 sg13g2_nor2b_2 _5942_ (.A(net1977),
    .B_N(net2242),
    .Y(_1558_));
 sg13g2_nand2_2 _5943_ (.Y(_1559_),
    .A(net2242),
    .B(net1883));
 sg13g2_nor2_1 _5944_ (.A(net1807),
    .B(_1559_),
    .Y(_1560_));
 sg13g2_nor2_1 _5945_ (.A(net2034),
    .B(_1560_),
    .Y(_1561_));
 sg13g2_o21ai_1 _5946_ (.B1(_1561_),
    .Y(_1562_),
    .A1(net2238),
    .A2(_1555_));
 sg13g2_nand2_2 _5947_ (.Y(_1563_),
    .A(net2187),
    .B(net1869));
 sg13g2_o21ai_1 _5948_ (.B1(net2191),
    .Y(_1564_),
    .A1(net1983),
    .A2(net1870));
 sg13g2_nor2_2 _5949_ (.A(net2048),
    .B(_1564_),
    .Y(_1565_));
 sg13g2_a221oi_1 _5950_ (.B2(_1565_),
    .C1(net2052),
    .B1(_1562_),
    .A1(_1544_),
    .Y(_1566_),
    .A2(_1548_));
 sg13g2_o21ai_1 _5951_ (.B1(_1566_),
    .Y(_1567_),
    .A1(_1526_),
    .A2(_1542_));
 sg13g2_nand2_1 _5952_ (.Y(_1568_),
    .A(net2155),
    .B(net2162));
 sg13g2_nand2_2 _5953_ (.Y(_1569_),
    .A(net2149),
    .B(net2137));
 sg13g2_nor2_2 _5954_ (.A(net2140),
    .B(net1947),
    .Y(_1570_));
 sg13g2_nand2_2 _5955_ (.Y(_1571_),
    .A(net2139),
    .B(net1885));
 sg13g2_nand2_2 _5956_ (.Y(_1572_),
    .A(_1537_),
    .B(net1867));
 sg13g2_nor2b_2 _5957_ (.A(net2212),
    .B_N(net2226),
    .Y(_1573_));
 sg13g2_nand2_2 _5958_ (.Y(_1574_),
    .A(net2226),
    .B(net2034));
 sg13g2_o21ai_1 _5959_ (.B1(net2034),
    .Y(_1575_),
    .A1(net2226),
    .A2(_1572_));
 sg13g2_nor2_1 _5960_ (.A(net2036),
    .B(net1886),
    .Y(_1576_));
 sg13g2_nand2_2 _5961_ (.Y(_1577_),
    .A(net2210),
    .B(net1810));
 sg13g2_a21o_1 _5962_ (.A2(_1577_),
    .A1(_1575_),
    .B1(net1889),
    .X(_1578_));
 sg13g2_nor2_1 _5963_ (.A(net2218),
    .B(net1806),
    .Y(_1579_));
 sg13g2_nor2_2 _5964_ (.A(net1945),
    .B(_1579_),
    .Y(_1580_));
 sg13g2_nand2b_2 _5965_ (.Y(_1581_),
    .B(net1804),
    .A_N(net2240));
 sg13g2_nand4_1 _5966_ (.B(_1513_),
    .C(_1580_),
    .A(net2191),
    .Y(_1582_),
    .D(_1581_));
 sg13g2_nor2_2 _5967_ (.A(net2225),
    .B(net2032),
    .Y(_1583_));
 sg13g2_nand2b_1 _5968_ (.Y(_1584_),
    .B(net2200),
    .A_N(net2225));
 sg13g2_nor2_1 _5969_ (.A(net2186),
    .B(_1583_),
    .Y(_1585_));
 sg13g2_nand2_2 _5970_ (.Y(_1586_),
    .A(net1865),
    .B(_1585_));
 sg13g2_nand3_1 _5971_ (.B(_1582_),
    .C(_1586_),
    .A(net2178),
    .Y(_1587_));
 sg13g2_nor2_1 _5972_ (.A(net2155),
    .B(net2161),
    .Y(_1588_));
 sg13g2_or2_1 _5973_ (.X(_1589_),
    .B(net2161),
    .A(net2156));
 sg13g2_nor2_1 _5974_ (.A(net2175),
    .B(net2043),
    .Y(_1590_));
 sg13g2_nand2_1 _5975_ (.Y(_1591_),
    .A(net2050),
    .B(net2193));
 sg13g2_nand2_2 _5976_ (.Y(_1592_),
    .A(net2142),
    .B(net1977));
 sg13g2_nand2_2 _5977_ (.Y(_1593_),
    .A(net2026),
    .B(_1485_));
 sg13g2_nor2_2 _5978_ (.A(net2138),
    .B(net1886),
    .Y(_1594_));
 sg13g2_nand2_2 _5979_ (.Y(_1595_),
    .A(_1536_),
    .B(_1550_));
 sg13g2_nor2_2 _5980_ (.A(_1537_),
    .B(net1867),
    .Y(_1596_));
 sg13g2_o21ai_1 _5981_ (.B1(net1859),
    .Y(_1597_),
    .A1(_1583_),
    .A2(_1595_));
 sg13g2_nand4_1 _5982_ (.B(_1587_),
    .C(net1944),
    .A(_1578_),
    .Y(_1598_),
    .D(_1597_));
 sg13g2_and2_1 _5983_ (.A(net1948),
    .B(_1598_),
    .X(_1599_));
 sg13g2_a21oi_2 _5984_ (.B1(_1503_),
    .Y(_1600_),
    .A2(_1599_),
    .A1(_1567_));
 sg13g2_nand2_2 _5985_ (.Y(_1601_),
    .A(_1450_),
    .B(_1474_));
 sg13g2_nor2_2 _5986_ (.A(_1464_),
    .B(_1601_),
    .Y(_1602_));
 sg13g2_nand2_1 _5987_ (.Y(_1603_),
    .A(net1892),
    .B(net1808));
 sg13g2_a21oi_1 _5988_ (.A1(_1400_),
    .A2(net1807),
    .Y(_1604_),
    .B1(net2239));
 sg13g2_a21oi_1 _5989_ (.A1(net2239),
    .A2(_1572_),
    .Y(_1605_),
    .B1(net1887));
 sg13g2_nor2b_1 _5990_ (.A(_1604_),
    .B_N(_1605_),
    .Y(_1606_));
 sg13g2_o21ai_1 _5991_ (.B1(net1730),
    .Y(_1607_),
    .A1(net1949),
    .A2(_1606_));
 sg13g2_nor2_2 _5992_ (.A(net2048),
    .B(net2043),
    .Y(_1608_));
 sg13g2_nand2_1 _5993_ (.Y(_1609_),
    .A(net2180),
    .B(net2196));
 sg13g2_nor2b_2 _5994_ (.A(net1953),
    .B_N(net2247),
    .Y(_1610_));
 sg13g2_nand2_1 _5995_ (.Y(_1611_),
    .A(net1807),
    .B(_1610_));
 sg13g2_nand3_1 _5996_ (.B(net1853),
    .C(_1611_),
    .A(_1518_),
    .Y(_1612_));
 sg13g2_nor2_2 _5997_ (.A(net2151),
    .B(_1536_),
    .Y(_1613_));
 sg13g2_nand2_1 _5998_ (.Y(_1614_),
    .A(net2027),
    .B(_1537_));
 sg13g2_nor2_2 _5999_ (.A(net2207),
    .B(_1402_),
    .Y(_1615_));
 sg13g2_nor2_2 _6000_ (.A(net2043),
    .B(net2033),
    .Y(_1616_));
 sg13g2_nand2_1 _6001_ (.Y(_1617_),
    .A(net2193),
    .B(net2212));
 sg13g2_nor3_1 _6002_ (.A(_1490_),
    .B(net1859),
    .C(_1616_),
    .Y(_1618_));
 sg13g2_a221oi_1 _6003_ (.B2(net1909),
    .C1(_1618_),
    .B1(_1615_),
    .A1(net1859),
    .Y(_1619_),
    .A2(net1799));
 sg13g2_a21oi_1 _6004_ (.A1(_1612_),
    .A2(_1619_),
    .Y(_1620_),
    .B1(net1895));
 sg13g2_nand2_2 _6005_ (.Y(_1621_),
    .A(net2219),
    .B(_1603_));
 sg13g2_a21oi_1 _6006_ (.A1(_1575_),
    .A2(_1621_),
    .Y(_1622_),
    .B1(net1889));
 sg13g2_nor2_2 _6007_ (.A(net2177),
    .B(net1930),
    .Y(_1623_));
 sg13g2_nor2_2 _6008_ (.A(net2136),
    .B(net1810),
    .Y(_1624_));
 sg13g2_nand2_2 _6009_ (.Y(_1625_),
    .A(net2024),
    .B(net1807));
 sg13g2_nand2_1 _6010_ (.Y(_1626_),
    .A(_1558_),
    .B(net1790));
 sg13g2_o21ai_1 _6011_ (.B1(_1626_),
    .Y(_1627_),
    .A1(_1519_),
    .A2(net1801));
 sg13g2_nand2_1 _6012_ (.Y(_1628_),
    .A(_1623_),
    .B(_1627_));
 sg13g2_nor2_2 _6013_ (.A(net2034),
    .B(net1934),
    .Y(_1629_));
 sg13g2_nand2_2 _6014_ (.Y(_1630_),
    .A(net2212),
    .B(net1853));
 sg13g2_nor2_2 _6015_ (.A(net1959),
    .B(net1933),
    .Y(_1631_));
 sg13g2_nand2_2 _6016_ (.Y(_1632_),
    .A(net1965),
    .B(net1851));
 sg13g2_nor2b_1 _6017_ (.A(net2142),
    .B_N(net2132),
    .Y(_1633_));
 sg13g2_nor2_1 _6018_ (.A(net1876),
    .B(_1633_),
    .Y(_1634_));
 sg13g2_inv_1 _6019_ (.Y(_1635_),
    .A(_1634_));
 sg13g2_nor2_2 _6020_ (.A(net2246),
    .B(net2036),
    .Y(_1636_));
 sg13g2_a22oi_1 _6021_ (.Y(_1637_),
    .B1(_1635_),
    .B2(net1849),
    .A2(net1967),
    .A1(_1491_));
 sg13g2_nor2_1 _6022_ (.A(net1934),
    .B(_1637_),
    .Y(_1638_));
 sg13g2_nand3_1 _6023_ (.B(net2023),
    .C(net1953),
    .A(net2239),
    .Y(_1639_));
 sg13g2_nor2_1 _6024_ (.A(net2043),
    .B(net2212),
    .Y(_1640_));
 sg13g2_nand2_2 _6025_ (.Y(_1641_),
    .A(net2193),
    .B(net2033));
 sg13g2_nor2_1 _6026_ (.A(net2175),
    .B(_1641_),
    .Y(_1642_));
 sg13g2_nand2_1 _6027_ (.Y(_1643_),
    .A(net2048),
    .B(net1845));
 sg13g2_nand2_1 _6028_ (.Y(_1644_),
    .A(net2236),
    .B(net1971));
 sg13g2_nand2_2 _6029_ (.Y(_1645_),
    .A(net2036),
    .B(net1879));
 sg13g2_nand3_1 _6030_ (.B(_1639_),
    .C(net1798),
    .A(net1878),
    .Y(_1646_));
 sg13g2_nor2_2 _6031_ (.A(net2212),
    .B(net1934),
    .Y(_1647_));
 sg13g2_nand2_1 _6032_ (.Y(_1648_),
    .A(net2037),
    .B(net1855));
 sg13g2_nor2_1 _6033_ (.A(net2230),
    .B(net1868),
    .Y(_1649_));
 sg13g2_nand2b_1 _6034_ (.Y(_1650_),
    .B(net1951),
    .A_N(net2240));
 sg13g2_nor2_2 _6035_ (.A(net2246),
    .B(net2027),
    .Y(_1651_));
 sg13g2_nand2b_2 _6036_ (.Y(_1652_),
    .B(net2147),
    .A_N(net2232));
 sg13g2_nor2_2 _6037_ (.A(net2234),
    .B(_1506_),
    .Y(_1653_));
 sg13g2_nor2_2 _6038_ (.A(net2244),
    .B(net1875),
    .Y(_1654_));
 sg13g2_nand2_1 _6039_ (.Y(_1655_),
    .A(net1950),
    .B(_1654_));
 sg13g2_nor2b_2 _6040_ (.A(_1634_),
    .B_N(net2243),
    .Y(_1656_));
 sg13g2_a21oi_1 _6041_ (.A1(net1951),
    .A2(_1654_),
    .Y(_1657_),
    .B1(_1656_));
 sg13g2_o21ai_1 _6042_ (.B1(_1646_),
    .Y(_1658_),
    .A1(_1648_),
    .A2(_1657_));
 sg13g2_or3_1 _6043_ (.A(net2161),
    .B(_1638_),
    .C(_1658_),
    .X(_1659_));
 sg13g2_nand2_2 _6044_ (.Y(_1660_),
    .A(net2238),
    .B(net1799));
 sg13g2_o21ai_1 _6045_ (.B1(_1660_),
    .Y(_1661_),
    .A1(net2238),
    .A2(_1555_));
 sg13g2_nor2_2 _6046_ (.A(net2210),
    .B(_1661_),
    .Y(_1662_));
 sg13g2_nor3_1 _6047_ (.A(net1906),
    .B(_1613_),
    .C(_1662_),
    .Y(_1663_));
 sg13g2_nor3_1 _6048_ (.A(_1622_),
    .B(_1659_),
    .C(_1663_),
    .Y(_1664_));
 sg13g2_a21oi_1 _6049_ (.A1(_1628_),
    .A2(_1664_),
    .Y(_1665_),
    .B1(net2159));
 sg13g2_nor3_1 _6050_ (.A(_1607_),
    .B(_1620_),
    .C(_1665_),
    .Y(_1666_));
 sg13g2_and2_2 _6051_ (.A(_1449_),
    .B(_1474_),
    .X(_1667_));
 sg13g2_and2_2 _6052_ (.A(_1476_),
    .B(_1667_),
    .X(_1668_));
 sg13g2_nor2_2 _6053_ (.A(net2196),
    .B(net2220),
    .Y(_1669_));
 sg13g2_nand2_2 _6054_ (.Y(_1670_),
    .A(net2038),
    .B(net2032));
 sg13g2_a21oi_1 _6055_ (.A1(net1813),
    .A2(net1865),
    .Y(_1671_),
    .B1(net1949));
 sg13g2_nor2b_2 _6056_ (.A(_1671_),
    .B_N(_1668_),
    .Y(_1672_));
 sg13g2_nor2_2 _6057_ (.A(net1871),
    .B(net1865),
    .Y(_1673_));
 sg13g2_nand2_2 _6058_ (.Y(_1674_),
    .A(net1869),
    .B(net1861));
 sg13g2_nand2_2 _6059_ (.Y(_1675_),
    .A(net2045),
    .B(net1861));
 sg13g2_a21oi_1 _6060_ (.A1(net1991),
    .A2(net1945),
    .Y(_1676_),
    .B1(net2161));
 sg13g2_nand3_1 _6061_ (.B(_1675_),
    .C(_1676_),
    .A(_1674_),
    .Y(_1677_));
 sg13g2_nand2_2 _6062_ (.Y(_1678_),
    .A(net2166),
    .B(net1861));
 sg13g2_nor2_1 _6063_ (.A(net2186),
    .B(_1678_),
    .Y(_1679_));
 sg13g2_o21ai_1 _6064_ (.B1(net2051),
    .Y(_1680_),
    .A1(_1677_),
    .A2(_1679_));
 sg13g2_nor3_1 _6065_ (.A(net2190),
    .B(_1533_),
    .C(net1865),
    .Y(_1681_));
 sg13g2_nor2_1 _6066_ (.A(net2168),
    .B(_1681_),
    .Y(_1682_));
 sg13g2_nor2_2 _6067_ (.A(net2203),
    .B(net2148),
    .Y(_1683_));
 sg13g2_nand2_2 _6068_ (.Y(_1684_),
    .A(net2032),
    .B(net1971));
 sg13g2_nand2_2 _6069_ (.Y(_1685_),
    .A(net1868),
    .B(_1683_));
 sg13g2_nand2_1 _6070_ (.Y(_1686_),
    .A(net2186),
    .B(_1685_));
 sg13g2_nor2_2 _6071_ (.A(net2236),
    .B(net1971),
    .Y(_1687_));
 sg13g2_o21ai_1 _6072_ (.B1(net2199),
    .Y(_1688_),
    .A1(net2229),
    .A2(net1971));
 sg13g2_nor2_1 _6073_ (.A(_1536_),
    .B(_1688_),
    .Y(_1689_));
 sg13g2_o21ai_1 _6074_ (.B1(_1682_),
    .Y(_1690_),
    .A1(_1686_),
    .A2(_1689_));
 sg13g2_nand2_1 _6075_ (.Y(_1691_),
    .A(net2038),
    .B(_1536_));
 sg13g2_nand2_1 _6076_ (.Y(_1692_),
    .A(net2187),
    .B(net1863));
 sg13g2_nand2_2 _6077_ (.Y(_1693_),
    .A(net2211),
    .B(net1882));
 sg13g2_nand4_1 _6078_ (.B(_1691_),
    .C(_1692_),
    .A(net2170),
    .Y(_1694_),
    .D(_1693_));
 sg13g2_nand3_1 _6079_ (.B(_1690_),
    .C(_1694_),
    .A(net1898),
    .Y(_1695_));
 sg13g2_nand3_1 _6080_ (.B(_1680_),
    .C(_1695_),
    .A(_1672_),
    .Y(_1696_));
 sg13g2_nor2_2 _6081_ (.A(_1450_),
    .B(_1474_),
    .Y(_1697_));
 sg13g2_nor3_2 _6082_ (.A(_1450_),
    .B(_1464_),
    .C(_1474_),
    .Y(_1698_));
 sg13g2_nand2_2 _6083_ (.Y(_1699_),
    .A(net2238),
    .B(net1864));
 sg13g2_nand2_2 _6084_ (.Y(_1700_),
    .A(net2139),
    .B(net1975));
 sg13g2_nor2_2 _6085_ (.A(net2026),
    .B(net1876),
    .Y(_1701_));
 sg13g2_nand2_2 _6086_ (.Y(_1702_),
    .A(net2134),
    .B(net1809));
 sg13g2_nand2_1 _6087_ (.Y(_1703_),
    .A(_1593_),
    .B(_1702_));
 sg13g2_a21oi_1 _6088_ (.A1(_1593_),
    .A2(_1702_),
    .Y(_1704_),
    .B1(net2235));
 sg13g2_a21oi_1 _6089_ (.A1(net2235),
    .A2(_1556_),
    .Y(_1705_),
    .B1(_1704_));
 sg13g2_a21oi_1 _6090_ (.A1(net2235),
    .A2(net1977),
    .Y(_1706_),
    .B1(net2031));
 sg13g2_nand2_1 _6091_ (.Y(_1707_),
    .A(_1556_),
    .B(_1706_));
 sg13g2_o21ai_1 _6092_ (.B1(_1707_),
    .Y(_1708_),
    .A1(net2208),
    .A2(_1705_));
 sg13g2_nor2_2 _6093_ (.A(net2231),
    .B(net1996),
    .Y(_1709_));
 sg13g2_nor3_2 _6094_ (.A(net2231),
    .B(net2029),
    .C(net1996),
    .Y(_1710_));
 sg13g2_a21oi_1 _6095_ (.A1(_1550_),
    .A2(_1710_),
    .Y(_1711_),
    .B1(_1703_));
 sg13g2_o21ai_1 _6096_ (.B1(net1943),
    .Y(_1712_),
    .A1(net1903),
    .A2(_1711_));
 sg13g2_nor2_2 _6097_ (.A(net2036),
    .B(net1954),
    .Y(_1713_));
 sg13g2_o21ai_1 _6098_ (.B1(_1550_),
    .Y(_1714_),
    .A1(net2022),
    .A2(_1651_));
 sg13g2_nor2_2 _6099_ (.A(net2219),
    .B(net1952),
    .Y(_1715_));
 sg13g2_nand2_2 _6100_ (.Y(_1716_),
    .A(net2030),
    .B(net1883));
 sg13g2_nand2_2 _6101_ (.Y(_1717_),
    .A(net1882),
    .B(_1715_));
 sg13g2_a21oi_2 _6102_ (.B1(net2184),
    .Y(_1718_),
    .A2(_1714_),
    .A1(net2216));
 sg13g2_nand2_1 _6103_ (.Y(_1719_),
    .A(_1717_),
    .B(_1718_));
 sg13g2_a221oi_1 _6104_ (.B2(net2047),
    .C1(_1712_),
    .B1(_1719_),
    .A1(net1855),
    .Y(_1720_),
    .A2(_1708_));
 sg13g2_nor2_2 _6105_ (.A(net2248),
    .B(net1977),
    .Y(_1721_));
 sg13g2_or2_2 _6106_ (.X(_1722_),
    .B(net1977),
    .A(net2241));
 sg13g2_a21oi_2 _6107_ (.B1(net1882),
    .Y(_1723_),
    .A2(net2143),
    .A1(net2227));
 sg13g2_nor2_2 _6108_ (.A(net2203),
    .B(net1996),
    .Y(_1724_));
 sg13g2_nor2_2 _6109_ (.A(net2221),
    .B(_1553_),
    .Y(_1725_));
 sg13g2_nor3_1 _6110_ (.A(_1483_),
    .B(net1801),
    .C(_1723_),
    .Y(_1726_));
 sg13g2_and2_1 _6111_ (.A(net2134),
    .B(net2145),
    .X(_1727_));
 sg13g2_nand2_1 _6112_ (.Y(_1728_),
    .A(net2138),
    .B(net2145));
 sg13g2_nor2_1 _6113_ (.A(_1594_),
    .B(_1727_),
    .Y(_1729_));
 sg13g2_nand2_2 _6114_ (.Y(_1730_),
    .A(_1593_),
    .B(_1728_));
 sg13g2_nor2_2 _6115_ (.A(net2248),
    .B(_1554_),
    .Y(_1731_));
 sg13g2_nor2_2 _6116_ (.A(net2035),
    .B(net1890),
    .Y(_1732_));
 sg13g2_nand2_2 _6117_ (.Y(_1733_),
    .A(net2216),
    .B(net1995));
 sg13g2_a221oi_1 _6118_ (.B2(net2234),
    .C1(_1733_),
    .B1(_1729_),
    .A1(net1996),
    .Y(_1734_),
    .A2(_1651_));
 sg13g2_o21ai_1 _6119_ (.B1(net1855),
    .Y(_1735_),
    .A1(net1983),
    .A2(net1867));
 sg13g2_nand2_2 _6120_ (.Y(_1736_),
    .A(net1901),
    .B(_1735_));
 sg13g2_nor2b_2 _6121_ (.A(net2137),
    .B_N(net2146),
    .Y(_1737_));
 sg13g2_nand2_1 _6122_ (.Y(_1738_),
    .A(net2024),
    .B(net2146));
 sg13g2_nand2_1 _6123_ (.Y(_1739_),
    .A(_1700_),
    .B(net1842));
 sg13g2_a22oi_1 _6124_ (.Y(_1740_),
    .B1(net1955),
    .B2(net1797),
    .A2(net1986),
    .A1(net2145));
 sg13g2_a22oi_1 _6125_ (.Y(_1741_),
    .B1(net1798),
    .B2(_1730_),
    .A2(_1623_),
    .A1(net2145));
 sg13g2_o21ai_1 _6126_ (.B1(net2208),
    .Y(_1742_),
    .A1(_1549_),
    .A2(_1709_));
 sg13g2_a21oi_1 _6127_ (.A1(_1740_),
    .A2(_1742_),
    .Y(_1743_),
    .B1(net1903));
 sg13g2_nand2b_1 _6128_ (.Y(_1744_),
    .B(_1741_),
    .A_N(_1736_));
 sg13g2_nor4_1 _6129_ (.A(_1726_),
    .B(_1734_),
    .C(_1743_),
    .D(_1744_),
    .Y(_1745_));
 sg13g2_o21ai_1 _6130_ (.B1(_1698_),
    .Y(_1746_),
    .A1(_1720_),
    .A2(_1745_));
 sg13g2_nor2_2 _6131_ (.A(_1463_),
    .B(_1475_),
    .Y(_1747_));
 sg13g2_and2_2 _6132_ (.A(net2132),
    .B(net1972),
    .X(_1748_));
 sg13g2_nand2_2 _6133_ (.Y(_1749_),
    .A(net2131),
    .B(net1971));
 sg13g2_nor2_1 _6134_ (.A(net2034),
    .B(_1748_),
    .Y(_1750_));
 sg13g2_a21o_1 _6135_ (.A2(net1841),
    .A1(net1966),
    .B1(_1710_),
    .X(_1751_));
 sg13g2_o21ai_1 _6136_ (.B1(net1852),
    .Y(_1752_),
    .A1(_1724_),
    .A2(_1751_));
 sg13g2_nor2_2 _6137_ (.A(net2027),
    .B(_1537_),
    .Y(_1753_));
 sg13g2_nand2_2 _6138_ (.Y(_1754_),
    .A(net2148),
    .B(_1536_));
 sg13g2_nor3_1 _6139_ (.A(net2230),
    .B(_1710_),
    .C(_1754_),
    .Y(_1755_));
 sg13g2_nor2_1 _6140_ (.A(_1752_),
    .B(_1755_),
    .Y(_1756_));
 sg13g2_nand2_1 _6141_ (.Y(_1757_),
    .A(net2171),
    .B(net1943));
 sg13g2_nor2_2 _6142_ (.A(net2184),
    .B(net1940),
    .Y(_1758_));
 sg13g2_nand2b_2 _6143_ (.Y(_1759_),
    .B(net1943),
    .A_N(net2184));
 sg13g2_a21oi_1 _6144_ (.A1(_1592_),
    .A2(_1724_),
    .Y(_1760_),
    .B1(_1759_));
 sg13g2_nor2_1 _6145_ (.A(net2233),
    .B(net1841),
    .Y(_1761_));
 sg13g2_nor2_1 _6146_ (.A(net1967),
    .B(_1750_),
    .Y(_1762_));
 sg13g2_and2_2 _6147_ (.A(net2246),
    .B(_1485_),
    .X(_1763_));
 sg13g2_nand2_2 _6148_ (.Y(_1764_),
    .A(net2244),
    .B(net1878));
 sg13g2_nand2b_1 _6149_ (.Y(_1765_),
    .B(_1594_),
    .A_N(_1764_));
 sg13g2_nand2b_2 _6150_ (.Y(_1766_),
    .B(_1765_),
    .A_N(_1762_));
 sg13g2_a22oi_1 _6151_ (.Y(_1767_),
    .B1(_1760_),
    .B2(_1766_),
    .A2(net1943),
    .A1(net2171));
 sg13g2_nand2b_1 _6152_ (.Y(_1768_),
    .B(net2149),
    .A_N(net2133));
 sg13g2_nor2_2 _6153_ (.A(net2131),
    .B(net1974),
    .Y(_1769_));
 sg13g2_or2_1 _6154_ (.X(_1770_),
    .B(net1975),
    .A(net2131));
 sg13g2_nor2_1 _6155_ (.A(net2031),
    .B(_1769_),
    .Y(_1771_));
 sg13g2_a22oi_1 _6156_ (.Y(_1772_),
    .B1(net1796),
    .B2(net1838),
    .A2(_1500_),
    .A1(_1496_));
 sg13g2_nor2_1 _6157_ (.A(net1902),
    .B(_1772_),
    .Y(_1773_));
 sg13g2_nor3_2 _6158_ (.A(_1756_),
    .B(_1767_),
    .C(_1773_),
    .Y(_1774_));
 sg13g2_nor2_1 _6159_ (.A(net2215),
    .B(_1748_),
    .Y(_1775_));
 sg13g2_nor2_1 _6160_ (.A(net2195),
    .B(_1775_),
    .Y(_1776_));
 sg13g2_or2_1 _6161_ (.X(_1777_),
    .B(net2146),
    .A(net2141));
 sg13g2_o21ai_1 _6162_ (.B1(_1777_),
    .Y(_1778_),
    .A1(net2021),
    .A2(net2132));
 sg13g2_and2_1 _6163_ (.A(net2248),
    .B(_1778_),
    .X(_1779_));
 sg13g2_o21ai_1 _6164_ (.B1(_1776_),
    .Y(_1780_),
    .A1(_1762_),
    .A2(_1779_));
 sg13g2_nor2_2 _6165_ (.A(net2042),
    .B(net1984),
    .Y(_1781_));
 sg13g2_nand2_2 _6166_ (.Y(_1782_),
    .A(net2188),
    .B(net1985));
 sg13g2_a21oi_1 _6167_ (.A1(_1778_),
    .A2(_1781_),
    .Y(_1783_),
    .B1(net2049));
 sg13g2_nor2_2 _6168_ (.A(net2044),
    .B(_1579_),
    .Y(_1784_));
 sg13g2_o21ai_1 _6169_ (.B1(net1796),
    .Y(_1785_),
    .A1(net2244),
    .A2(net1805));
 sg13g2_o21ai_1 _6170_ (.B1(net2218),
    .Y(_1786_),
    .A1(net2226),
    .A2(net1805));
 sg13g2_a22oi_1 _6171_ (.Y(_1787_),
    .B1(_1786_),
    .B2(_1776_),
    .A2(_1785_),
    .A1(_1784_));
 sg13g2_a221oi_1 _6172_ (.B2(net2050),
    .C1(net1896),
    .B1(_1787_),
    .A1(_1780_),
    .Y(_1788_),
    .A2(_1783_));
 sg13g2_o21ai_1 _6173_ (.B1(_1747_),
    .Y(_1789_),
    .A1(_1774_),
    .A2(_1788_));
 sg13g2_and2_1 _6174_ (.A(_1462_),
    .B(_1697_),
    .X(_1790_));
 sg13g2_o21ai_1 _6175_ (.B1(net2214),
    .Y(_1791_),
    .A1(net2142),
    .A2(_1722_));
 sg13g2_nand2_1 _6176_ (.Y(_1792_),
    .A(net1910),
    .B(_1791_));
 sg13g2_a21oi_1 _6177_ (.A1(net2243),
    .A2(net1954),
    .Y(_1793_),
    .B1(_1556_));
 sg13g2_a221oi_1 _6178_ (.B2(net2031),
    .C1(_1792_),
    .B1(_1793_),
    .A1(net1956),
    .Y(_1794_),
    .A2(net1873));
 sg13g2_nor2_2 _6179_ (.A(net2247),
    .B(net2025),
    .Y(_1795_));
 sg13g2_nand2b_2 _6180_ (.Y(_1796_),
    .B(net2137),
    .A_N(net2243));
 sg13g2_o21ai_1 _6181_ (.B1(_1728_),
    .Y(_1797_),
    .A1(net2138),
    .A2(net1876));
 sg13g2_nand3_1 _6182_ (.B(_1796_),
    .C(_1797_),
    .A(net2214),
    .Y(_1798_));
 sg13g2_nand2_2 _6183_ (.Y(_1799_),
    .A(net2138),
    .B(_1494_));
 sg13g2_a21oi_1 _6184_ (.A1(net1842),
    .A2(_1799_),
    .Y(_1800_),
    .B1(net2214));
 sg13g2_nor2_1 _6185_ (.A(net1890),
    .B(_1800_),
    .Y(_1801_));
 sg13g2_and2_1 _6186_ (.A(net2230),
    .B(net1973),
    .X(_1802_));
 sg13g2_nand2_2 _6187_ (.Y(_1803_),
    .A(net2243),
    .B(net1973));
 sg13g2_nand3_1 _6188_ (.B(_1797_),
    .C(_1803_),
    .A(net2214),
    .Y(_1804_));
 sg13g2_a21oi_1 _6189_ (.A1(net2142),
    .A2(net2146),
    .Y(_1805_),
    .B1(_1633_));
 sg13g2_nor2_1 _6190_ (.A(net2207),
    .B(_1805_),
    .Y(_1806_));
 sg13g2_nor2_2 _6191_ (.A(net1857),
    .B(_1806_),
    .Y(_1807_));
 sg13g2_a221oi_1 _6192_ (.B2(_1807_),
    .C1(_1794_),
    .B1(_1804_),
    .A1(_1798_),
    .Y(_1808_),
    .A2(_1801_));
 sg13g2_nor2_1 _6193_ (.A(net1896),
    .B(_1808_),
    .Y(_1809_));
 sg13g2_nor2_2 _6194_ (.A(_0091_),
    .B(net1938),
    .Y(_1810_));
 sg13g2_nand2b_2 _6195_ (.Y(_1811_),
    .B(net1942),
    .A_N(_0091_));
 sg13g2_nor2_1 _6196_ (.A(_1551_),
    .B(_1737_),
    .Y(_1812_));
 sg13g2_a22oi_1 _6197_ (.Y(_1813_),
    .B1(_1812_),
    .B2(_1616_),
    .A2(net1846),
    .A1(net1800));
 sg13g2_nor2_1 _6198_ (.A(net2140),
    .B(_1768_),
    .Y(_1814_));
 sg13g2_nand2b_2 _6199_ (.Y(_1815_),
    .B(net2021),
    .A_N(_1768_));
 sg13g2_nor2_2 _6200_ (.A(net2229),
    .B(net1834),
    .Y(_1816_));
 sg13g2_a21oi_1 _6201_ (.A1(net1989),
    .A2(_1815_),
    .Y(_1817_),
    .B1(net1811));
 sg13g2_or2_2 _6202_ (.X(_1818_),
    .B(net2130),
    .A(net2147));
 sg13g2_a22oi_1 _6203_ (.Y(_1819_),
    .B1(_1818_),
    .B2(net1913),
    .A2(_1817_),
    .A1(net2042));
 sg13g2_a21oi_1 _6204_ (.A1(_1813_),
    .A2(_1819_),
    .Y(_1820_),
    .B1(_1811_));
 sg13g2_o21ai_1 _6205_ (.B1(net1729),
    .Y(_1821_),
    .A1(_1809_),
    .A2(_1820_));
 sg13g2_and2_1 _6206_ (.A(_1462_),
    .B(_1667_),
    .X(_1822_));
 sg13g2_nand2_1 _6207_ (.Y(_1823_),
    .A(net2024),
    .B(_0096_));
 sg13g2_nand2_1 _6208_ (.Y(_1824_),
    .A(net1789),
    .B(net1833));
 sg13g2_a22oi_1 _6209_ (.Y(_1825_),
    .B1(_1824_),
    .B2(net1966),
    .A2(net1848),
    .A1(net1975));
 sg13g2_inv_1 _6210_ (.Y(_1826_),
    .A(_1825_));
 sg13g2_nand2_2 _6211_ (.Y(_1827_),
    .A(net2134),
    .B(_0096_));
 sg13g2_o21ai_1 _6212_ (.B1(_1827_),
    .Y(_1828_),
    .A1(net2134),
    .A2(net1876));
 sg13g2_nor2b_1 _6213_ (.A(net2231),
    .B_N(_1828_),
    .Y(_1829_));
 sg13g2_a21o_1 _6214_ (.A2(net1975),
    .A1(net2231),
    .B1(_1829_),
    .X(_1830_));
 sg13g2_a21oi_2 _6215_ (.B1(net2172),
    .Y(_1831_),
    .A2(_1828_),
    .A1(net1846));
 sg13g2_a21oi_1 _6216_ (.A1(net2026),
    .A2(net1974),
    .Y(_1832_),
    .B1(net1971));
 sg13g2_o21ai_1 _6217_ (.B1(_1831_),
    .Y(_1833_),
    .A1(_1670_),
    .A2(_1832_));
 sg13g2_a221oi_1 _6218_ (.B2(net1912),
    .C1(_1833_),
    .B1(_1830_),
    .A1(net2188),
    .Y(_1834_),
    .A2(_1826_));
 sg13g2_a21oi_1 _6219_ (.A1(net1789),
    .A2(net1833),
    .Y(_1835_),
    .B1(net1981));
 sg13g2_nor2_2 _6220_ (.A(net1874),
    .B(net1868),
    .Y(_1836_));
 sg13g2_nand2_2 _6221_ (.Y(_1837_),
    .A(net1947),
    .B(_1836_));
 sg13g2_nor2_1 _6222_ (.A(net2130),
    .B(_1519_),
    .Y(_1838_));
 sg13g2_nor2_1 _6223_ (.A(net2029),
    .B(_1838_),
    .Y(_1839_));
 sg13g2_o21ai_1 _6224_ (.B1(net1908),
    .Y(_1840_),
    .A1(_1521_),
    .A2(_1837_));
 sg13g2_nor3_1 _6225_ (.A(_1835_),
    .B(_1839_),
    .C(_1840_),
    .Y(_1841_));
 sg13g2_o21ai_1 _6226_ (.B1(net1899),
    .Y(_1842_),
    .A1(_1834_),
    .A2(_1841_));
 sg13g2_nand2_2 _6227_ (.Y(_1843_),
    .A(net2245),
    .B(_1595_));
 sg13g2_nand2_1 _6228_ (.Y(_1844_),
    .A(net2219),
    .B(_1843_));
 sg13g2_nand3b_1 _6229_ (.B(_1592_),
    .C(net1833),
    .Y(_1845_),
    .A_N(net2235));
 sg13g2_nand3_1 _6230_ (.B(_1843_),
    .C(_1845_),
    .A(net2208),
    .Y(_1846_));
 sg13g2_o21ai_1 _6231_ (.B1(_1728_),
    .Y(_1847_),
    .A1(net2138),
    .A2(net1880));
 sg13g2_a22oi_1 _6232_ (.Y(_1848_),
    .B1(_1847_),
    .B2(net1956),
    .A2(net1838),
    .A1(net1986));
 sg13g2_a21oi_1 _6233_ (.A1(_1846_),
    .A2(_1848_),
    .Y(_1849_),
    .B1(net2189));
 sg13g2_nand2_2 _6234_ (.Y(_1850_),
    .A(net1974),
    .B(net1950));
 sg13g2_nor2_2 _6235_ (.A(net1810),
    .B(net1868),
    .Y(_1851_));
 sg13g2_nor2_1 _6236_ (.A(_1521_),
    .B(_1805_),
    .Y(_1852_));
 sg13g2_a221oi_1 _6237_ (.B2(net1986),
    .C1(_1852_),
    .B1(_1851_),
    .A1(net2207),
    .Y(_1853_),
    .A2(_1797_));
 sg13g2_o21ai_1 _6238_ (.B1(_1810_),
    .Y(_1854_),
    .A1(net2040),
    .A2(_1853_));
 sg13g2_o21ai_1 _6239_ (.B1(_1842_),
    .Y(_1855_),
    .A1(_1849_),
    .A2(_1854_));
 sg13g2_and2_1 _6240_ (.A(net1742),
    .B(_1855_),
    .X(_1856_));
 sg13g2_nand3_1 _6241_ (.B(_1462_),
    .C(_1474_),
    .A(_1450_),
    .Y(_1857_));
 sg13g2_nor2_1 _6242_ (.A(net2132),
    .B(net1810),
    .Y(_1858_));
 sg13g2_nand2b_2 _6243_ (.Y(_1859_),
    .B(net1807),
    .A_N(net2132));
 sg13g2_nand2_2 _6244_ (.Y(_1860_),
    .A(net2229),
    .B(net1869));
 sg13g2_and2_2 _6245_ (.A(net2227),
    .B(net1869),
    .X(_1861_));
 sg13g2_nor2_1 _6246_ (.A(net2201),
    .B(_1861_),
    .Y(_1862_));
 sg13g2_nor2_2 _6247_ (.A(net1973),
    .B(_1536_),
    .Y(_1863_));
 sg13g2_nand2_2 _6248_ (.Y(_1864_),
    .A(_1402_),
    .B(_1850_));
 sg13g2_nand2_1 _6249_ (.Y(_1865_),
    .A(_1558_),
    .B(_1864_));
 sg13g2_a21oi_1 _6250_ (.A1(net1804),
    .A2(_1816_),
    .Y(_1866_),
    .B1(net2202));
 sg13g2_nand2_1 _6251_ (.Y(_1867_),
    .A(net2203),
    .B(_1850_));
 sg13g2_a22oi_1 _6252_ (.Y(_1868_),
    .B1(_1865_),
    .B2(_1866_),
    .A2(_1863_),
    .A1(net2202));
 sg13g2_nand2_1 _6253_ (.Y(_1869_),
    .A(_1717_),
    .B(_1758_));
 sg13g2_o21ai_1 _6254_ (.B1(net1839),
    .Y(_1870_),
    .A1(net1796),
    .A2(_1869_));
 sg13g2_nor2_1 _6255_ (.A(net1904),
    .B(_1748_),
    .Y(_1871_));
 sg13g2_nand2_2 _6256_ (.Y(_1872_),
    .A(net1907),
    .B(net1841));
 sg13g2_o21ai_1 _6257_ (.B1(_1749_),
    .Y(_1873_),
    .A1(net1965),
    .A2(net1837));
 sg13g2_nor2_1 _6258_ (.A(net1904),
    .B(_1873_),
    .Y(_1874_));
 sg13g2_a21oi_1 _6259_ (.A1(net1851),
    .A2(_1868_),
    .Y(_1875_),
    .B1(_1874_));
 sg13g2_a21oi_1 _6260_ (.A1(net2234),
    .A2(net1947),
    .Y(_1876_),
    .B1(net2208));
 sg13g2_o21ai_1 _6261_ (.B1(_1876_),
    .Y(_1877_),
    .A1(net2234),
    .A2(_1729_));
 sg13g2_nand2b_1 _6262_ (.Y(_1878_),
    .B(net1947),
    .A_N(net2232));
 sg13g2_nand2_2 _6263_ (.Y(_1879_),
    .A(net2207),
    .B(_1769_));
 sg13g2_nand2b_2 _6264_ (.Y(_1880_),
    .B(_1879_),
    .A_N(net1847));
 sg13g2_a21oi_1 _6265_ (.A1(_1878_),
    .A2(_1880_),
    .Y(_1881_),
    .B1(net2039));
 sg13g2_nand2_1 _6266_ (.Y(_1882_),
    .A(_1877_),
    .B(_1881_));
 sg13g2_nor2_1 _6267_ (.A(_1594_),
    .B(_1764_),
    .Y(_1883_));
 sg13g2_nor2_1 _6268_ (.A(_1838_),
    .B(_1883_),
    .Y(_1884_));
 sg13g2_a22oi_1 _6269_ (.Y(_1885_),
    .B1(_1884_),
    .B2(net1927),
    .A2(_1730_),
    .A1(net1912));
 sg13g2_a21oi_1 _6270_ (.A1(_1882_),
    .A2(_1885_),
    .Y(_1886_),
    .B1(net2173));
 sg13g2_o21ai_1 _6271_ (.B1(net1851),
    .Y(_1887_),
    .A1(net1982),
    .A2(_1837_));
 sg13g2_nand2_2 _6272_ (.Y(_1888_),
    .A(net1899),
    .B(_1887_));
 sg13g2_nand2b_2 _6273_ (.Y(_1889_),
    .B(net1884),
    .A_N(net2130));
 sg13g2_nor2_1 _6274_ (.A(net2130),
    .B(net1809),
    .Y(_1890_));
 sg13g2_nand2b_2 _6275_ (.Y(_1891_),
    .B(net1811),
    .A_N(net2133));
 sg13g2_nor2_2 _6276_ (.A(net2234),
    .B(_1890_),
    .Y(_1892_));
 sg13g2_a21oi_1 _6277_ (.A1(net1982),
    .A2(_1684_),
    .Y(_1893_),
    .B1(_1892_));
 sg13g2_a22oi_1 _6278_ (.Y(_1894_),
    .B1(_1577_),
    .B2(net1961),
    .A2(net1867),
    .A1(net1892));
 sg13g2_nor3_1 _6279_ (.A(net1904),
    .B(_1893_),
    .C(_1894_),
    .Y(_1895_));
 sg13g2_nor3_1 _6280_ (.A(_1886_),
    .B(_1888_),
    .C(_1895_),
    .Y(_1896_));
 sg13g2_a21oi_1 _6281_ (.A1(_1870_),
    .A2(_1875_),
    .Y(_1897_),
    .B1(_1896_));
 sg13g2_nor2_1 _6282_ (.A(_1857_),
    .B(_1897_),
    .Y(_1898_));
 sg13g2_nand2b_2 _6283_ (.Y(_1899_),
    .B(_1667_),
    .A_N(_1464_));
 sg13g2_nand2_2 _6284_ (.Y(_1900_),
    .A(net2142),
    .B(_1550_));
 sg13g2_nand2_2 _6285_ (.Y(_1901_),
    .A(net2136),
    .B(net1810));
 sg13g2_nand2_2 _6286_ (.Y(_1902_),
    .A(net1869),
    .B(net1789));
 sg13g2_inv_1 _6287_ (.Y(_1903_),
    .A(_1902_));
 sg13g2_nor2_1 _6288_ (.A(_1521_),
    .B(_1902_),
    .Y(_1904_));
 sg13g2_a21oi_2 _6289_ (.B1(_1904_),
    .Y(_1905_),
    .A2(net1787),
    .A1(net1987));
 sg13g2_nand2_1 _6290_ (.Y(_1906_),
    .A(net2223),
    .B(_1859_));
 sg13g2_a21oi_1 _6291_ (.A1(_1905_),
    .A2(_1906_),
    .Y(_1907_),
    .B1(net1906));
 sg13g2_nand2_1 _6292_ (.Y(_1908_),
    .A(net2227),
    .B(net1787));
 sg13g2_nand2_2 _6293_ (.Y(_1909_),
    .A(net1968),
    .B(net1787));
 sg13g2_nand2_1 _6294_ (.Y(_1910_),
    .A(net1964),
    .B(_1595_));
 sg13g2_a21oi_1 _6295_ (.A1(_1909_),
    .A2(_1910_),
    .Y(_1911_),
    .B1(net1857));
 sg13g2_nand2b_2 _6296_ (.Y(_1912_),
    .B(net1884),
    .A_N(net2241));
 sg13g2_nor2_2 _6297_ (.A(_1484_),
    .B(_1519_),
    .Y(_1913_));
 sg13g2_a21oi_1 _6298_ (.A1(net1808),
    .A2(_1715_),
    .Y(_1914_),
    .B1(net1936));
 sg13g2_o21ai_1 _6299_ (.B1(_1914_),
    .Y(_1915_),
    .A1(_1844_),
    .A2(_1913_));
 sg13g2_nor2_1 _6300_ (.A(_1514_),
    .B(_1553_),
    .Y(_1916_));
 sg13g2_nor2_2 _6301_ (.A(net2226),
    .B(_1512_),
    .Y(_1917_));
 sg13g2_nor2_1 _6302_ (.A(net2219),
    .B(_1917_),
    .Y(_1918_));
 sg13g2_nor2_1 _6303_ (.A(_1916_),
    .B(_1918_),
    .Y(_1919_));
 sg13g2_o21ai_1 _6304_ (.B1(_1915_),
    .Y(_1920_),
    .A1(net1890),
    .A2(_1919_));
 sg13g2_nor4_1 _6305_ (.A(net1939),
    .B(_1907_),
    .C(_1911_),
    .D(_1920_),
    .Y(_1921_));
 sg13g2_nand2_2 _6306_ (.Y(_1922_),
    .A(net2236),
    .B(net1804));
 sg13g2_o21ai_1 _6307_ (.B1(_1922_),
    .Y(_1923_),
    .A1(_1519_),
    .A2(net1801));
 sg13g2_a21oi_1 _6308_ (.A1(_1509_),
    .A2(_1923_),
    .Y(_1924_),
    .B1(net1887));
 sg13g2_nand2_1 _6309_ (.Y(_1925_),
    .A(net2158),
    .B(net1813));
 sg13g2_nor2_2 _6310_ (.A(net1887),
    .B(net1948),
    .Y(_1926_));
 sg13g2_or2_2 _6311_ (.X(_1927_),
    .B(net1948),
    .A(net1887));
 sg13g2_a21oi_1 _6312_ (.A1(_1509_),
    .A2(_1923_),
    .Y(_1928_),
    .B1(_1927_));
 sg13g2_nor2_2 _6313_ (.A(net2245),
    .B(_1596_),
    .Y(_1929_));
 sg13g2_o21ai_1 _6314_ (.B1(_1922_),
    .Y(_1930_),
    .A1(net2240),
    .A2(_1596_));
 sg13g2_nor2_2 _6315_ (.A(net2239),
    .B(net1872),
    .Y(_1931_));
 sg13g2_nand2_2 _6316_ (.Y(_1932_),
    .A(net1870),
    .B(_1721_));
 sg13g2_nand2_2 _6317_ (.Y(_1933_),
    .A(_1865_),
    .B(_1932_));
 sg13g2_nand2_1 _6318_ (.Y(_1934_),
    .A(net1850),
    .B(_1933_));
 sg13g2_nor2_1 _6319_ (.A(net2213),
    .B(net1872),
    .Y(_1935_));
 sg13g2_nand2_1 _6320_ (.Y(_1936_),
    .A(net2029),
    .B(net1870));
 sg13g2_nor2_1 _6321_ (.A(_1563_),
    .B(_1716_),
    .Y(_1937_));
 sg13g2_a221oi_1 _6322_ (.B2(net1928),
    .C1(_1937_),
    .B1(_1930_),
    .A1(net1913),
    .Y(_1938_),
    .A2(_1900_));
 sg13g2_a21oi_1 _6323_ (.A1(_1934_),
    .A2(_1938_),
    .Y(_1939_),
    .B1(net2176));
 sg13g2_nor2_2 _6324_ (.A(net1906),
    .B(net1868),
    .Y(_1940_));
 sg13g2_o21ai_1 _6325_ (.B1(net1787),
    .Y(_1941_),
    .A1(_1393_),
    .A2(_1940_));
 sg13g2_nand2_2 _6326_ (.Y(_1942_),
    .A(net2248),
    .B(_1554_));
 sg13g2_nor2_1 _6327_ (.A(_1514_),
    .B(_1942_),
    .Y(_1943_));
 sg13g2_nand2_1 _6328_ (.Y(_1944_),
    .A(net2245),
    .B(_1916_));
 sg13g2_a21oi_1 _6329_ (.A1(net2213),
    .A2(_1929_),
    .Y(_1945_),
    .B1(_1943_));
 sg13g2_o21ai_1 _6330_ (.B1(_1941_),
    .Y(_1946_),
    .A1(net1934),
    .A2(_1945_));
 sg13g2_a21oi_1 _6331_ (.A1(_1581_),
    .A2(_1843_),
    .Y(_1947_),
    .B1(_1648_));
 sg13g2_nor4_1 _6332_ (.A(net1895),
    .B(_1939_),
    .C(_1946_),
    .D(_1947_),
    .Y(_1948_));
 sg13g2_nor3_1 _6333_ (.A(_1921_),
    .B(_1928_),
    .C(_1948_),
    .Y(_1949_));
 sg13g2_nor2_1 _6334_ (.A(_1899_),
    .B(_1949_),
    .Y(_1950_));
 sg13g2_nand2_2 _6335_ (.Y(_1951_),
    .A(_1476_),
    .B(_1697_));
 sg13g2_a21oi_1 _6336_ (.A1(net1813),
    .A2(_1674_),
    .Y(_1952_),
    .B1(net1948));
 sg13g2_nor2_1 _6337_ (.A(_1951_),
    .B(_1952_),
    .Y(_1953_));
 sg13g2_or2_1 _6338_ (.X(_1954_),
    .B(_1952_),
    .A(_1951_));
 sg13g2_nor2_2 _6339_ (.A(net2195),
    .B(net1946),
    .Y(_1955_));
 sg13g2_o21ai_1 _6340_ (.B1(net2049),
    .Y(_1956_),
    .A1(_1781_),
    .A2(_1955_));
 sg13g2_or3_1 _6341_ (.A(net2046),
    .B(_0093_),
    .C(net2183),
    .X(_1957_));
 sg13g2_a221oi_1 _6342_ (.B2(_1957_),
    .C1(net2160),
    .B1(_1956_),
    .A1(net1870),
    .Y(_1958_),
    .A2(net1864));
 sg13g2_nor2_1 _6343_ (.A(net2158),
    .B(_1958_),
    .Y(_1959_));
 sg13g2_a21oi_2 _6344_ (.B1(net1866),
    .Y(_1960_),
    .A2(net1872),
    .A1(net2238));
 sg13g2_o21ai_1 _6345_ (.B1(net1854),
    .Y(_1961_),
    .A1(net2198),
    .A2(_1960_));
 sg13g2_o21ai_1 _6346_ (.B1(net2169),
    .Y(_1962_),
    .A1(net2187),
    .A2(net1874));
 sg13g2_nor2_2 _6347_ (.A(net2190),
    .B(net1965),
    .Y(_1963_));
 sg13g2_nand2_2 _6348_ (.Y(_1964_),
    .A(net2039),
    .B(net1960));
 sg13g2_nand3_1 _6349_ (.B(net1959),
    .C(_1674_),
    .A(net1993),
    .Y(_1965_));
 sg13g2_nor2_2 _6350_ (.A(net2038),
    .B(net2198),
    .Y(_1966_));
 sg13g2_nand2_1 _6351_ (.Y(_1967_),
    .A(net1874),
    .B(_1966_));
 sg13g2_nand3_1 _6352_ (.B(_1965_),
    .C(_1967_),
    .A(_1962_),
    .Y(_1968_));
 sg13g2_a21oi_1 _6353_ (.A1(_1961_),
    .A2(_1968_),
    .Y(_1969_),
    .B1(net1893));
 sg13g2_nor3_2 _6354_ (.A(_1954_),
    .B(_1959_),
    .C(_1969_),
    .Y(_1970_));
 sg13g2_nor3_2 _6355_ (.A(_1600_),
    .B(_1666_),
    .C(_1950_),
    .Y(_1971_));
 sg13g2_and3_1 _6356_ (.X(_1972_),
    .A(_1696_),
    .B(_1789_),
    .C(_1821_));
 sg13g2_nor4_1 _6357_ (.A(net1732),
    .B(_1856_),
    .C(_1898_),
    .D(_1970_),
    .Y(_1973_));
 sg13g2_nand4_1 _6358_ (.B(_1971_),
    .C(_1972_),
    .A(_1746_),
    .Y(_1974_),
    .D(_1973_));
 sg13g2_o21ai_1 _6359_ (.B1(_1565_),
    .Y(_1975_),
    .A1(_1584_),
    .A2(_1673_));
 sg13g2_a21oi_1 _6360_ (.A1(net1865),
    .A2(net1929),
    .Y(_1976_),
    .B1(net2166));
 sg13g2_nor2_1 _6361_ (.A(net2191),
    .B(net1872),
    .Y(_1977_));
 sg13g2_nor2_1 _6362_ (.A(net1904),
    .B(net1871),
    .Y(_1978_));
 sg13g2_nor3_1 _6363_ (.A(net1893),
    .B(_1976_),
    .C(_1978_),
    .Y(_1979_));
 sg13g2_o21ai_1 _6364_ (.B1(_1927_),
    .Y(_1980_),
    .A1(net1939),
    .A2(_1956_));
 sg13g2_a22oi_1 _6365_ (.Y(_1981_),
    .B1(_1980_),
    .B2(_1674_),
    .A2(_1979_),
    .A1(_1975_));
 sg13g2_nand2_1 _6366_ (.Y(_1982_),
    .A(net1731),
    .B(_1981_));
 sg13g2_a21oi_1 _6367_ (.A1(_1974_),
    .A2(_1982_),
    .Y(_1983_),
    .B1(\draw_game_inst.board_x[1] ));
 sg13g2_nand2_2 _6368_ (.Y(_1984_),
    .A(net2192),
    .B(net1964));
 sg13g2_nor2_1 _6369_ (.A(net1804),
    .B(_1984_),
    .Y(_1985_));
 sg13g2_nor2_1 _6370_ (.A(net2238),
    .B(_1613_),
    .Y(_1986_));
 sg13g2_a21oi_2 _6371_ (.B1(_1986_),
    .Y(_1987_),
    .A2(net1864),
    .A1(net2238));
 sg13g2_inv_1 _6372_ (.Y(_1988_),
    .A(_1987_));
 sg13g2_nor3_1 _6373_ (.A(net2199),
    .B(_1802_),
    .C(_1987_),
    .Y(_1989_));
 sg13g2_nor3_1 _6374_ (.A(net1796),
    .B(_1964_),
    .C(_1989_),
    .Y(_1990_));
 sg13g2_o21ai_1 _6375_ (.B1(_1667_),
    .Y(_1991_),
    .A1(_1985_),
    .A2(_1990_));
 sg13g2_a21o_2 _6376_ (.A2(_1683_),
    .A1(net1950),
    .B1(net2188),
    .X(_1992_));
 sg13g2_nor2_2 _6377_ (.A(net2225),
    .B(net1929),
    .Y(_1993_));
 sg13g2_o21ai_1 _6378_ (.B1(net2187),
    .Y(_1994_),
    .A1(net1862),
    .A2(_1583_));
 sg13g2_nand3_1 _6379_ (.B(_1992_),
    .C(_1994_),
    .A(_1697_),
    .Y(_1995_));
 sg13g2_a21oi_1 _6380_ (.A1(_1991_),
    .A2(_1995_),
    .Y(_1996_),
    .B1(_1811_));
 sg13g2_nand2_1 _6381_ (.Y(_1997_),
    .A(net2131),
    .B(net1847));
 sg13g2_nand3_1 _6382_ (.B(net1885),
    .C(_1997_),
    .A(net1908),
    .Y(_1998_));
 sg13g2_nand2_1 _6383_ (.Y(_1999_),
    .A(net1843),
    .B(_1901_));
 sg13g2_a21oi_2 _6384_ (.B1(net2244),
    .Y(_2000_),
    .A2(_1901_),
    .A1(net1843));
 sg13g2_o21ai_1 _6385_ (.B1(net1843),
    .Y(_2001_),
    .A1(net2025),
    .A2(net1881));
 sg13g2_a21oi_1 _6386_ (.A1(net2245),
    .A2(net1795),
    .Y(_2002_),
    .B1(_2000_));
 sg13g2_o21ai_1 _6387_ (.B1(net2180),
    .Y(_2003_),
    .A1(net1931),
    .A2(_1929_));
 sg13g2_a21oi_2 _6388_ (.B1(_2003_),
    .Y(_2004_),
    .A2(_2002_),
    .A1(net1845));
 sg13g2_a21oi_1 _6389_ (.A1(net1789),
    .A2(_1710_),
    .Y(_2005_),
    .B1(net2184));
 sg13g2_a22oi_1 _6390_ (.Y(_2006_),
    .B1(_1837_),
    .B2(_1480_),
    .A2(net1966),
    .A1(net1884));
 sg13g2_o21ai_1 _6391_ (.B1(_2006_),
    .Y(_2007_),
    .A1(net2171),
    .A2(_2005_));
 sg13g2_o21ai_1 _6392_ (.B1(_1998_),
    .Y(_2008_),
    .A1(_2004_),
    .A2(_2007_));
 sg13g2_nand2_1 _6393_ (.Y(_2009_),
    .A(net1892),
    .B(net1789));
 sg13g2_nand3_1 _6394_ (.B(net1789),
    .C(_1861_),
    .A(net1892),
    .Y(_2010_));
 sg13g2_o21ai_1 _6395_ (.B1(_2010_),
    .Y(_2011_),
    .A1(net2227),
    .A2(net1788));
 sg13g2_nor2_2 _6396_ (.A(net2241),
    .B(net1952),
    .Y(_2012_));
 sg13g2_o21ai_1 _6397_ (.B1(net2201),
    .Y(_2013_),
    .A1(net2228),
    .A2(net1954));
 sg13g2_a21oi_2 _6398_ (.B1(_2013_),
    .Y(_2014_),
    .A2(_1763_),
    .A1(net1879));
 sg13g2_nor3_1 _6399_ (.A(net2143),
    .B(_1497_),
    .C(_2014_),
    .Y(_2015_));
 sg13g2_nand2_1 _6400_ (.Y(_2016_),
    .A(net2227),
    .B(_1815_));
 sg13g2_a21oi_1 _6401_ (.A1(_1650_),
    .A2(_2016_),
    .Y(_2017_),
    .B1(net2201));
 sg13g2_nor2_2 _6402_ (.A(net2166),
    .B(_1686_),
    .Y(_2018_));
 sg13g2_nand2_2 _6403_ (.Y(_2019_),
    .A(_1402_),
    .B(_1713_));
 sg13g2_a221oi_1 _6404_ (.B2(_2019_),
    .C1(_1888_),
    .B1(_2018_),
    .A1(_1871_),
    .Y(_2020_),
    .A2(_2017_));
 sg13g2_o21ai_1 _6405_ (.B1(_2020_),
    .Y(_2021_),
    .A1(net1888),
    .A2(_2015_));
 sg13g2_a21oi_1 _6406_ (.A1(_1393_),
    .A2(_2011_),
    .Y(_2022_),
    .B1(_2021_));
 sg13g2_a21oi_1 _6407_ (.A1(net1942),
    .A2(_2008_),
    .Y(_2023_),
    .B1(_2022_));
 sg13g2_nor2_2 _6408_ (.A(net1902),
    .B(net1966),
    .Y(_2024_));
 sg13g2_nand2_2 _6409_ (.Y(_2025_),
    .A(net1910),
    .B(net1963));
 sg13g2_nand2_2 _6410_ (.Y(_2026_),
    .A(_1574_),
    .B(net1794));
 sg13g2_a21oi_1 _6411_ (.A1(net2199),
    .A2(net1862),
    .Y(_2027_),
    .B1(net2167));
 sg13g2_nor2_1 _6412_ (.A(net2183),
    .B(_1583_),
    .Y(_2028_));
 sg13g2_nand3_1 _6413_ (.B(_2027_),
    .C(_2028_),
    .A(_1716_),
    .Y(_2029_));
 sg13g2_o21ai_1 _6414_ (.B1(_2029_),
    .Y(_2030_),
    .A1(net1800),
    .A2(_2026_));
 sg13g2_nand2_1 _6415_ (.Y(_2031_),
    .A(net2188),
    .B(_1684_));
 sg13g2_nor2_2 _6416_ (.A(net2199),
    .B(net1804),
    .Y(_2032_));
 sg13g2_nand2_1 _6417_ (.Y(_2033_),
    .A(net2035),
    .B(net1806));
 sg13g2_nor2_2 _6418_ (.A(net2186),
    .B(_2032_),
    .Y(_2034_));
 sg13g2_nor2_1 _6419_ (.A(net2167),
    .B(_2034_),
    .Y(_2035_));
 sg13g2_o21ai_1 _6420_ (.B1(_2035_),
    .Y(_2036_),
    .A1(_1761_),
    .A2(_2031_));
 sg13g2_nor3_1 _6421_ (.A(net2045),
    .B(net1965),
    .C(net1945),
    .Y(_2037_));
 sg13g2_nand3_1 _6422_ (.B(net1950),
    .C(_2037_),
    .A(net2028),
    .Y(_2038_));
 sg13g2_a21oi_1 _6423_ (.A1(_2036_),
    .A2(_2038_),
    .Y(_2039_),
    .B1(net1851));
 sg13g2_a22oi_1 _6424_ (.Y(_2040_),
    .B1(_2039_),
    .B2(_1697_),
    .A2(_2030_),
    .A1(_1667_));
 sg13g2_nand2b_1 _6425_ (.Y(_2041_),
    .B(net1898),
    .A_N(_2040_));
 sg13g2_o21ai_1 _6426_ (.B1(_2041_),
    .Y(_2042_),
    .A1(_1601_),
    .A2(_2023_));
 sg13g2_o21ai_1 _6427_ (.B1(_1462_),
    .Y(_2043_),
    .A1(_1996_),
    .A2(_2042_));
 sg13g2_nand2_2 _6428_ (.Y(_2044_),
    .A(net2164),
    .B(net1813));
 sg13g2_nor2_2 _6429_ (.A(net1807),
    .B(_1722_),
    .Y(_2045_));
 sg13g2_a221oi_1 _6430_ (.B2(_1818_),
    .C1(_2044_),
    .B1(_1763_),
    .A1(net1810),
    .Y(_2046_),
    .A2(_1721_));
 sg13g2_nor2_2 _6431_ (.A(net2219),
    .B(net1874),
    .Y(_2047_));
 sg13g2_nand2_2 _6432_ (.Y(_2048_),
    .A(net2035),
    .B(_1509_));
 sg13g2_nor2b_1 _6433_ (.A(_2047_),
    .B_N(_1955_),
    .Y(_2049_));
 sg13g2_a21oi_1 _6434_ (.A1(net2244),
    .A2(_1570_),
    .Y(_2050_),
    .B1(net1875));
 sg13g2_nand2_1 _6435_ (.Y(_2051_),
    .A(net2218),
    .B(_2050_));
 sg13g2_nand2_1 _6436_ (.Y(_2052_),
    .A(net2218),
    .B(_1815_));
 sg13g2_nor2_2 _6437_ (.A(net1988),
    .B(net1836),
    .Y(_2053_));
 sg13g2_nand2b_1 _6438_ (.Y(_2054_),
    .B(_1572_),
    .A_N(net2240));
 sg13g2_a21oi_1 _6439_ (.A1(net1988),
    .A2(_1572_),
    .Y(_2055_),
    .B1(_2053_));
 sg13g2_a221oi_1 _6440_ (.B2(net2195),
    .C1(net2180),
    .B1(_2055_),
    .A1(_2049_),
    .Y(_2056_),
    .A2(_2051_));
 sg13g2_o21ai_1 _6441_ (.B1(net2211),
    .Y(_2057_),
    .A1(_1560_),
    .A2(_1986_));
 sg13g2_nor2_1 _6442_ (.A(net2218),
    .B(net1972),
    .Y(_2058_));
 sg13g2_nand2_1 _6443_ (.Y(_2059_),
    .A(_1803_),
    .B(_2058_));
 sg13g2_a21oi_1 _6444_ (.A1(_2057_),
    .A2(_2059_),
    .Y(_2060_),
    .B1(net1935));
 sg13g2_nor2_1 _6445_ (.A(net2228),
    .B(_1815_),
    .Y(_2061_));
 sg13g2_o21ai_1 _6446_ (.B1(_1775_),
    .Y(_2062_),
    .A1(net2244),
    .A2(_1815_));
 sg13g2_o21ai_1 _6447_ (.B1(_1644_),
    .Y(_2063_),
    .A1(net1967),
    .A2(net1796));
 sg13g2_a21oi_1 _6448_ (.A1(_2062_),
    .A2(_2063_),
    .Y(_2064_),
    .B1(net1905));
 sg13g2_nor4_2 _6449_ (.A(net2164),
    .B(_2056_),
    .C(_2060_),
    .Y(_2065_),
    .D(_2064_));
 sg13g2_o21ai_1 _6450_ (.B1(net1743),
    .Y(_2066_),
    .A1(_2046_),
    .A2(_2065_));
 sg13g2_a21oi_1 _6451_ (.A1(net1969),
    .A2(net1804),
    .Y(_2067_),
    .B1(net2194));
 sg13g2_o21ai_1 _6452_ (.B1(_2067_),
    .Y(_2068_),
    .A1(net1976),
    .A2(net1969));
 sg13g2_nor2_1 _6453_ (.A(net2176),
    .B(_2068_),
    .Y(_2069_));
 sg13g2_nor2_2 _6454_ (.A(net2218),
    .B(_1491_),
    .Y(_2070_));
 sg13g2_nor3_1 _6455_ (.A(net2033),
    .B(_1651_),
    .C(_1836_),
    .Y(_2071_));
 sg13g2_o21ai_1 _6456_ (.B1(net1853),
    .Y(_2072_),
    .A1(_2070_),
    .A2(_2071_));
 sg13g2_a21oi_1 _6457_ (.A1(_1513_),
    .A2(net1934),
    .Y(_2073_),
    .B1(_2069_));
 sg13g2_a21oi_1 _6458_ (.A1(_2072_),
    .A2(_2073_),
    .Y(_2074_),
    .B1(net2163));
 sg13g2_a221oi_1 _6459_ (.B2(net1951),
    .C1(_2044_),
    .B1(_1654_),
    .A1(net2239),
    .Y(_2075_),
    .A2(_1572_));
 sg13g2_o21ai_1 _6460_ (.B1(net1730),
    .Y(_2076_),
    .A1(_2074_),
    .A2(_2075_));
 sg13g2_a21oi_2 _6461_ (.B1(net2052),
    .Y(_2077_),
    .A2(_2076_),
    .A1(_2066_));
 sg13g2_nor2_1 _6462_ (.A(_1748_),
    .B(net1834),
    .Y(_2078_));
 sg13g2_nand2_1 _6463_ (.Y(_2079_),
    .A(net1841),
    .B(_1815_));
 sg13g2_a221oi_1 _6464_ (.B2(net1965),
    .C1(net2183),
    .B1(_2078_),
    .A1(net1847),
    .Y(_2080_),
    .A2(_1859_));
 sg13g2_a21o_1 _6465_ (.A2(_2080_),
    .A1(_1905_),
    .B1(net2170),
    .X(_2081_));
 sg13g2_o21ai_1 _6466_ (.B1(_1940_),
    .Y(_2082_),
    .A1(net2210),
    .A2(_1749_));
 sg13g2_nor3_1 _6467_ (.A(net2032),
    .B(net1806),
    .C(_2061_),
    .Y(_2083_));
 sg13g2_o21ai_1 _6468_ (.B1(net1854),
    .Y(_2084_),
    .A1(_2017_),
    .A2(_2083_));
 sg13g2_and4_1 _6469_ (.A(net1942),
    .B(_2081_),
    .C(_2082_),
    .D(_2084_),
    .X(_2085_));
 sg13g2_nand2_2 _6470_ (.Y(_2086_),
    .A(net2227),
    .B(net1802));
 sg13g2_nor2b_1 _6471_ (.A(_1816_),
    .B_N(_2086_),
    .Y(_2087_));
 sg13g2_and2_1 _6472_ (.A(_1545_),
    .B(_1799_),
    .X(_2088_));
 sg13g2_nand2_2 _6473_ (.Y(_2089_),
    .A(net1985),
    .B(net1851));
 sg13g2_a21oi_1 _6474_ (.A1(net1883),
    .A2(net1958),
    .Y(_2090_),
    .B1(_2089_));
 sg13g2_a221oi_1 _6475_ (.B2(net1833),
    .C1(_2090_),
    .B1(_2088_),
    .A1(net1836),
    .Y(_2091_),
    .A2(_2024_));
 sg13g2_nand2b_1 _6476_ (.Y(_2092_),
    .B(net1803),
    .A_N(net2228));
 sg13g2_nor2_2 _6477_ (.A(net2032),
    .B(_1931_),
    .Y(_2093_));
 sg13g2_a22oi_1 _6478_ (.Y(_2094_),
    .B1(_2093_),
    .B2(_2016_),
    .A2(_2092_),
    .A1(_1862_));
 sg13g2_nor2_1 _6479_ (.A(net2041),
    .B(_2094_),
    .Y(_2095_));
 sg13g2_a221oi_1 _6480_ (.B2(net1912),
    .C1(_2095_),
    .B1(_2087_),
    .A1(net1927),
    .Y(_2096_),
    .A2(net1788));
 sg13g2_o21ai_1 _6481_ (.B1(_2091_),
    .Y(_2097_),
    .A1(net2170),
    .A2(_2096_));
 sg13g2_a21oi_1 _6482_ (.A1(net1898),
    .A2(_2097_),
    .Y(_2098_),
    .B1(_2085_));
 sg13g2_nor2b_1 _6483_ (.A(_2098_),
    .B_N(_1698_),
    .Y(_2099_));
 sg13g2_nand2_1 _6484_ (.Y(_2100_),
    .A(net2039),
    .B(net1873));
 sg13g2_o21ai_1 _6485_ (.B1(net2167),
    .Y(_2101_),
    .A1(net1869),
    .A2(_1964_));
 sg13g2_nor2_2 _6486_ (.A(_1506_),
    .B(net1866),
    .Y(_2102_));
 sg13g2_nand2_1 _6487_ (.Y(_2103_),
    .A(net1958),
    .B(net1861));
 sg13g2_nor2_1 _6488_ (.A(_1654_),
    .B(_2102_),
    .Y(_2104_));
 sg13g2_nor3_2 _6489_ (.A(net2042),
    .B(net1946),
    .C(_2047_),
    .Y(_2105_));
 sg13g2_o21ai_1 _6490_ (.B1(_2105_),
    .Y(_2106_),
    .A1(net2032),
    .A2(_2104_));
 sg13g2_nand2b_1 _6491_ (.Y(_2107_),
    .B(_2106_),
    .A_N(_2101_));
 sg13g2_nand2_2 _6492_ (.Y(_2108_),
    .A(net1983),
    .B(net1872));
 sg13g2_a22oi_1 _6493_ (.Y(_2109_),
    .B1(_2108_),
    .B2(net1858),
    .A2(_1685_),
    .A1(net1991));
 sg13g2_a21oi_1 _6494_ (.A1(_2107_),
    .A2(_2109_),
    .Y(_2110_),
    .B1(net1893));
 sg13g2_a21oi_2 _6495_ (.B1(net1949),
    .Y(_2111_),
    .A2(_2103_),
    .A1(net1813));
 sg13g2_nand2_2 _6496_ (.Y(_2112_),
    .A(net2211),
    .B(net1866));
 sg13g2_and2_1 _6497_ (.A(_2108_),
    .B(_2112_),
    .X(_2113_));
 sg13g2_a21oi_2 _6498_ (.B1(net2160),
    .Y(_2114_),
    .A2(_2113_),
    .A1(net1993));
 sg13g2_a21oi_1 _6499_ (.A1(net1874),
    .A2(_1963_),
    .Y(_2115_),
    .B1(_1678_));
 sg13g2_a221oi_1 _6500_ (.B2(net1863),
    .C1(_2115_),
    .B1(net1798),
    .A1(net1800),
    .Y(_2116_),
    .A2(_1623_));
 sg13g2_a21oi_1 _6501_ (.A1(_2114_),
    .A2(_2116_),
    .Y(_2117_),
    .B1(net2156));
 sg13g2_nor3_1 _6502_ (.A(_2110_),
    .B(_2111_),
    .C(_2117_),
    .Y(_2118_));
 sg13g2_a21oi_1 _6503_ (.A1(net2142),
    .A2(_1549_),
    .Y(_2119_),
    .B1(net1963));
 sg13g2_a22oi_1 _6504_ (.Y(_2120_),
    .B1(_2119_),
    .B2(_1552_),
    .A2(_1703_),
    .A1(net1961));
 sg13g2_a21oi_1 _6505_ (.A1(_1506_),
    .A2(net1927),
    .Y(_2121_),
    .B1(_1678_));
 sg13g2_nand3_1 _6506_ (.B(_1652_),
    .C(_2103_),
    .A(net2200),
    .Y(_2122_));
 sg13g2_o21ai_1 _6507_ (.B1(_2122_),
    .Y(_2123_),
    .A1(net2200),
    .A2(net1800));
 sg13g2_nor2_1 _6508_ (.A(net2166),
    .B(_2123_),
    .Y(_2124_));
 sg13g2_nor2_1 _6509_ (.A(_2121_),
    .B(_2124_),
    .Y(_2125_));
 sg13g2_o21ai_1 _6510_ (.B1(_2125_),
    .Y(_2126_),
    .A1(net1888),
    .A2(_2120_));
 sg13g2_nor2_2 _6511_ (.A(net1861),
    .B(net1945),
    .Y(_2127_));
 sg13g2_nor2_1 _6512_ (.A(net2186),
    .B(_2127_),
    .Y(_2128_));
 sg13g2_a21oi_1 _6513_ (.A1(_1544_),
    .A2(net1862),
    .Y(_2129_),
    .B1(_2128_));
 sg13g2_nand2_1 _6514_ (.Y(_2130_),
    .A(net1871),
    .B(net1929));
 sg13g2_nor2b_1 _6515_ (.A(_1678_),
    .B_N(_2130_),
    .Y(_2131_));
 sg13g2_nor2_1 _6516_ (.A(net2161),
    .B(_2131_),
    .Y(_2132_));
 sg13g2_o21ai_1 _6517_ (.B1(_2132_),
    .Y(_2133_),
    .A1(net2167),
    .A2(_2129_));
 sg13g2_a22oi_1 _6518_ (.Y(_2134_),
    .B1(_2133_),
    .B2(net2051),
    .A2(_2126_),
    .A1(net1898));
 sg13g2_nand2_1 _6519_ (.Y(_2135_),
    .A(_1672_),
    .B(_2134_));
 sg13g2_a21oi_1 _6520_ (.A1(net2230),
    .A2(_2009_),
    .Y(_2136_),
    .B1(_1791_));
 sg13g2_o21ai_1 _6521_ (.B1(net1908),
    .Y(_2137_),
    .A1(net2203),
    .A2(net1885));
 sg13g2_nor2_1 _6522_ (.A(_2136_),
    .B(_2137_),
    .Y(_2138_));
 sg13g2_nor2_1 _6523_ (.A(net2215),
    .B(_1596_),
    .Y(_2139_));
 sg13g2_nor3_1 _6524_ (.A(net1891),
    .B(_1517_),
    .C(_2139_),
    .Y(_2140_));
 sg13g2_a21oi_1 _6525_ (.A1(_1500_),
    .A2(net1789),
    .Y(_2141_),
    .B1(_2089_));
 sg13g2_nor3_1 _6526_ (.A(_2138_),
    .B(_2140_),
    .C(_2141_),
    .Y(_2142_));
 sg13g2_o21ai_1 _6527_ (.B1(_2086_),
    .Y(_2143_),
    .A1(net2229),
    .A2(_1902_));
 sg13g2_a21oi_1 _6528_ (.A1(net2199),
    .A2(_2143_),
    .Y(_2144_),
    .B1(net2183));
 sg13g2_nand2_1 _6529_ (.Y(_2145_),
    .A(_1592_),
    .B(_1709_));
 sg13g2_a21oi_1 _6530_ (.A1(_2010_),
    .A2(_2145_),
    .Y(_2146_),
    .B1(_1481_));
 sg13g2_nor2_2 _6531_ (.A(net2186),
    .B(net1834),
    .Y(_2147_));
 sg13g2_nor2_2 _6532_ (.A(net1904),
    .B(net1834),
    .Y(_2148_));
 sg13g2_and2_1 _6533_ (.A(net1884),
    .B(_1724_),
    .X(_2149_));
 sg13g2_nand3_1 _6534_ (.B(net1947),
    .C(_1796_),
    .A(_1536_),
    .Y(_2150_));
 sg13g2_nor3_1 _6535_ (.A(net1945),
    .B(_2149_),
    .C(_2150_),
    .Y(_2151_));
 sg13g2_nor2_1 _6536_ (.A(net1932),
    .B(_2151_),
    .Y(_2152_));
 sg13g2_nor4_1 _6537_ (.A(net1938),
    .B(_2146_),
    .C(_2148_),
    .D(_2152_),
    .Y(_2153_));
 sg13g2_o21ai_1 _6538_ (.B1(_2153_),
    .Y(_2154_),
    .A1(net2167),
    .A2(_2144_));
 sg13g2_o21ai_1 _6539_ (.B1(_2154_),
    .Y(_2155_),
    .A1(net1893),
    .A2(_2142_));
 sg13g2_nor2_1 _6540_ (.A(net2242),
    .B(_1624_),
    .Y(_2156_));
 sg13g2_nand2b_1 _6541_ (.Y(_2157_),
    .B(net1790),
    .A_N(net2243));
 sg13g2_o21ai_1 _6542_ (.B1(_1626_),
    .Y(_2158_),
    .A1(net1866),
    .A2(_2157_));
 sg13g2_nand3_1 _6543_ (.B(_1516_),
    .C(_1764_),
    .A(net1877),
    .Y(_2159_));
 sg13g2_nand4_1 _6544_ (.B(net1951),
    .C(net1790),
    .A(net2243),
    .Y(_2160_),
    .D(_1732_));
 sg13g2_or4_1 _6545_ (.A(net2179),
    .B(net1877),
    .C(net1930),
    .D(_1731_),
    .X(_2161_));
 sg13g2_nand2_1 _6546_ (.Y(_2162_),
    .A(_2160_),
    .B(_2161_));
 sg13g2_a221oi_1 _6547_ (.B2(net1911),
    .C1(_2162_),
    .B1(_2159_),
    .A1(net1798),
    .Y(_2163_),
    .A2(_2158_));
 sg13g2_a21oi_1 _6548_ (.A1(_1575_),
    .A2(_2054_),
    .Y(_2164_),
    .B1(net1889));
 sg13g2_nand3_1 _6549_ (.B(_1660_),
    .C(_2054_),
    .A(net2210),
    .Y(_2165_));
 sg13g2_o21ai_1 _6550_ (.B1(net2191),
    .Y(_2166_),
    .A1(net2210),
    .A2(_1572_));
 sg13g2_nor2_1 _6551_ (.A(net2048),
    .B(_2166_),
    .Y(_2167_));
 sg13g2_a21oi_1 _6552_ (.A1(_2165_),
    .A2(_2167_),
    .Y(_2168_),
    .B1(_2164_));
 sg13g2_nand3_1 _6553_ (.B(_2163_),
    .C(_2168_),
    .A(net1730),
    .Y(_2169_));
 sg13g2_o21ai_1 _6554_ (.B1(_1645_),
    .Y(_2170_),
    .A1(net2033),
    .A2(_1513_));
 sg13g2_nand2_1 _6555_ (.Y(_2171_),
    .A(net1854),
    .B(_2170_));
 sg13g2_nor2_2 _6556_ (.A(net1886),
    .B(_1733_),
    .Y(_2172_));
 sg13g2_nor2_2 _6557_ (.A(net1976),
    .B(net1856),
    .Y(_2173_));
 sg13g2_a21oi_1 _6558_ (.A1(net2248),
    .A2(_1507_),
    .Y(_2174_),
    .B1(_2012_));
 sg13g2_o21ai_1 _6559_ (.B1(_2160_),
    .Y(_2175_),
    .A1(net1877),
    .A2(net1856));
 sg13g2_a221oi_1 _6560_ (.B2(_1623_),
    .C1(_2175_),
    .B1(_2174_),
    .A1(_1654_),
    .Y(_2176_),
    .A2(_2172_));
 sg13g2_a21oi_1 _6561_ (.A1(net1884),
    .A2(_2047_),
    .Y(_2177_),
    .B1(net1946));
 sg13g2_nor2_1 _6562_ (.A(net1889),
    .B(_2177_),
    .Y(_2178_));
 sg13g2_nand2_1 _6563_ (.Y(_2179_),
    .A(net1969),
    .B(net1806));
 sg13g2_nand3_1 _6564_ (.B(net1882),
    .C(_1749_),
    .A(net1909),
    .Y(_2180_));
 sg13g2_nand2_1 _6565_ (.Y(_2181_),
    .A(_1546_),
    .B(_2180_));
 sg13g2_a21oi_1 _6566_ (.A1(_2179_),
    .A2(_2181_),
    .Y(_2182_),
    .B1(_2178_));
 sg13g2_nand4_1 _6567_ (.B(_2171_),
    .C(_2176_),
    .A(net1743),
    .Y(_2183_),
    .D(_2182_));
 sg13g2_a21oi_2 _6568_ (.B1(net1938),
    .Y(_2184_),
    .A2(_2183_),
    .A1(_2169_));
 sg13g2_nor2_2 _6569_ (.A(_1673_),
    .B(_1931_),
    .Y(_2185_));
 sg13g2_nor2_1 _6570_ (.A(_1670_),
    .B(_2185_),
    .Y(_2186_));
 sg13g2_a21oi_1 _6571_ (.A1(net1800),
    .A2(_1670_),
    .Y(_2187_),
    .B1(_2186_));
 sg13g2_or2_1 _6572_ (.X(_2188_),
    .B(_2122_),
    .A(net2038));
 sg13g2_nand2_1 _6573_ (.Y(_2189_),
    .A(_1613_),
    .B(net1929));
 sg13g2_nand2_1 _6574_ (.Y(_2190_),
    .A(net2168),
    .B(_2189_));
 sg13g2_nand3_1 _6575_ (.B(_2188_),
    .C(_2189_),
    .A(net2168),
    .Y(_2191_));
 sg13g2_a21oi_2 _6576_ (.B1(_1530_),
    .Y(_2192_),
    .A2(net2140),
    .A1(net2216));
 sg13g2_o21ai_1 _6577_ (.B1(net2155),
    .Y(_2193_),
    .A1(_3995_),
    .A2(_2192_));
 sg13g2_o21ai_1 _6578_ (.B1(_2191_),
    .Y(_2194_),
    .A1(net2168),
    .A2(_2187_));
 sg13g2_nor2_2 _6579_ (.A(net1869),
    .B(net1930),
    .Y(_2195_));
 sg13g2_nor2_1 _6580_ (.A(net1929),
    .B(_1960_),
    .Y(_2196_));
 sg13g2_a221oi_1 _6581_ (.B2(net2201),
    .C1(net1888),
    .B1(_2185_),
    .A1(net1957),
    .Y(_2197_),
    .A2(net1871));
 sg13g2_o21ai_1 _6582_ (.B1(net1942),
    .Y(_2198_),
    .A1(net1857),
    .A2(_1613_));
 sg13g2_nor2_1 _6583_ (.A(_2197_),
    .B(_2198_),
    .Y(_2199_));
 sg13g2_o21ai_1 _6584_ (.B1(_2199_),
    .Y(_2200_),
    .A1(_2190_),
    .A2(_2196_));
 sg13g2_o21ai_1 _6585_ (.B1(_2200_),
    .Y(_2201_),
    .A1(_2193_),
    .A2(_2194_));
 sg13g2_nor2b_1 _6586_ (.A(_1951_),
    .B_N(_2201_),
    .Y(_2202_));
 sg13g2_nor4_2 _6587_ (.A(net2134),
    .B(net1876),
    .C(net1966),
    .Y(_2203_),
    .D(_1724_));
 sg13g2_nor3_2 _6588_ (.A(net1932),
    .B(_1802_),
    .C(_2203_),
    .Y(_2204_));
 sg13g2_nor2_2 _6589_ (.A(net1987),
    .B(net1841),
    .Y(_2205_));
 sg13g2_a21oi_2 _6590_ (.B1(_2205_),
    .Y(_2206_),
    .A2(net1836),
    .A1(net1960));
 sg13g2_a22oi_1 _6591_ (.Y(_2207_),
    .B1(_2052_),
    .B2(net2195),
    .A2(_1955_),
    .A1(_1624_));
 sg13g2_a21oi_1 _6592_ (.A1(net2049),
    .A2(_2207_),
    .Y(_2208_),
    .B1(_2204_));
 sg13g2_a221oi_1 _6593_ (.B2(net1910),
    .C1(net1940),
    .B1(_2206_),
    .A1(net1798),
    .Y(_2209_),
    .A2(_2050_));
 sg13g2_nand3_1 _6594_ (.B(_1942_),
    .C(_2157_),
    .A(_1926_),
    .Y(_2210_));
 sg13g2_a21oi_1 _6595_ (.A1(net2232),
    .A2(net1975),
    .Y(_2211_),
    .B1(net2030));
 sg13g2_a221oi_1 _6596_ (.B2(net2243),
    .C1(net2035),
    .B1(_1701_),
    .A1(net2132),
    .Y(_2212_),
    .A2(net1971));
 sg13g2_o21ai_1 _6597_ (.B1(net1860),
    .Y(_2213_),
    .A1(_2058_),
    .A2(_2212_));
 sg13g2_o21ai_1 _6598_ (.B1(net2214),
    .Y(_2214_),
    .A1(_1625_),
    .A2(_1651_));
 sg13g2_a21oi_1 _6599_ (.A1(_2048_),
    .A2(_2214_),
    .Y(_2215_),
    .B1(net1935));
 sg13g2_a21oi_1 _6600_ (.A1(net2035),
    .A2(_1701_),
    .Y(_2216_),
    .B1(_1872_));
 sg13g2_nor3_1 _6601_ (.A(net2219),
    .B(net2149),
    .C(net2137),
    .Y(_2217_));
 sg13g2_nor3_1 _6602_ (.A(net1889),
    .B(net1972),
    .C(_2217_),
    .Y(_2218_));
 sg13g2_nor4_1 _6603_ (.A(net1896),
    .B(_2215_),
    .C(_2216_),
    .D(_2218_),
    .Y(_2219_));
 sg13g2_a22oi_1 _6604_ (.Y(_2220_),
    .B1(_2213_),
    .B2(_2219_),
    .A2(_2209_),
    .A1(_2208_));
 sg13g2_a21oi_2 _6605_ (.B1(_1899_),
    .Y(_2221_),
    .A2(_2220_),
    .A1(_2210_));
 sg13g2_nor2_1 _6606_ (.A(_2202_),
    .B(_2221_),
    .Y(_2222_));
 sg13g2_a22oi_1 _6607_ (.Y(_2223_),
    .B1(_2155_),
    .B2(_1747_),
    .A2(_2118_),
    .A1(net1731));
 sg13g2_nand4_1 _6608_ (.B(_2135_),
    .C(_2222_),
    .A(\draw_game_inst.board_x[0] ),
    .Y(_2224_),
    .D(_2223_));
 sg13g2_nor4_1 _6609_ (.A(_2077_),
    .B(_2099_),
    .C(_2184_),
    .D(_2224_),
    .Y(_2225_));
 sg13g2_nand2b_1 _6610_ (.Y(_2226_),
    .B(net998),
    .A_N(net995));
 sg13g2_a21oi_1 _6611_ (.A1(_2043_),
    .A2(_2225_),
    .Y(_2227_),
    .B1(_1983_));
 sg13g2_a221oi_1 _6612_ (.B2(net2134),
    .C1(net2189),
    .B1(net1848),
    .A1(net2204),
    .Y(_2228_),
    .A2(net1974));
 sg13g2_a221oi_1 _6613_ (.B2(net1882),
    .C1(net2171),
    .B1(_1715_),
    .A1(net1996),
    .Y(_2229_),
    .A2(net1955));
 sg13g2_nor2_1 _6614_ (.A(net1981),
    .B(net1973),
    .Y(_2230_));
 sg13g2_a22oi_1 _6615_ (.Y(_2231_),
    .B1(_2230_),
    .B2(_1799_),
    .A2(_1850_),
    .A1(net1955));
 sg13g2_nand3_1 _6616_ (.B(_2024_),
    .C(_2231_),
    .A(_1867_),
    .Y(_2232_));
 sg13g2_o21ai_1 _6617_ (.B1(net2203),
    .Y(_2233_),
    .A1(net1885),
    .A2(net1877));
 sg13g2_a22oi_1 _6618_ (.Y(_2234_),
    .B1(_2233_),
    .B2(_1807_),
    .A2(_2229_),
    .A1(_2228_));
 sg13g2_nand2_1 _6619_ (.Y(_2235_),
    .A(_2232_),
    .B(_2234_));
 sg13g2_nor2_2 _6620_ (.A(net1928),
    .B(_1977_),
    .Y(_2236_));
 sg13g2_a21oi_1 _6621_ (.A1(net2200),
    .A2(net1871),
    .Y(_2237_),
    .B1(net2186));
 sg13g2_o21ai_1 _6622_ (.B1(_1908_),
    .Y(_2238_),
    .A1(net2229),
    .A2(_1902_));
 sg13g2_o21ai_1 _6623_ (.B1(_2237_),
    .Y(_2239_),
    .A1(net2200),
    .A2(_2238_));
 sg13g2_nor2_1 _6624_ (.A(net1872),
    .B(net1930),
    .Y(_2240_));
 sg13g2_nand2_1 _6625_ (.Y(_2241_),
    .A(net1850),
    .B(_1673_));
 sg13g2_nand3_1 _6626_ (.B(_2239_),
    .C(_2241_),
    .A(_1831_),
    .Y(_2242_));
 sg13g2_o21ai_1 _6627_ (.B1(net1794),
    .Y(_2243_),
    .A1(net2199),
    .A2(_1652_));
 sg13g2_o21ai_1 _6628_ (.B1(_2242_),
    .Y(_2244_),
    .A1(_1836_),
    .A2(_2243_));
 sg13g2_a22oi_1 _6629_ (.Y(_2245_),
    .B1(_2244_),
    .B2(net1742),
    .A2(_2235_),
    .A1(net1729));
 sg13g2_or2_1 _6630_ (.X(_2246_),
    .B(_1572_),
    .A(net1887));
 sg13g2_nor2_2 _6631_ (.A(_1570_),
    .B(_1764_),
    .Y(_2247_));
 sg13g2_a21oi_1 _6632_ (.A1(net1878),
    .A2(_1721_),
    .Y(_2248_),
    .B1(_1630_));
 sg13g2_nand2b_1 _6633_ (.Y(_2249_),
    .B(_2248_),
    .A_N(_2247_));
 sg13g2_a21oi_1 _6634_ (.A1(net1877),
    .A2(_1630_),
    .Y(_2250_),
    .B1(net2164));
 sg13g2_a22oi_1 _6635_ (.Y(_2251_),
    .B1(_2249_),
    .B2(_2250_),
    .A2(_2246_),
    .A1(net2163));
 sg13g2_nand2_1 _6636_ (.Y(_2252_),
    .A(_1516_),
    .B(_1524_));
 sg13g2_nand2_1 _6637_ (.Y(_2253_),
    .A(_2034_),
    .B(_2252_));
 sg13g2_nand2_1 _6638_ (.Y(_2254_),
    .A(_1574_),
    .B(net1835));
 sg13g2_a21oi_1 _6639_ (.A1(net2191),
    .A2(_2254_),
    .Y(_2255_),
    .B1(net2174));
 sg13g2_o21ai_1 _6640_ (.B1(_1562_),
    .Y(_2256_),
    .A1(net2226),
    .A2(_1685_));
 sg13g2_nand2_1 _6641_ (.Y(_2257_),
    .A(net1853),
    .B(_2256_));
 sg13g2_a221oi_1 _6642_ (.B2(_2255_),
    .C1(net2163),
    .B1(_2253_),
    .A1(net1834),
    .Y(_2258_),
    .A2(net1794));
 sg13g2_a22oi_1 _6643_ (.Y(_2259_),
    .B1(_2257_),
    .B2(_2258_),
    .A2(_1501_),
    .A1(net2163));
 sg13g2_a22oi_1 _6644_ (.Y(_2260_),
    .B1(_2259_),
    .B2(net1743),
    .A2(_2251_),
    .A1(_1602_));
 sg13g2_o21ai_1 _6645_ (.B1(_2260_),
    .Y(_2261_),
    .A1(net2165),
    .A2(_2245_));
 sg13g2_nand2_1 _6646_ (.Y(_2262_),
    .A(net2155),
    .B(_2261_));
 sg13g2_a21oi_1 _6647_ (.A1(net2213),
    .A2(net1810),
    .Y(_2263_),
    .B1(net2192));
 sg13g2_nand2_1 _6648_ (.Y(_2264_),
    .A(net2037),
    .B(_1923_));
 sg13g2_nand3_1 _6649_ (.B(_1693_),
    .C(_2264_),
    .A(net2192),
    .Y(_2265_));
 sg13g2_a21oi_1 _6650_ (.A1(_2177_),
    .A2(_2263_),
    .Y(_2266_),
    .B1(net2176));
 sg13g2_nand2_1 _6651_ (.Y(_2267_),
    .A(_2265_),
    .B(_2266_));
 sg13g2_o21ai_1 _6652_ (.B1(_1784_),
    .Y(_2268_),
    .A1(net2037),
    .A2(_1513_));
 sg13g2_nand3_1 _6653_ (.B(_2068_),
    .C(_2268_),
    .A(net2176),
    .Y(_2269_));
 sg13g2_nand4_1 _6654_ (.B(net1944),
    .C(_2267_),
    .A(net1743),
    .Y(_2270_),
    .D(_2269_));
 sg13g2_a21oi_2 _6655_ (.B1(_1737_),
    .Y(_2271_),
    .A2(net1884),
    .A1(net2136));
 sg13g2_o21ai_1 _6656_ (.B1(net1843),
    .Y(_2272_),
    .A1(net2024),
    .A2(net1886));
 sg13g2_nand2b_2 _6657_ (.Y(_2273_),
    .B(_2272_),
    .A_N(net2247));
 sg13g2_nor2_1 _6658_ (.A(net2216),
    .B(_1763_),
    .Y(_2274_));
 sg13g2_nand2_2 _6659_ (.Y(_2275_),
    .A(_1530_),
    .B(_1558_));
 sg13g2_and2_1 _6660_ (.A(net2216),
    .B(_1912_),
    .X(_2276_));
 sg13g2_a221oi_1 _6661_ (.B2(_2276_),
    .C1(net1905),
    .B1(_2275_),
    .A1(_2273_),
    .Y(_2277_),
    .A2(_2274_));
 sg13g2_nor2_1 _6662_ (.A(net1989),
    .B(_2272_),
    .Y(_2278_));
 sg13g2_o21ai_1 _6663_ (.B1(net1860),
    .Y(_2279_),
    .A1(net1983),
    .A2(net1884));
 sg13g2_nand2_2 _6664_ (.Y(_2280_),
    .A(net1881),
    .B(_1795_));
 sg13g2_nand3_1 _6665_ (.B(_1725_),
    .C(_2280_),
    .A(net1994),
    .Y(_2281_));
 sg13g2_o21ai_1 _6666_ (.B1(_2281_),
    .Y(_2282_),
    .A1(_2278_),
    .A2(_2279_));
 sg13g2_nor4_1 _6667_ (.A(_1736_),
    .B(_2172_),
    .C(_2277_),
    .D(_2282_),
    .Y(_2283_));
 sg13g2_a21oi_1 _6668_ (.A1(net1973),
    .A2(net1967),
    .Y(_2284_),
    .B1(net2140));
 sg13g2_nor2_1 _6669_ (.A(net2197),
    .B(_2284_),
    .Y(_2285_));
 sg13g2_o21ai_1 _6670_ (.B1(net2197),
    .Y(_2286_),
    .A1(net1883),
    .A2(net1963));
 sg13g2_o21ai_1 _6671_ (.B1(net2181),
    .Y(_2287_),
    .A1(_1555_),
    .A2(_2286_));
 sg13g2_nor2_1 _6672_ (.A(_2285_),
    .B(_2287_),
    .Y(_2288_));
 sg13g2_a21oi_1 _6673_ (.A1(net2049),
    .A2(_1718_),
    .Y(_2289_),
    .B1(_2288_));
 sg13g2_nand2b_2 _6674_ (.Y(_2290_),
    .B(_2001_),
    .A_N(net2247));
 sg13g2_nand2b_1 _6675_ (.Y(_2291_),
    .B(_2290_),
    .A_N(_1610_));
 sg13g2_a21oi_1 _6676_ (.A1(_2275_),
    .A2(_2290_),
    .Y(_2292_),
    .B1(_1481_));
 sg13g2_nor3_1 _6677_ (.A(net1941),
    .B(_2289_),
    .C(_2292_),
    .Y(_2293_));
 sg13g2_o21ai_1 _6678_ (.B1(_1698_),
    .Y(_2294_),
    .A1(_2283_),
    .A2(_2293_));
 sg13g2_a21oi_1 _6679_ (.A1(_1583_),
    .A2(_1748_),
    .Y(_2295_),
    .B1(_2032_));
 sg13g2_nor3_1 _6680_ (.A(net1981),
    .B(net1812),
    .C(net1973),
    .Y(_2296_));
 sg13g2_a221oi_1 _6681_ (.B2(_2295_),
    .C1(net1897),
    .B1(net1858),
    .A1(net1992),
    .Y(_2297_),
    .A2(_1517_));
 sg13g2_o21ai_1 _6682_ (.B1(_2297_),
    .Y(_2298_),
    .A1(net1933),
    .A2(_2296_));
 sg13g2_a221oi_1 _6683_ (.B2(net1908),
    .C1(_2298_),
    .B1(_2136_),
    .A1(net1927),
    .Y(_2299_),
    .A2(net1841));
 sg13g2_o21ai_1 _6684_ (.B1(net2203),
    .Y(_2300_),
    .A1(net2135),
    .A2(net1809));
 sg13g2_nand2_1 _6685_ (.Y(_2301_),
    .A(_1760_),
    .B(_2300_));
 sg13g2_nor2_1 _6686_ (.A(net1877),
    .B(_1753_),
    .Y(_2302_));
 sg13g2_nor2_1 _6687_ (.A(net1981),
    .B(_2302_),
    .Y(_2303_));
 sg13g2_o21ai_1 _6688_ (.B1(net1908),
    .Y(_2304_),
    .A1(_2053_),
    .A2(_2303_));
 sg13g2_o21ai_1 _6689_ (.B1(_1752_),
    .Y(_2305_),
    .A1(_2205_),
    .A2(_2304_));
 sg13g2_a21oi_1 _6690_ (.A1(net1839),
    .A2(_2301_),
    .Y(_2306_),
    .B1(_2305_));
 sg13g2_o21ai_1 _6691_ (.B1(_1747_),
    .Y(_2307_),
    .A1(_2299_),
    .A2(_2306_));
 sg13g2_nor3_2 _6692_ (.A(net1880),
    .B(net1963),
    .C(_1570_),
    .Y(_2308_));
 sg13g2_a221oi_1 _6693_ (.B2(net1993),
    .C1(_2164_),
    .B1(_2308_),
    .A1(_1647_),
    .Y(_2309_),
    .A2(_1836_));
 sg13g2_a22oi_1 _6694_ (.Y(_2310_),
    .B1(net1790),
    .B2(_2173_),
    .A2(net1859),
    .A1(net1988));
 sg13g2_a21oi_1 _6695_ (.A1(net1988),
    .A2(_1851_),
    .Y(_2311_),
    .B1(_2310_));
 sg13g2_nand2_1 _6696_ (.Y(_2312_),
    .A(net2218),
    .B(net1800));
 sg13g2_o21ai_1 _6697_ (.B1(_2312_),
    .Y(_2313_),
    .A1(net1877),
    .A2(_1731_));
 sg13g2_nor2_1 _6698_ (.A(net1938),
    .B(_1638_),
    .Y(_2314_));
 sg13g2_a21oi_1 _6699_ (.A1(net1909),
    .A2(_2313_),
    .Y(_2315_),
    .B1(_2311_));
 sg13g2_nand4_1 _6700_ (.B(_2309_),
    .C(_2314_),
    .A(net1730),
    .Y(_2316_),
    .D(_2315_));
 sg13g2_nand4_1 _6701_ (.B(_2294_),
    .C(_2307_),
    .A(_2270_),
    .Y(_2317_),
    .D(_2316_));
 sg13g2_a21o_1 _6702_ (.A2(_2188_),
    .A1(_1976_),
    .B1(_2121_),
    .X(_2318_));
 sg13g2_a21oi_1 _6703_ (.A1(net1907),
    .A2(_2192_),
    .Y(_2319_),
    .B1(_1677_));
 sg13g2_o21ai_1 _6704_ (.B1(_1672_),
    .Y(_2320_),
    .A1(net2155),
    .A2(_2319_));
 sg13g2_a21oi_1 _6705_ (.A1(net1898),
    .A2(_2318_),
    .Y(_2321_),
    .B1(_2320_));
 sg13g2_a221oi_1 _6706_ (.B2(_1700_),
    .C1(net1929),
    .B1(_1931_),
    .A1(net1950),
    .Y(_2322_),
    .A2(_1763_));
 sg13g2_a21oi_2 _6707_ (.B1(net2187),
    .Y(_2323_),
    .A2(net1834),
    .A1(net1987));
 sg13g2_a221oi_1 _6708_ (.B2(_2323_),
    .C1(_2322_),
    .B1(_2079_),
    .A1(net1846),
    .Y(_2324_),
    .A2(_1902_));
 sg13g2_nor2_1 _6709_ (.A(net1839),
    .B(_2324_),
    .Y(_2325_));
 sg13g2_a21oi_1 _6710_ (.A1(net2229),
    .A2(_1837_),
    .Y(_2326_),
    .B1(_1688_));
 sg13g2_a22oi_1 _6711_ (.Y(_2327_),
    .B1(net1841),
    .B2(_1649_),
    .A2(_1684_),
    .A1(net1982));
 sg13g2_nor2_1 _6712_ (.A(_2326_),
    .B(_2327_),
    .Y(_2328_));
 sg13g2_a21oi_1 _6713_ (.A1(net2039),
    .A2(net1885),
    .Y(_2329_),
    .B1(net1868));
 sg13g2_a221oi_1 _6714_ (.B2(net2045),
    .C1(_1888_),
    .B1(_2329_),
    .A1(net1907),
    .Y(_2330_),
    .A2(_2328_));
 sg13g2_nor2b_1 _6715_ (.A(_1717_),
    .B_N(_1644_),
    .Y(_2331_));
 sg13g2_nor4_1 _6716_ (.A(net2171),
    .B(_1751_),
    .C(_1759_),
    .D(_2331_),
    .Y(_2332_));
 sg13g2_nor3_1 _6717_ (.A(_2325_),
    .B(_2330_),
    .C(_2332_),
    .Y(_2333_));
 sg13g2_nor2_1 _6718_ (.A(_1857_),
    .B(_2333_),
    .Y(_2334_));
 sg13g2_nor4_1 _6719_ (.A(net1731),
    .B(_2317_),
    .C(_2321_),
    .D(_2334_),
    .Y(_2335_));
 sg13g2_a21oi_1 _6720_ (.A1(net2144),
    .A2(net2145),
    .Y(_2336_),
    .B1(_1557_));
 sg13g2_a21oi_1 _6721_ (.A1(net1960),
    .A2(_1867_),
    .Y(_2337_),
    .B1(_2336_));
 sg13g2_o21ai_1 _6722_ (.B1(net2039),
    .Y(_2338_),
    .A1(_1645_),
    .A2(_1802_));
 sg13g2_nor2_1 _6723_ (.A(_2337_),
    .B(_2338_),
    .Y(_2339_));
 sg13g2_nand3_1 _6724_ (.B(_1700_),
    .C(net1842),
    .A(net2029),
    .Y(_2340_));
 sg13g2_nand2b_2 _6725_ (.Y(_2341_),
    .B(_1739_),
    .A_N(net2232));
 sg13g2_nand3_1 _6726_ (.B(_2275_),
    .C(_2341_),
    .A(net1850),
    .Y(_2342_));
 sg13g2_o21ai_1 _6727_ (.B1(_2342_),
    .Y(_2343_),
    .A1(net1844),
    .A2(net1797));
 sg13g2_o21ai_1 _6728_ (.B1(net1729),
    .Y(_2344_),
    .A1(_2339_),
    .A2(_2343_));
 sg13g2_a21oi_1 _6729_ (.A1(_1537_),
    .A2(_1650_),
    .Y(_2345_),
    .B1(_1497_));
 sg13g2_a21o_1 _6730_ (.A2(net1874),
    .A1(net2240),
    .B1(_2345_),
    .X(_2346_));
 sg13g2_nand2b_2 _6731_ (.Y(_2347_),
    .B(_1660_),
    .A_N(_1654_));
 sg13g2_nand2_1 _6732_ (.Y(_2348_),
    .A(_1908_),
    .B(_2093_));
 sg13g2_nand3_1 _6733_ (.B(net1803),
    .C(_2348_),
    .A(net2187),
    .Y(_2349_));
 sg13g2_a22oi_1 _6734_ (.Y(_2350_),
    .B1(_2347_),
    .B2(net1927),
    .A2(_2346_),
    .A1(net1912));
 sg13g2_nand3_1 _6735_ (.B(_2349_),
    .C(_2350_),
    .A(_1822_),
    .Y(_2351_));
 sg13g2_a21oi_1 _6736_ (.A1(_2344_),
    .A2(_2351_),
    .Y(_2352_),
    .B1(_1811_));
 sg13g2_o21ai_1 _6737_ (.B1(net2176),
    .Y(_2353_),
    .A1(net2192),
    .A2(_1858_));
 sg13g2_a21oi_1 _6738_ (.A1(net1878),
    .A2(_1763_),
    .Y(_2354_),
    .B1(_1604_));
 sg13g2_nor2_2 _6739_ (.A(net1801),
    .B(net1930),
    .Y(_2355_));
 sg13g2_a21oi_1 _6740_ (.A1(net1878),
    .A2(_2355_),
    .Y(_2356_),
    .B1(_2353_));
 sg13g2_o21ai_1 _6741_ (.B1(_2356_),
    .Y(_2357_),
    .A1(_1641_),
    .A2(_2354_));
 sg13g2_nand2_1 _6742_ (.Y(_2358_),
    .A(_1519_),
    .B(net1788));
 sg13g2_a221oi_1 _6743_ (.B2(_1616_),
    .C1(net2176),
    .B1(_2358_),
    .A1(_1595_),
    .Y(_2359_),
    .A2(net1845));
 sg13g2_o21ai_1 _6744_ (.B1(_2359_),
    .Y(_2360_),
    .A1(net2192),
    .A2(_1919_));
 sg13g2_a21oi_1 _6745_ (.A1(_2357_),
    .A2(_2360_),
    .Y(_2361_),
    .B1(net1939));
 sg13g2_nor2_2 _6746_ (.A(net2188),
    .B(_1517_),
    .Y(_2362_));
 sg13g2_o21ai_1 _6747_ (.B1(_2362_),
    .Y(_2363_),
    .A1(net2214),
    .A2(_1701_));
 sg13g2_nand2b_1 _6748_ (.Y(_2364_),
    .B(_1784_),
    .A_N(_1916_));
 sg13g2_nand3_1 _6749_ (.B(_2363_),
    .C(_2364_),
    .A(net2181),
    .Y(_2365_));
 sg13g2_nor3_2 _6750_ (.A(net2143),
    .B(_1515_),
    .C(_1651_),
    .Y(_2366_));
 sg13g2_nor2b_1 _6751_ (.A(_2366_),
    .B_N(_2173_),
    .Y(_2367_));
 sg13g2_nand2_1 _6752_ (.Y(_2368_),
    .A(net1883),
    .B(net1967));
 sg13g2_a22oi_1 _6753_ (.Y(_2369_),
    .B1(_1558_),
    .B2(net2215),
    .A2(net1804),
    .A1(net1963));
 sg13g2_o21ai_1 _6754_ (.B1(_2365_),
    .Y(_2370_),
    .A1(net1890),
    .A2(_2369_));
 sg13g2_nor3_1 _6755_ (.A(net1896),
    .B(_2367_),
    .C(_2370_),
    .Y(_2371_));
 sg13g2_nor3_1 _6756_ (.A(net1810),
    .B(_1534_),
    .C(_1927_),
    .Y(_2372_));
 sg13g2_nor3_1 _6757_ (.A(_2361_),
    .B(_2371_),
    .C(_2372_),
    .Y(_2373_));
 sg13g2_nor2_1 _6758_ (.A(_1899_),
    .B(_2373_),
    .Y(_2374_));
 sg13g2_o21ai_1 _6759_ (.B1(_1953_),
    .Y(_2375_),
    .A1(net1948),
    .A2(_1860_));
 sg13g2_nand2_1 _6760_ (.Y(_2376_),
    .A(net1846),
    .B(_2347_));
 sg13g2_a21oi_1 _6761_ (.A1(net1850),
    .A2(_1960_),
    .Y(_2377_),
    .B1(_1962_));
 sg13g2_nand2_2 _6762_ (.Y(_2378_),
    .A(net2189),
    .B(_1509_));
 sg13g2_a221oi_1 _6763_ (.B2(_1682_),
    .C1(net1894),
    .B1(_2378_),
    .A1(_2376_),
    .Y(_2379_),
    .A2(_2377_));
 sg13g2_a21oi_1 _6764_ (.A1(_1574_),
    .A2(_1674_),
    .Y(_2380_),
    .B1(net1888));
 sg13g2_nor3_1 _6765_ (.A(net2161),
    .B(_2018_),
    .C(_2380_),
    .Y(_2381_));
 sg13g2_o21ai_1 _6766_ (.B1(_1574_),
    .Y(_2382_),
    .A1(_1543_),
    .A2(net1865));
 sg13g2_o21ai_1 _6767_ (.B1(net2168),
    .Y(_2383_),
    .A1(net2183),
    .A2(_2382_));
 sg13g2_a21oi_1 _6768_ (.A1(_2381_),
    .A2(_2383_),
    .Y(_2384_),
    .B1(net2156));
 sg13g2_nor3_1 _6769_ (.A(_2375_),
    .B(_2379_),
    .C(_2384_),
    .Y(_2385_));
 sg13g2_nor3_1 _6770_ (.A(_2352_),
    .B(_2374_),
    .C(_2385_),
    .Y(_2386_));
 sg13g2_nand3_1 _6771_ (.B(_2335_),
    .C(_2386_),
    .A(_2262_),
    .Y(_2387_));
 sg13g2_nor4_1 _6772_ (.A(net2225),
    .B(net2198),
    .C(net2183),
    .D(net1862),
    .Y(_2388_));
 sg13g2_nand2b_1 _6773_ (.Y(_2389_),
    .B(net2167),
    .A_N(_2388_));
 sg13g2_a21oi_1 _6774_ (.A1(_2381_),
    .A2(_2389_),
    .Y(_2390_),
    .B1(net2156));
 sg13g2_nor2_1 _6775_ (.A(net2225),
    .B(net2198),
    .Y(_2391_));
 sg13g2_nand2_1 _6776_ (.Y(_2392_),
    .A(_2103_),
    .B(_2391_));
 sg13g2_a21oi_1 _6777_ (.A1(net1991),
    .A2(net1861),
    .Y(_2393_),
    .B1(_1978_));
 sg13g2_and3_2 _6778_ (.X(_2394_),
    .A(net2225),
    .B(net2198),
    .C(net1865));
 sg13g2_nor2_1 _6779_ (.A(_1543_),
    .B(_2394_),
    .Y(_2395_));
 sg13g2_a22oi_1 _6780_ (.Y(_2396_),
    .B1(_2395_),
    .B2(net1858),
    .A2(_2392_),
    .A1(net1851));
 sg13g2_a21oi_1 _6781_ (.A1(_2393_),
    .A2(_2396_),
    .Y(_2397_),
    .B1(net1893));
 sg13g2_or3_1 _6782_ (.A(_2111_),
    .B(_2390_),
    .C(_2397_),
    .X(_2398_));
 sg13g2_a21oi_1 _6783_ (.A1(net1731),
    .A2(_2398_),
    .Y(_2399_),
    .B1(_2226_));
 sg13g2_a22oi_1 _6784_ (.Y(_2400_),
    .B1(_2387_),
    .B2(_2399_),
    .A2(_2227_),
    .A1(_2226_));
 sg13g2_nand2_1 _6785_ (.Y(_2401_),
    .A(net2174),
    .B(_2048_));
 sg13g2_a21oi_1 _6786_ (.A1(net2211),
    .A2(_2347_),
    .Y(_2402_),
    .B1(_2401_));
 sg13g2_nand2_1 _6787_ (.Y(_2403_),
    .A(_1613_),
    .B(_1650_));
 sg13g2_a221oi_1 _6788_ (.B2(_2403_),
    .C1(_2186_),
    .B1(net1912),
    .A1(net2174),
    .Y(_2404_),
    .A2(net2043));
 sg13g2_a21oi_1 _6789_ (.A1(net2239),
    .A2(net1872),
    .Y(_2405_),
    .B1(_1630_));
 sg13g2_nor2_1 _6790_ (.A(_1516_),
    .B(net1856),
    .Y(_2406_));
 sg13g2_a221oi_1 _6791_ (.B2(_2405_),
    .C1(_2406_),
    .B1(_1988_),
    .A1(net1799),
    .Y(_2407_),
    .A2(net1845));
 sg13g2_o21ai_1 _6792_ (.B1(_2407_),
    .Y(_2408_),
    .A1(_2402_),
    .A2(_2404_));
 sg13g2_a221oi_1 _6793_ (.B2(net2238),
    .C1(_1643_),
    .B1(net1874),
    .A1(net2023),
    .Y(_2409_),
    .A2(net1976));
 sg13g2_a21oi_1 _6794_ (.A1(net1909),
    .A2(net1799),
    .Y(_2410_),
    .B1(_2409_));
 sg13g2_nand2_1 _6795_ (.Y(_2411_),
    .A(_1647_),
    .B(_1988_));
 sg13g2_a22oi_1 _6796_ (.Y(_2412_),
    .B1(_1629_),
    .B2(_1960_),
    .A2(_1623_),
    .A1(net1799));
 sg13g2_nand4_1 _6797_ (.B(_2410_),
    .C(_2411_),
    .A(_2114_),
    .Y(_2413_),
    .D(_2412_));
 sg13g2_a221oi_1 _6798_ (.B2(net2051),
    .C1(_2375_),
    .B1(_2413_),
    .A1(net1900),
    .Y(_2414_),
    .A2(_2408_));
 sg13g2_a21oi_1 _6799_ (.A1(net2230),
    .A2(net1806),
    .Y(_2415_),
    .B1(net2206));
 sg13g2_nor2_2 _6800_ (.A(net1804),
    .B(_1782_),
    .Y(_2416_));
 sg13g2_and2_1 _6801_ (.A(_1761_),
    .B(_2362_),
    .X(_2417_));
 sg13g2_nand2b_1 _6802_ (.Y(_2418_),
    .B(_2415_),
    .A_N(_1761_));
 sg13g2_a21oi_1 _6803_ (.A1(_2362_),
    .A2(_2418_),
    .Y(_2419_),
    .B1(_2416_));
 sg13g2_nor4_1 _6804_ (.A(net1902),
    .B(net1945),
    .C(_2136_),
    .D(_2149_),
    .Y(_2420_));
 sg13g2_nand2b_1 _6805_ (.Y(_2421_),
    .B(_2009_),
    .A_N(_2089_));
 sg13g2_o21ai_1 _6806_ (.B1(_2421_),
    .Y(_2422_),
    .A1(net2171),
    .A2(_2419_));
 sg13g2_o21ai_1 _6807_ (.B1(net1899),
    .Y(_2423_),
    .A1(_2420_),
    .A2(_2422_));
 sg13g2_a221oi_1 _6808_ (.B2(net2230),
    .C1(net2203),
    .B1(_1837_),
    .A1(_1592_),
    .Y(_2424_),
    .A2(_1709_));
 sg13g2_a21oi_1 _6809_ (.A1(net2203),
    .A2(_2302_),
    .Y(_2425_),
    .B1(_2424_));
 sg13g2_o21ai_1 _6810_ (.B1(net2047),
    .Y(_2426_),
    .A1(net2184),
    .A2(_2425_));
 sg13g2_nor3_1 _6811_ (.A(net1892),
    .B(net1945),
    .C(_1683_),
    .Y(_2427_));
 sg13g2_nor2_1 _6812_ (.A(net1932),
    .B(_2427_),
    .Y(_2428_));
 sg13g2_nand3_1 _6813_ (.B(_2304_),
    .C(_2426_),
    .A(net1942),
    .Y(_2429_));
 sg13g2_o21ai_1 _6814_ (.B1(_2423_),
    .Y(_2430_),
    .A1(_2428_),
    .A2(_2429_));
 sg13g2_nor2_1 _6815_ (.A(_1850_),
    .B(_2026_),
    .Y(_2431_));
 sg13g2_a21oi_1 _6816_ (.A1(net2227),
    .A2(net1787),
    .Y(_2432_),
    .B1(net2201));
 sg13g2_a21oi_1 _6817_ (.A1(_1932_),
    .A2(_2432_),
    .Y(_2433_),
    .B1(_2236_));
 sg13g2_o21ai_1 _6818_ (.B1(net1796),
    .Y(_2434_),
    .A1(net2236),
    .A2(net1837));
 sg13g2_a22oi_1 _6819_ (.Y(_2435_),
    .B1(_1864_),
    .B2(net1987),
    .A2(_1851_),
    .A1(net1957));
 sg13g2_a21oi_1 _6820_ (.A1(_2434_),
    .A2(_2435_),
    .Y(_2436_),
    .B1(net2040));
 sg13g2_nor3_1 _6821_ (.A(net2170),
    .B(_2433_),
    .C(_2436_),
    .Y(_2437_));
 sg13g2_o21ai_1 _6822_ (.B1(net1901),
    .Y(_2438_),
    .A1(_2431_),
    .A2(_2437_));
 sg13g2_nand2_1 _6823_ (.Y(_2439_),
    .A(net2210),
    .B(_1748_));
 sg13g2_nand2_1 _6824_ (.Y(_2440_),
    .A(net1964),
    .B(_2439_));
 sg13g2_a21oi_1 _6825_ (.A1(_1942_),
    .A2(_2440_),
    .Y(_2441_),
    .B1(_1992_));
 sg13g2_nor3_1 _6826_ (.A(net1867),
    .B(_1645_),
    .C(_1709_),
    .Y(_2442_));
 sg13g2_nand2_1 _6827_ (.Y(_2443_),
    .A(net1844),
    .B(_1692_));
 sg13g2_o21ai_1 _6828_ (.B1(_2443_),
    .Y(_2444_),
    .A1(_1861_),
    .A2(_2013_));
 sg13g2_o21ai_1 _6829_ (.B1(_1810_),
    .Y(_2445_),
    .A1(_2442_),
    .A2(_2444_));
 sg13g2_o21ai_1 _6830_ (.B1(_2438_),
    .Y(_2446_),
    .A1(_2441_),
    .A2(_2445_));
 sg13g2_and2_1 _6831_ (.A(net1729),
    .B(_2446_),
    .X(_2447_));
 sg13g2_a21oi_1 _6832_ (.A1(net1991),
    .A2(net1861),
    .Y(_2448_),
    .B1(_2121_));
 sg13g2_o21ai_1 _6833_ (.B1(_2448_),
    .Y(_2449_),
    .A1(net1857),
    .A2(_2123_));
 sg13g2_a21oi_1 _6834_ (.A1(net1982),
    .A2(net1871),
    .Y(_2450_),
    .B1(net2186));
 sg13g2_nand2_2 _6835_ (.Y(_2451_),
    .A(net2191),
    .B(net1969));
 sg13g2_nand2_2 _6836_ (.Y(_2452_),
    .A(_1563_),
    .B(_2451_));
 sg13g2_o21ai_1 _6837_ (.B1(net1861),
    .Y(_2453_),
    .A1(_2450_),
    .A2(_2452_));
 sg13g2_nand3_1 _6838_ (.B(_1676_),
    .C(_2453_),
    .A(_1675_),
    .Y(_2454_));
 sg13g2_a22oi_1 _6839_ (.Y(_2455_),
    .B1(_2454_),
    .B2(net2051),
    .A2(_2449_),
    .A1(net1898));
 sg13g2_nor3_1 _6840_ (.A(_1710_),
    .B(_1759_),
    .C(_2331_),
    .Y(_2456_));
 sg13g2_o21ai_1 _6841_ (.B1(_2456_),
    .Y(_2457_),
    .A1(net1959),
    .A2(_2079_));
 sg13g2_a21oi_2 _6842_ (.B1(_2000_),
    .Y(_2458_),
    .A2(_1763_),
    .A1(net1951));
 sg13g2_nand3_1 _6843_ (.B(net1987),
    .C(net1971),
    .A(net2131),
    .Y(_2459_));
 sg13g2_a22oi_1 _6844_ (.Y(_2460_),
    .B1(_2147_),
    .B2(_2459_),
    .A2(_1903_),
    .A1(net1846));
 sg13g2_o21ai_1 _6845_ (.B1(_2460_),
    .Y(_2461_),
    .A1(net1929),
    .A2(_2458_));
 sg13g2_a22oi_1 _6846_ (.Y(_2462_),
    .B1(_2461_),
    .B2(net2167),
    .A2(_2457_),
    .A1(net1839));
 sg13g2_o21ai_1 _6847_ (.B1(net1858),
    .Y(_2463_),
    .A1(net1959),
    .A2(net1841));
 sg13g2_a21oi_1 _6848_ (.A1(net1885),
    .A2(net1959),
    .Y(_2464_),
    .B1(net1888));
 sg13g2_o21ai_1 _6849_ (.B1(_2463_),
    .Y(_2465_),
    .A1(net2199),
    .A2(_1872_));
 sg13g2_o21ai_1 _6850_ (.B1(net1950),
    .Y(_2466_),
    .A1(_2464_),
    .A2(_2465_));
 sg13g2_a22oi_1 _6851_ (.Y(_2467_),
    .B1(_1837_),
    .B2(net1965),
    .A2(_1816_),
    .A1(net1796));
 sg13g2_o21ai_1 _6852_ (.B1(_2466_),
    .Y(_2468_),
    .A1(net1904),
    .A2(_2467_));
 sg13g2_nor2_1 _6853_ (.A(_1888_),
    .B(_2468_),
    .Y(_2469_));
 sg13g2_nor2_1 _6854_ (.A(_2462_),
    .B(_2469_),
    .Y(_2470_));
 sg13g2_nor2_1 _6855_ (.A(_1857_),
    .B(_2470_),
    .Y(_2471_));
 sg13g2_nand2_1 _6856_ (.Y(_2472_),
    .A(net2033),
    .B(net1864));
 sg13g2_a21oi_1 _6857_ (.A1(_2057_),
    .A2(_2472_),
    .Y(_2473_),
    .B1(net1937));
 sg13g2_nand2_2 _6858_ (.Y(_2474_),
    .A(net2034),
    .B(net1835));
 sg13g2_o21ai_1 _6859_ (.B1(_1872_),
    .Y(_2475_),
    .A1(net1856),
    .A2(net1835));
 sg13g2_a221oi_1 _6860_ (.B2(_2475_),
    .C1(_2473_),
    .B1(_2474_),
    .A1(net1994),
    .Y(_2476_),
    .A2(_2252_));
 sg13g2_a21oi_1 _6861_ (.A1(net1790),
    .A2(_2173_),
    .Y(_2477_),
    .B1(_0090_));
 sg13g2_o21ai_1 _6862_ (.B1(_2172_),
    .Y(_2478_),
    .A1(net1878),
    .A2(_1795_));
 sg13g2_nand2_1 _6863_ (.Y(_2479_),
    .A(net1983),
    .B(_2173_));
 sg13g2_nand4_1 _6864_ (.B(_2477_),
    .C(_2478_),
    .A(_2269_),
    .Y(_2480_),
    .D(_2479_));
 sg13g2_o21ai_1 _6865_ (.B1(net2052),
    .Y(_2481_),
    .A1(_2178_),
    .A2(_2480_));
 sg13g2_o21ai_1 _6866_ (.B1(_2481_),
    .Y(_2482_),
    .A1(net1895),
    .A2(_2476_));
 sg13g2_o21ai_1 _6867_ (.B1(_1655_),
    .Y(_2483_),
    .A1(net1880),
    .A2(_1559_));
 sg13g2_nand2_1 _6868_ (.Y(_2484_),
    .A(_1629_),
    .B(_2483_));
 sg13g2_nand3b_1 _6869_ (.B(net1909),
    .C(net1799),
    .Y(_2485_),
    .A_N(_2070_));
 sg13g2_nand4_1 _6870_ (.B(_2477_),
    .C(_2484_),
    .A(_2309_),
    .Y(_2486_),
    .D(_2485_));
 sg13g2_a21oi_1 _6871_ (.A1(net1877),
    .A2(_1632_),
    .Y(_2487_),
    .B1(net1893));
 sg13g2_o21ai_1 _6872_ (.B1(_2487_),
    .Y(_2488_),
    .A1(_1632_),
    .A2(_1836_));
 sg13g2_nand3_1 _6873_ (.B(net2163),
    .C(_2246_),
    .A(net2158),
    .Y(_2489_));
 sg13g2_nand3_1 _6874_ (.B(_2488_),
    .C(_2489_),
    .A(net1730),
    .Y(_2490_));
 sg13g2_a21oi_1 _6875_ (.A1(net2051),
    .A2(_2486_),
    .Y(_2491_),
    .B1(_2490_));
 sg13g2_nand2b_1 _6876_ (.Y(_2492_),
    .B(net2147),
    .A_N(_0096_));
 sg13g2_and2_1 _6877_ (.A(_1818_),
    .B(_2492_),
    .X(_2493_));
 sg13g2_a21o_1 _6878_ (.A2(_2493_),
    .A1(net2231),
    .B1(_1829_),
    .X(_2494_));
 sg13g2_o21ai_1 _6879_ (.B1(_2100_),
    .Y(_2495_),
    .A1(_1670_),
    .A2(_2280_));
 sg13g2_a21oi_1 _6880_ (.A1(net1866),
    .A2(net1850),
    .Y(_2496_),
    .B1(_2495_));
 sg13g2_o21ai_1 _6881_ (.B1(_2496_),
    .Y(_2497_),
    .A1(net1844),
    .A2(_2494_));
 sg13g2_nand2_1 _6882_ (.Y(_2498_),
    .A(net2047),
    .B(_2497_));
 sg13g2_o21ai_1 _6883_ (.B1(_2498_),
    .Y(_2499_),
    .A1(_1836_),
    .A2(_2026_));
 sg13g2_a21o_1 _6884_ (.A2(_2078_),
    .A1(net2227),
    .B1(_1687_),
    .X(_2500_));
 sg13g2_a21oi_1 _6885_ (.A1(net1912),
    .A2(_2500_),
    .Y(_2501_),
    .B1(_1811_));
 sg13g2_a221oi_1 _6886_ (.B2(net2199),
    .C1(_1904_),
    .B1(_2238_),
    .A1(net1987),
    .Y(_2502_),
    .A2(_1815_));
 sg13g2_o21ai_1 _6887_ (.B1(_2501_),
    .Y(_2503_),
    .A1(net2039),
    .A2(_2502_));
 sg13g2_a21oi_1 _6888_ (.A1(net2039),
    .A2(_1989_),
    .Y(_2504_),
    .B1(_2503_));
 sg13g2_a21oi_1 _6889_ (.A1(net1898),
    .A2(_2499_),
    .Y(_2505_),
    .B1(_2504_));
 sg13g2_nor2b_1 _6890_ (.A(_2505_),
    .B_N(net1742),
    .Y(_2506_));
 sg13g2_nand2_1 _6891_ (.Y(_2507_),
    .A(_3963_),
    .B(net995));
 sg13g2_nand2_1 _6892_ (.Y(_2508_),
    .A(net2036),
    .B(net1795));
 sg13g2_o21ai_1 _6893_ (.B1(net2021),
    .Y(_2509_),
    .A1(net2246),
    .A2(net2137));
 sg13g2_nand2_1 _6894_ (.Y(_2510_),
    .A(_1576_),
    .B(_2509_));
 sg13g2_nand3_1 _6895_ (.B(_2508_),
    .C(_2510_),
    .A(_1758_),
    .Y(_2511_));
 sg13g2_nand2_2 _6896_ (.Y(_2512_),
    .A(_1554_),
    .B(_1721_));
 sg13g2_a21oi_1 _6897_ (.A1(_1843_),
    .A2(_2512_),
    .Y(_2513_),
    .B1(net1930));
 sg13g2_nor3_1 _6898_ (.A(_1484_),
    .B(net1868),
    .C(net1844),
    .Y(_2514_));
 sg13g2_or3_1 _6899_ (.A(_2285_),
    .B(_2513_),
    .C(_2514_),
    .X(_2515_));
 sg13g2_a22oi_1 _6900_ (.Y(_2516_),
    .B1(_2515_),
    .B2(net2179),
    .A2(_2511_),
    .A1(net1840));
 sg13g2_o21ai_1 _6901_ (.B1(_1669_),
    .Y(_2517_),
    .A1(_1763_),
    .A2(_1929_));
 sg13g2_nand2_1 _6902_ (.Y(_2518_),
    .A(net2196),
    .B(_2271_));
 sg13g2_o21ai_1 _6903_ (.B1(_2518_),
    .Y(_2519_),
    .A1(net2196),
    .A2(_1576_));
 sg13g2_a21oi_1 _6904_ (.A1(_2517_),
    .A2(_2519_),
    .Y(_2520_),
    .B1(net2179));
 sg13g2_nor2_1 _6905_ (.A(net1886),
    .B(_2025_),
    .Y(_2521_));
 sg13g2_a21oi_1 _6906_ (.A1(net1842),
    .A2(_1799_),
    .Y(_2522_),
    .B1(_1546_));
 sg13g2_nor4_1 _6907_ (.A(_1736_),
    .B(_2520_),
    .C(_2521_),
    .D(_2522_),
    .Y(_2523_));
 sg13g2_o21ai_1 _6908_ (.B1(_1698_),
    .Y(_2524_),
    .A1(_2516_),
    .A2(_2523_));
 sg13g2_nand2_1 _6909_ (.Y(_2525_),
    .A(net2046),
    .B(_1692_));
 sg13g2_nor2_1 _6910_ (.A(_1993_),
    .B(_2525_),
    .Y(_2526_));
 sg13g2_a221oi_1 _6911_ (.B2(net1851),
    .C1(_2526_),
    .B1(_2127_),
    .A1(net1874),
    .Y(_2527_),
    .A2(net1794));
 sg13g2_nand2b_1 _6912_ (.Y(_2528_),
    .B(_2114_),
    .A_N(_2527_));
 sg13g2_nor2_1 _6913_ (.A(net2166),
    .B(_2195_),
    .Y(_2529_));
 sg13g2_a21oi_1 _6914_ (.A1(_1966_),
    .A2(_2104_),
    .Y(_2530_),
    .B1(_2101_));
 sg13g2_a21o_1 _6915_ (.A2(_2529_),
    .A1(_1586_),
    .B1(_2530_),
    .X(_2531_));
 sg13g2_a221oi_1 _6916_ (.B2(net1898),
    .C1(_2111_),
    .B1(_2531_),
    .A1(net2051),
    .Y(_2532_),
    .A2(_2528_));
 sg13g2_nand2_2 _6917_ (.Y(_2533_),
    .A(_1512_),
    .B(net1849));
 sg13g2_inv_1 _6918_ (.Y(_2534_),
    .A(_2533_));
 sg13g2_nand3_1 _6919_ (.B(_1944_),
    .C(_2533_),
    .A(_1784_),
    .Y(_2535_));
 sg13g2_nand2_1 _6920_ (.Y(_2536_),
    .A(_2363_),
    .B(_2535_));
 sg13g2_o21ai_1 _6921_ (.B1(net2181),
    .Y(_2537_),
    .A1(_2417_),
    .A2(_2536_));
 sg13g2_a21oi_1 _6922_ (.A1(net2028),
    .A2(_1649_),
    .Y(_2538_),
    .B1(_2205_));
 sg13g2_a221oi_1 _6923_ (.B2(_2538_),
    .C1(net1888),
    .B1(_2415_),
    .A1(net1882),
    .Y(_2539_),
    .A2(net1796));
 sg13g2_nor3_1 _6924_ (.A(net1976),
    .B(_1748_),
    .C(_2366_),
    .Y(_2540_));
 sg13g2_o21ai_1 _6925_ (.B1(_2537_),
    .Y(_2541_),
    .A1(net1856),
    .A2(_2540_));
 sg13g2_o21ai_1 _6926_ (.B1(net1901),
    .Y(_2542_),
    .A1(_2539_),
    .A2(_2541_));
 sg13g2_nand3_1 _6927_ (.B(_1906_),
    .C(_2264_),
    .A(net1859),
    .Y(_2543_));
 sg13g2_nand3_1 _6928_ (.B(_1574_),
    .C(_1851_),
    .A(net1994),
    .Y(_2544_));
 sg13g2_nand3_1 _6929_ (.B(_2543_),
    .C(_2544_),
    .A(_2353_),
    .Y(_2545_));
 sg13g2_a21oi_1 _6930_ (.A1(_1399_),
    .A2(net1984),
    .Y(_2546_),
    .B1(net1880));
 sg13g2_a21oi_2 _6931_ (.B1(net1940),
    .Y(_2547_),
    .A2(_2546_),
    .A1(net1855));
 sg13g2_a21oi_1 _6932_ (.A1(_2545_),
    .A2(_2547_),
    .Y(_2548_),
    .B1(_2372_));
 sg13g2_a21oi_1 _6933_ (.A1(_2542_),
    .A2(_2548_),
    .Y(_2549_),
    .B1(_1899_));
 sg13g2_a21oi_1 _6934_ (.A1(net1731),
    .A2(_2532_),
    .Y(_2550_),
    .B1(_2507_));
 sg13g2_a22oi_1 _6935_ (.Y(_2551_),
    .B1(_2455_),
    .B2(_1672_),
    .A2(_2430_),
    .A1(_1747_));
 sg13g2_o21ai_1 _6936_ (.B1(_2524_),
    .Y(_2552_),
    .A1(_1503_),
    .A2(_2482_));
 sg13g2_nor4_1 _6937_ (.A(_2471_),
    .B(_2491_),
    .C(_2506_),
    .D(_2552_),
    .Y(_2553_));
 sg13g2_nor3_2 _6938_ (.A(_2414_),
    .B(_2447_),
    .C(_2549_),
    .Y(_2554_));
 sg13g2_and3_1 _6939_ (.X(_2555_),
    .A(_2551_),
    .B(_2553_),
    .C(_2554_));
 sg13g2_and2_1 _6940_ (.A(_2550_),
    .B(_2555_),
    .X(_2556_));
 sg13g2_a21oi_1 _6941_ (.A1(net2143),
    .A2(net1867),
    .Y(_2557_),
    .B1(net2210));
 sg13g2_o21ai_1 _6942_ (.B1(_1577_),
    .Y(_2558_),
    .A1(_1515_),
    .A2(_1763_));
 sg13g2_o21ai_1 _6943_ (.B1(net2042),
    .Y(_2559_),
    .A1(_2557_),
    .A2(_2558_));
 sg13g2_a21oi_1 _6944_ (.A1(net1805),
    .A2(net1850),
    .Y(_2560_),
    .B1(net2181));
 sg13g2_o21ai_1 _6945_ (.B1(net1845),
    .Y(_2561_),
    .A1(_1656_),
    .A2(_2045_));
 sg13g2_nand3_1 _6946_ (.B(_2560_),
    .C(_2561_),
    .A(_2559_),
    .Y(_2562_));
 sg13g2_o21ai_1 _6947_ (.B1(_2562_),
    .Y(_2563_),
    .A1(net1797),
    .A2(_2026_));
 sg13g2_a21oi_1 _6948_ (.A1(net1989),
    .A2(net1801),
    .Y(_2564_),
    .B1(_2278_));
 sg13g2_and2_1 _6949_ (.A(_1593_),
    .B(_1827_),
    .X(_2565_));
 sg13g2_nand2_1 _6950_ (.Y(_2566_),
    .A(_1593_),
    .B(_1827_));
 sg13g2_a22oi_1 _6951_ (.Y(_2567_),
    .B1(_2566_),
    .B2(_1522_),
    .A2(_1913_),
    .A1(net1947));
 sg13g2_a221oi_1 _6952_ (.B2(net2025),
    .C1(net2196),
    .B1(net1808),
    .A1(net2221),
    .Y(_2568_),
    .A2(net1886));
 sg13g2_nor3_1 _6953_ (.A(net2179),
    .B(_2355_),
    .C(_2568_),
    .Y(_2569_));
 sg13g2_o21ai_1 _6954_ (.B1(_2569_),
    .Y(_2570_),
    .A1(net1844),
    .A2(_2567_));
 sg13g2_o21ai_1 _6955_ (.B1(_2570_),
    .Y(_2571_),
    .A1(_2025_),
    .A2(_2564_));
 sg13g2_a22oi_1 _6956_ (.Y(_2572_),
    .B1(_2571_),
    .B2(net1742),
    .A2(_2563_),
    .A1(net1729));
 sg13g2_nor2_1 _6957_ (.A(net1893),
    .B(_2572_),
    .Y(_2573_));
 sg13g2_o21ai_1 _6958_ (.B1(_1953_),
    .Y(_2574_),
    .A1(net1948),
    .A2(_1699_));
 sg13g2_nand2b_2 _6959_ (.Y(_2575_),
    .B(_2086_),
    .A_N(_1931_));
 sg13g2_a22oi_1 _6960_ (.Y(_2576_),
    .B1(_2575_),
    .B2(net1912),
    .A2(_1960_),
    .A1(net1927));
 sg13g2_nand3_1 _6961_ (.B(net1802),
    .C(net1854),
    .A(net1959),
    .Y(_2577_));
 sg13g2_a21oi_1 _6962_ (.A1(_1631_),
    .A2(_1673_),
    .Y(_2578_),
    .B1(_2148_));
 sg13g2_nand2_1 _6963_ (.Y(_2579_),
    .A(_2577_),
    .B(_2578_));
 sg13g2_nand2_1 _6964_ (.Y(_2580_),
    .A(net1987),
    .B(net1802));
 sg13g2_nand2b_1 _6965_ (.Y(_2581_),
    .B(_2580_),
    .A_N(_2053_));
 sg13g2_a21oi_1 _6966_ (.A1(net1858),
    .A2(_2581_),
    .Y(_2582_),
    .B1(_2579_));
 sg13g2_o21ai_1 _6967_ (.B1(_2582_),
    .Y(_2583_),
    .A1(net2174),
    .A2(_2576_));
 sg13g2_nor2_1 _6968_ (.A(net1931),
    .B(_2185_),
    .Y(_2584_));
 sg13g2_a21oi_1 _6969_ (.A1(net1802),
    .A2(net1931),
    .Y(_2585_),
    .B1(_2584_));
 sg13g2_nor2_2 _6970_ (.A(_1538_),
    .B(net1856),
    .Y(_2586_));
 sg13g2_nand2b_1 _6971_ (.Y(_2587_),
    .B(_2237_),
    .A_N(_2127_));
 sg13g2_nor2_1 _6972_ (.A(net2169),
    .B(_2587_),
    .Y(_2588_));
 sg13g2_nor3_1 _6973_ (.A(net2160),
    .B(_2586_),
    .C(_2588_),
    .Y(_2589_));
 sg13g2_o21ai_1 _6974_ (.B1(_2589_),
    .Y(_2590_),
    .A1(net2048),
    .A2(_2585_));
 sg13g2_a221oi_1 _6975_ (.B2(net2052),
    .C1(_2574_),
    .B1(_2590_),
    .A1(net1900),
    .Y(_2591_),
    .A2(_2583_));
 sg13g2_a21o_1 _6976_ (.A2(_2341_),
    .A1(_1860_),
    .B1(net2206),
    .X(_2592_));
 sg13g2_o21ai_1 _6977_ (.B1(net1960),
    .Y(_2593_),
    .A1(net2030),
    .A2(_1402_));
 sg13g2_or2_1 _6978_ (.X(_2594_),
    .B(_1769_),
    .A(net2236));
 sg13g2_a21oi_1 _6979_ (.A1(net2233),
    .A2(_1402_),
    .Y(_2595_),
    .B1(net2206));
 sg13g2_a22oi_1 _6980_ (.Y(_2596_),
    .B1(_2594_),
    .B2(_2595_),
    .A2(_2593_),
    .A1(_1922_));
 sg13g2_o21ai_1 _6981_ (.B1(net2171),
    .Y(_2597_),
    .A1(net2039),
    .A2(_2596_));
 sg13g2_a21oi_1 _6982_ (.A1(_2228_),
    .A2(_2592_),
    .Y(_2598_),
    .B1(_2597_));
 sg13g2_o21ai_1 _6983_ (.B1(net2243),
    .Y(_2599_),
    .A1(_1570_),
    .A2(_1594_));
 sg13g2_nand2b_1 _6984_ (.Y(_2600_),
    .B(net2031),
    .A_N(_2599_));
 sg13g2_a21oi_1 _6985_ (.A1(net1965),
    .A2(net1797),
    .Y(_2601_),
    .B1(net2185));
 sg13g2_or2_1 _6986_ (.X(_2602_),
    .B(_2019_),
    .A(net2235));
 sg13g2_a21oi_1 _6987_ (.A1(net1986),
    .A2(_1889_),
    .Y(_2603_),
    .B1(net1940));
 sg13g2_nand4_1 _6988_ (.B(_2601_),
    .C(_2602_),
    .A(_2600_),
    .Y(_2604_),
    .D(_2603_));
 sg13g2_a21oi_1 _6989_ (.A1(net1839),
    .A2(_2604_),
    .Y(_2605_),
    .B1(_2598_));
 sg13g2_nand2_2 _6990_ (.Y(_2606_),
    .A(net2204),
    .B(_2494_));
 sg13g2_a21oi_1 _6991_ (.A1(net2130),
    .A2(net1985),
    .Y(_2607_),
    .B1(_1496_));
 sg13g2_nand2_1 _6992_ (.Y(_2608_),
    .A(_2606_),
    .B(_2607_));
 sg13g2_a21o_1 _6993_ (.A2(net1852),
    .A1(net1996),
    .B1(_1736_),
    .X(_2609_));
 sg13g2_nand2_1 _6994_ (.Y(_2610_),
    .A(net2208),
    .B(_1891_));
 sg13g2_a221oi_1 _6995_ (.B2(_1889_),
    .C1(net2189),
    .B1(net1955),
    .A1(_1402_),
    .Y(_2611_),
    .A2(net1986));
 sg13g2_a22oi_1 _6996_ (.Y(_2612_),
    .B1(_2610_),
    .B2(_2611_),
    .A2(_2394_),
    .A1(net2189));
 sg13g2_a221oi_1 _6997_ (.B2(net2047),
    .C1(_2609_),
    .B1(_2612_),
    .A1(net1907),
    .Y(_2613_),
    .A2(_2608_));
 sg13g2_o21ai_1 _6998_ (.B1(_1698_),
    .Y(_2614_),
    .A1(_2605_),
    .A2(_2613_));
 sg13g2_a21oi_1 _6999_ (.A1(net1847),
    .A2(_1889_),
    .Y(_2615_),
    .B1(net2184));
 sg13g2_nand2_1 _7000_ (.Y(_2616_),
    .A(net1967),
    .B(_1891_));
 sg13g2_a21oi_1 _7001_ (.A1(_2615_),
    .A2(_2616_),
    .Y(_2617_),
    .B1(net2181));
 sg13g2_nor3_1 _7002_ (.A(_1481_),
    .B(_1490_),
    .C(_1753_),
    .Y(_2618_));
 sg13g2_a21oi_1 _7003_ (.A1(net1866),
    .A2(_1636_),
    .Y(_2619_),
    .B1(net1905));
 sg13g2_o21ai_1 _7004_ (.B1(_2619_),
    .Y(_2620_),
    .A1(net1848),
    .A2(_1891_));
 sg13g2_o21ai_1 _7005_ (.B1(_2620_),
    .Y(_2621_),
    .A1(net1935),
    .A2(_2120_));
 sg13g2_nor4_2 _7006_ (.A(net1940),
    .B(_2617_),
    .C(_2618_),
    .Y(_2622_),
    .D(_2621_));
 sg13g2_a221oi_1 _7007_ (.B2(_2047_),
    .C1(net2195),
    .B1(_1901_),
    .A1(net2219),
    .Y(_2623_),
    .A2(net1799));
 sg13g2_nor3_1 _7008_ (.A(net2042),
    .B(_1491_),
    .C(_1615_),
    .Y(_2624_));
 sg13g2_nor3_1 _7009_ (.A(net2180),
    .B(_2623_),
    .C(_2624_),
    .Y(_2625_));
 sg13g2_nor3_1 _7010_ (.A(net1983),
    .B(_1570_),
    .C(_1594_),
    .Y(_2626_));
 sg13g2_o21ai_1 _7011_ (.B1(net1901),
    .Y(_2627_),
    .A1(net1935),
    .A2(_2626_));
 sg13g2_nand2_1 _7012_ (.Y(_2628_),
    .A(net1963),
    .B(_2112_));
 sg13g2_and2_1 _7013_ (.A(_2599_),
    .B(_2628_),
    .X(_2629_));
 sg13g2_nor2_1 _7014_ (.A(net1905),
    .B(_2629_),
    .Y(_2630_));
 sg13g2_nor3_1 _7015_ (.A(net1905),
    .B(_2070_),
    .C(_2629_),
    .Y(_2631_));
 sg13g2_nor3_1 _7016_ (.A(_2625_),
    .B(_2627_),
    .C(_2631_),
    .Y(_2632_));
 sg13g2_o21ai_1 _7017_ (.B1(_1747_),
    .Y(_2633_),
    .A1(_2622_),
    .A2(_2632_));
 sg13g2_a21o_1 _7018_ (.A2(_1621_),
    .A1(_1580_),
    .B1(net2191),
    .X(_2634_));
 sg13g2_a21oi_1 _7019_ (.A1(_2166_),
    .A2(_2634_),
    .Y(_2635_),
    .B1(net2178));
 sg13g2_nor2_2 _7020_ (.A(net2177),
    .B(net1939),
    .Y(_2636_));
 sg13g2_a21oi_1 _7021_ (.A1(net1987),
    .A2(net1879),
    .Y(_2637_),
    .B1(_1759_));
 sg13g2_a21oi_1 _7022_ (.A1(net1788),
    .A2(_2637_),
    .Y(_2638_),
    .B1(_2636_));
 sg13g2_nor4_2 _7023_ (.A(_0091_),
    .B(net2198),
    .C(net2185),
    .Y(_2639_),
    .D(net1894));
 sg13g2_o21ai_1 _7024_ (.B1(net1788),
    .Y(_2640_),
    .A1(_1926_),
    .A2(_2639_));
 sg13g2_o21ai_1 _7025_ (.B1(_2640_),
    .Y(_2641_),
    .A1(_2635_),
    .A2(_2638_));
 sg13g2_nand2_1 _7026_ (.Y(_2642_),
    .A(net1730),
    .B(_2641_));
 sg13g2_o21ai_1 _7027_ (.B1(net2169),
    .Y(_2643_),
    .A1(_1670_),
    .A2(_1864_));
 sg13g2_nand2_2 _7028_ (.Y(_2644_),
    .A(net1900),
    .B(_2643_));
 sg13g2_a21oi_1 _7029_ (.A1(_1863_),
    .A2(_1993_),
    .Y(_2645_),
    .B1(net2168));
 sg13g2_a21oi_1 _7030_ (.A1(_2130_),
    .A2(_2645_),
    .Y(_2646_),
    .B1(_2644_));
 sg13g2_nand3_1 _7031_ (.B(_1758_),
    .C(_2127_),
    .A(net2046),
    .Y(_2647_));
 sg13g2_o21ai_1 _7032_ (.B1(_2647_),
    .Y(_2648_),
    .A1(_1586_),
    .A2(net1839));
 sg13g2_o21ai_1 _7033_ (.B1(_1668_),
    .Y(_2649_),
    .A1(_2646_),
    .A2(_2648_));
 sg13g2_nand4_1 _7034_ (.B(_2633_),
    .C(_2642_),
    .A(_2614_),
    .Y(_2650_),
    .D(_2649_));
 sg13g2_nor3_2 _7035_ (.A(_2573_),
    .B(_2591_),
    .C(_2650_),
    .Y(_2651_));
 sg13g2_nand2_1 _7036_ (.Y(_2652_),
    .A(net2230),
    .B(net2145));
 sg13g2_nand2_1 _7037_ (.Y(_2653_),
    .A(_2341_),
    .B(_2652_));
 sg13g2_a22oi_1 _7038_ (.Y(_2654_),
    .B1(_2378_),
    .B2(_1782_),
    .A2(net1836),
    .A1(net1985));
 sg13g2_a221oi_1 _7039_ (.B2(net1928),
    .C1(_2654_),
    .B1(_2653_),
    .A1(net1912),
    .Y(_2655_),
    .A2(_1815_));
 sg13g2_a21oi_1 _7040_ (.A1(_2273_),
    .A2(_2652_),
    .Y(_2656_),
    .B1(_1670_));
 sg13g2_o21ai_1 _7041_ (.B1(_1754_),
    .Y(_2657_),
    .A1(net1913),
    .A2(_1781_));
 sg13g2_o21ai_1 _7042_ (.B1(_2657_),
    .Y(_2658_),
    .A1(_1527_),
    .A2(_1624_));
 sg13g2_nor2_2 _7043_ (.A(_2656_),
    .B(_2658_),
    .Y(_2659_));
 sg13g2_a22oi_1 _7044_ (.Y(_2660_),
    .B1(_2659_),
    .B2(_1667_),
    .A2(_2655_),
    .A1(_1697_));
 sg13g2_or2_1 _7045_ (.X(_2661_),
    .B(_2660_),
    .A(_0091_));
 sg13g2_nor2_2 _7046_ (.A(net1955),
    .B(net1847),
    .Y(_2662_));
 sg13g2_a21oi_1 _7047_ (.A1(_1571_),
    .A2(net1833),
    .Y(_2663_),
    .B1(_2662_));
 sg13g2_a21oi_1 _7048_ (.A1(net1986),
    .A2(_2102_),
    .Y(_2664_),
    .B1(_2663_));
 sg13g2_nand3_1 _7049_ (.B(net1842),
    .C(_2280_),
    .A(_1571_),
    .Y(_2665_));
 sg13g2_nand3_1 _7050_ (.B(_1700_),
    .C(net1833),
    .A(net1985),
    .Y(_2666_));
 sg13g2_a21oi_1 _7051_ (.A1(net1981),
    .A2(_1506_),
    .Y(_2667_),
    .B1(net1902));
 sg13g2_nand2_1 _7052_ (.Y(_2668_),
    .A(_1631_),
    .B(_1828_));
 sg13g2_a21oi_1 _7053_ (.A1(net2204),
    .A2(_0096_),
    .Y(_2669_),
    .B1(net2184));
 sg13g2_o21ai_1 _7054_ (.B1(_2668_),
    .Y(_2670_),
    .A1(net2172),
    .A2(_2669_));
 sg13g2_a221oi_1 _7055_ (.B2(_2667_),
    .C1(_2670_),
    .B1(_2666_),
    .A1(_1480_),
    .Y(_2671_),
    .A2(_2665_));
 sg13g2_o21ai_1 _7056_ (.B1(_2671_),
    .Y(_2672_),
    .A1(net1932),
    .A2(_2664_));
 sg13g2_o21ai_1 _7057_ (.B1(_2661_),
    .Y(_2673_),
    .A1(_1601_),
    .A2(_2672_));
 sg13g2_nand3_1 _7058_ (.B(net1942),
    .C(_2673_),
    .A(_1462_),
    .Y(_2674_));
 sg13g2_nand2_1 _7059_ (.Y(_2675_),
    .A(_1645_),
    .B(_1955_));
 sg13g2_o21ai_1 _7060_ (.B1(_1823_),
    .Y(_2676_),
    .A1(net2025),
    .A2(net1880));
 sg13g2_nand2_1 _7061_ (.Y(_2677_),
    .A(net1968),
    .B(_2676_));
 sg13g2_nand3_1 _7062_ (.B(_1571_),
    .C(_2676_),
    .A(net2209),
    .Y(_2678_));
 sg13g2_a21oi_1 _7063_ (.A1(_1603_),
    .A2(_1636_),
    .Y(_2679_),
    .B1(_2675_));
 sg13g2_o21ai_1 _7064_ (.B1(_2679_),
    .Y(_2680_),
    .A1(_1570_),
    .A2(_2677_));
 sg13g2_o21ai_1 _7065_ (.B1(net2192),
    .Y(_2681_),
    .A1(net2213),
    .A2(_2271_));
 sg13g2_o21ai_1 _7066_ (.B1(_2680_),
    .Y(_2682_),
    .A1(_1713_),
    .A2(_2681_));
 sg13g2_o21ai_1 _7067_ (.B1(net1953),
    .Y(_2683_),
    .A1(net2143),
    .A2(net1964));
 sg13g2_o21ai_1 _7068_ (.B1(net2175),
    .Y(_2684_),
    .A1(_2452_),
    .A2(_2683_));
 sg13g2_o21ai_1 _7069_ (.B1(_2684_),
    .Y(_2685_),
    .A1(net2176),
    .A2(_2682_));
 sg13g2_o21ai_1 _7070_ (.B1(net2052),
    .Y(_2686_),
    .A1(_0090_),
    .A2(_2685_));
 sg13g2_nand2_1 _7071_ (.Y(_2687_),
    .A(net1849),
    .B(_2676_));
 sg13g2_nand2_2 _7072_ (.Y(_2688_),
    .A(_1909_),
    .B(_2687_));
 sg13g2_a21oi_1 _7073_ (.A1(net1994),
    .A2(_2688_),
    .Y(_2689_),
    .B1(net2164));
 sg13g2_o21ai_1 _7074_ (.B1(_1669_),
    .Y(_2690_),
    .A1(_1512_),
    .A2(_1795_));
 sg13g2_a22oi_1 _7075_ (.Y(_2691_),
    .B1(_2240_),
    .B2(_2280_),
    .A2(net1787),
    .A1(net1845));
 sg13g2_nand2_1 _7076_ (.Y(_2692_),
    .A(_2690_),
    .B(_2691_));
 sg13g2_a21oi_1 _7077_ (.A1(net1962),
    .A2(_2271_),
    .Y(_2693_),
    .B1(net1935));
 sg13g2_nand2_1 _7078_ (.Y(_2694_),
    .A(net2221),
    .B(_1499_));
 sg13g2_o21ai_1 _7079_ (.B1(_2693_),
    .Y(_2695_),
    .A1(net1972),
    .A2(net1962));
 sg13g2_a21oi_1 _7080_ (.A1(net1989),
    .A2(net1954),
    .Y(_2696_),
    .B1(_2278_));
 sg13g2_a22oi_1 _7081_ (.Y(_2697_),
    .B1(_2696_),
    .B2(net1910),
    .A2(_2692_),
    .A1(net2049));
 sg13g2_nand3_1 _7082_ (.B(_2695_),
    .C(_2697_),
    .A(_2689_),
    .Y(_2698_));
 sg13g2_o21ai_1 _7083_ (.B1(_1768_),
    .Y(_2699_),
    .A1(net2149),
    .A2(_0096_));
 sg13g2_inv_1 _7084_ (.Y(_2700_),
    .A(_2699_));
 sg13g2_nand3_1 _7085_ (.B(net1814),
    .C(_2699_),
    .A(net2164),
    .Y(_2701_));
 sg13g2_nand3_1 _7086_ (.B(_2698_),
    .C(_2701_),
    .A(net2159),
    .Y(_2702_));
 sg13g2_and3_2 _7087_ (.X(_2703_),
    .A(_1479_),
    .B(_2686_),
    .C(_2702_));
 sg13g2_o21ai_1 _7088_ (.B1(net2196),
    .Y(_2704_),
    .A1(net2221),
    .A2(net1952));
 sg13g2_o21ai_1 _7089_ (.B1(net2241),
    .Y(_2705_),
    .A1(net1866),
    .A2(_1737_));
 sg13g2_nor2_1 _7090_ (.A(net2179),
    .B(_2012_),
    .Y(_2706_));
 sg13g2_a221oi_1 _7091_ (.B2(_2706_),
    .C1(net2036),
    .B1(_2705_),
    .A1(net2179),
    .Y(_2707_),
    .A2(_2174_));
 sg13g2_nand2_1 _7092_ (.Y(_2708_),
    .A(net1968),
    .B(net1952));
 sg13g2_o21ai_1 _7093_ (.B1(_2708_),
    .Y(_2709_),
    .A1(net1968),
    .A2(_2272_));
 sg13g2_a21oi_1 _7094_ (.A1(net1864),
    .A2(net1842),
    .Y(_2710_),
    .B1(net2220));
 sg13g2_nor3_1 _7095_ (.A(net1905),
    .B(_1713_),
    .C(_2710_),
    .Y(_2711_));
 sg13g2_a21oi_1 _7096_ (.A1(net1994),
    .A2(_2709_),
    .Y(_2712_),
    .B1(_2711_));
 sg13g2_o21ai_1 _7097_ (.B1(_2712_),
    .Y(_2713_),
    .A1(_2704_),
    .A2(_2707_));
 sg13g2_nand2_1 _7098_ (.Y(_2714_),
    .A(net2246),
    .B(_2272_));
 sg13g2_a22oi_1 _7099_ (.Y(_2715_),
    .B1(_2272_),
    .B2(net2246),
    .A2(_1777_),
    .A1(_1653_));
 sg13g2_nor2_1 _7100_ (.A(net2221),
    .B(_2156_),
    .Y(_2716_));
 sg13g2_nand2_1 _7101_ (.Y(_2717_),
    .A(net1884),
    .B(_1522_));
 sg13g2_a221oi_1 _7102_ (.B2(_2717_),
    .C1(net1936),
    .B1(_2716_),
    .A1(net2220),
    .Y(_2718_),
    .A2(_2715_));
 sg13g2_nand2_1 _7103_ (.Y(_2719_),
    .A(_2533_),
    .B(_2677_));
 sg13g2_nor3_1 _7104_ (.A(net1946),
    .B(_2047_),
    .C(_2719_),
    .Y(_2720_));
 sg13g2_nor2_1 _7105_ (.A(net1889),
    .B(_2720_),
    .Y(_2721_));
 sg13g2_nand3_1 _7106_ (.B(net1798),
    .C(net1795),
    .A(net2247),
    .Y(_2722_));
 sg13g2_a22oi_1 _7107_ (.Y(_2723_),
    .B1(_2291_),
    .B2(net1850),
    .A2(_1900_),
    .A1(_1781_));
 sg13g2_o21ai_1 _7108_ (.B1(_2722_),
    .Y(_2724_),
    .A1(net1906),
    .A2(_2192_));
 sg13g2_nor4_1 _7109_ (.A(net1940),
    .B(_2718_),
    .C(_2721_),
    .D(_2724_),
    .Y(_2725_));
 sg13g2_o21ai_1 _7110_ (.B1(_2725_),
    .Y(_2726_),
    .A1(net2180),
    .A2(_2723_));
 sg13g2_a22oi_1 _7111_ (.Y(_2727_),
    .B1(_2713_),
    .B2(net1901),
    .A2(_1926_),
    .A1(net1875));
 sg13g2_a21oi_2 _7112_ (.B1(_1899_),
    .Y(_2728_),
    .A2(_2727_),
    .A1(_2726_));
 sg13g2_o21ai_1 _7113_ (.B1(net2171),
    .Y(_2729_),
    .A1(_1782_),
    .A2(_2302_));
 sg13g2_nor2_2 _7114_ (.A(net1875),
    .B(_2599_),
    .Y(_2730_));
 sg13g2_o21ai_1 _7115_ (.B1(net2205),
    .Y(_2731_),
    .A1(_1829_),
    .A2(_2730_));
 sg13g2_nand2b_1 _7116_ (.Y(_2732_),
    .B(_2731_),
    .A_N(_1496_));
 sg13g2_nor2_1 _7117_ (.A(net2188),
    .B(_2732_),
    .Y(_2733_));
 sg13g2_nor2_1 _7118_ (.A(_2729_),
    .B(_2733_),
    .Y(_2734_));
 sg13g2_o21ai_1 _7119_ (.B1(net1954),
    .Y(_2735_),
    .A1(net2204),
    .A2(net2023));
 sg13g2_a221oi_1 _7120_ (.B2(_2735_),
    .C1(_1732_),
    .B1(net1860),
    .A1(net1992),
    .Y(_2736_),
    .A2(net1975));
 sg13g2_o21ai_1 _7121_ (.B1(_2736_),
    .Y(_2737_),
    .A1(net1932),
    .A2(_2732_));
 sg13g2_nor4_2 _7122_ (.A(net1894),
    .B(_1857_),
    .C(_2734_),
    .Y(_2738_),
    .D(_2737_));
 sg13g2_nor3_1 _7123_ (.A(_2703_),
    .B(_2728_),
    .C(_2738_),
    .Y(_2739_));
 sg13g2_nand3_1 _7124_ (.B(_2016_),
    .C(_2092_),
    .A(net2201),
    .Y(_2740_));
 sg13g2_nand2_1 _7125_ (.Y(_2741_),
    .A(_1394_),
    .B(_1547_));
 sg13g2_and2_1 _7126_ (.A(_2740_),
    .B(_2741_),
    .X(_2742_));
 sg13g2_nor2_1 _7127_ (.A(net1934),
    .B(net1835),
    .Y(_2743_));
 sg13g2_nor4_2 _7128_ (.A(net1939),
    .B(_2586_),
    .C(_2742_),
    .Y(_2744_),
    .D(_2743_));
 sg13g2_nand2_1 _7129_ (.Y(_2745_),
    .A(net1991),
    .B(_2382_));
 sg13g2_nand2_1 _7130_ (.Y(_2746_),
    .A(_2744_),
    .B(_2745_));
 sg13g2_o21ai_1 _7131_ (.B1(net1894),
    .Y(_2747_),
    .A1(_1864_),
    .A2(_1925_));
 sg13g2_o21ai_1 _7132_ (.B1(_1675_),
    .Y(_2748_),
    .A1(net1888),
    .A2(_2391_));
 sg13g2_nor2_1 _7133_ (.A(_1534_),
    .B(_1860_),
    .Y(_2749_));
 sg13g2_nand2b_2 _7134_ (.Y(_2750_),
    .B(_2093_),
    .A_N(_2749_));
 sg13g2_nor2_2 _7135_ (.A(net2043),
    .B(_1533_),
    .Y(_2751_));
 sg13g2_and2_1 _7136_ (.A(_2750_),
    .B(_2751_),
    .X(_2752_));
 sg13g2_a221oi_1 _7137_ (.B2(net2166),
    .C1(_2748_),
    .B1(_2752_),
    .A1(net1907),
    .Y(_2753_),
    .A2(_2395_));
 sg13g2_o21ai_1 _7138_ (.B1(_2747_),
    .Y(_2754_),
    .A1(net2162),
    .A2(_2753_));
 sg13g2_nand2_1 _7139_ (.Y(_2755_),
    .A(_2746_),
    .B(_2754_));
 sg13g2_a21oi_1 _7140_ (.A1(net1731),
    .A2(_2755_),
    .Y(_2756_),
    .B1(_2226_));
 sg13g2_and4_1 _7141_ (.A(_2651_),
    .B(_2674_),
    .C(_2739_),
    .D(_2756_),
    .X(_2757_));
 sg13g2_or2_1 _7142_ (.X(_2758_),
    .B(\draw_game_inst.board_x[1] ),
    .A(\draw_game_inst.board_x[0] ));
 sg13g2_a22oi_1 _7143_ (.Y(_2759_),
    .B1(_1771_),
    .B2(_1861_),
    .A2(net1797),
    .A1(net1847));
 sg13g2_nand3_1 _7144_ (.B(_1740_),
    .C(_2759_),
    .A(net1908),
    .Y(_2760_));
 sg13g2_a221oi_1 _7145_ (.B2(_1797_),
    .C1(net1857),
    .B1(net1956),
    .A1(net2207),
    .Y(_2761_),
    .A2(net2146));
 sg13g2_nand4_1 _7146_ (.B(_1574_),
    .C(_1645_),
    .A(net1995),
    .Y(_2762_),
    .D(_2678_));
 sg13g2_nor2_1 _7147_ (.A(net1974),
    .B(net1933),
    .Y(_2763_));
 sg13g2_a22oi_1 _7148_ (.Y(_2764_),
    .B1(_2763_),
    .B2(_1515_),
    .A2(_2761_),
    .A1(_2580_));
 sg13g2_nand3_1 _7149_ (.B(_2762_),
    .C(_2764_),
    .A(_2760_),
    .Y(_2765_));
 sg13g2_nand3_1 _7150_ (.B(_2054_),
    .C(_2634_),
    .A(_1880_),
    .Y(_2766_));
 sg13g2_o21ai_1 _7151_ (.B1(net1907),
    .Y(_2767_),
    .A1(net2201),
    .A2(net1837));
 sg13g2_nor3_1 _7152_ (.A(_1517_),
    .B(_1816_),
    .C(_2032_),
    .Y(_2768_));
 sg13g2_o21ai_1 _7153_ (.B1(net1854),
    .Y(_2769_),
    .A1(_1859_),
    .A2(_2768_));
 sg13g2_nand2_1 _7154_ (.Y(_2770_),
    .A(_2767_),
    .B(_2769_));
 sg13g2_a21oi_1 _7155_ (.A1(_2635_),
    .A2(_2766_),
    .Y(_2771_),
    .B1(_2770_));
 sg13g2_a22oi_1 _7156_ (.Y(_2772_),
    .B1(_2771_),
    .B2(_1602_),
    .A2(_2765_),
    .A1(_1479_));
 sg13g2_nor2_1 _7157_ (.A(net1938),
    .B(_2772_),
    .Y(_2773_));
 sg13g2_nand2_1 _7158_ (.Y(_2774_),
    .A(net1864),
    .B(net1833));
 sg13g2_nand2b_1 _7159_ (.Y(_2775_),
    .B(_2774_),
    .A_N(net2247));
 sg13g2_a21oi_1 _7160_ (.A1(net2244),
    .A2(_2700_),
    .Y(_2776_),
    .B1(_2044_));
 sg13g2_o21ai_1 _7161_ (.B1(_2693_),
    .Y(_2777_),
    .A1(net1962),
    .A2(_2774_));
 sg13g2_nand2_1 _7162_ (.Y(_2778_),
    .A(net1962),
    .B(_1900_));
 sg13g2_o21ai_1 _7163_ (.B1(_2778_),
    .Y(_2779_),
    .A1(net1964),
    .A2(net1806));
 sg13g2_o21ai_1 _7164_ (.B1(net1814),
    .Y(_2780_),
    .A1(_1507_),
    .A2(_1651_));
 sg13g2_o21ai_1 _7165_ (.B1(net1911),
    .Y(_2781_),
    .A1(_1576_),
    .A2(_1725_));
 sg13g2_nand3_1 _7166_ (.B(_2780_),
    .C(_2781_),
    .A(_2777_),
    .Y(_2782_));
 sg13g2_a21oi_1 _7167_ (.A1(net1860),
    .A2(_2779_),
    .Y(_2783_),
    .B1(_2782_));
 sg13g2_a22oi_1 _7168_ (.Y(_2784_),
    .B1(_2783_),
    .B2(_2689_),
    .A2(_2776_),
    .A1(_2775_));
 sg13g2_inv_1 _7169_ (.Y(_2785_),
    .A(_2784_));
 sg13g2_nand4_1 _7170_ (.B(net1814),
    .C(net1788),
    .A(net2163),
    .Y(_2786_),
    .D(_1922_));
 sg13g2_nand3_1 _7171_ (.B(_2179_),
    .C(_2254_),
    .A(net1853),
    .Y(_2787_));
 sg13g2_nand3_1 _7172_ (.B(_1879_),
    .C(_2323_),
    .A(net2045),
    .Y(_2788_));
 sg13g2_nand3_1 _7173_ (.B(net1934),
    .C(net1837),
    .A(net1889),
    .Y(_2789_));
 sg13g2_nand3_1 _7174_ (.B(_2788_),
    .C(_2789_),
    .A(_2787_),
    .Y(_2790_));
 sg13g2_o21ai_1 _7175_ (.B1(_2786_),
    .Y(_2791_),
    .A1(net2163),
    .A2(_2790_));
 sg13g2_a22oi_1 _7176_ (.Y(_2792_),
    .B1(_2791_),
    .B2(net1730),
    .A2(_2785_),
    .A1(net1743));
 sg13g2_nand2b_1 _7177_ (.Y(_2793_),
    .B(net2159),
    .A_N(_2792_));
 sg13g2_nand4_1 _7178_ (.B(net2191),
    .C(net1802),
    .A(net2174),
    .Y(_2794_),
    .D(_2750_));
 sg13g2_o21ai_1 _7179_ (.B1(net1887),
    .Y(_2795_),
    .A1(_1538_),
    .A2(net1854));
 sg13g2_o21ai_1 _7180_ (.B1(_2795_),
    .Y(_2796_),
    .A1(net1887),
    .A2(_1960_));
 sg13g2_nand2_1 _7181_ (.Y(_2797_),
    .A(_2794_),
    .B(_2796_));
 sg13g2_nand2_1 _7182_ (.Y(_2798_),
    .A(net1802),
    .B(_2451_));
 sg13g2_o21ai_1 _7183_ (.B1(_2798_),
    .Y(_2799_),
    .A1(net1930),
    .A2(_1699_));
 sg13g2_o21ai_1 _7184_ (.B1(net1993),
    .Y(_2800_),
    .A1(net2226),
    .A2(_1685_));
 sg13g2_a21oi_1 _7185_ (.A1(net1964),
    .A2(_2112_),
    .Y(_2801_),
    .B1(_2749_));
 sg13g2_a221oi_1 _7186_ (.B2(net2174),
    .C1(net2160),
    .B1(_2799_),
    .A1(net1802),
    .Y(_2802_),
    .A2(net1859));
 sg13g2_o21ai_1 _7187_ (.B1(_2802_),
    .Y(_2803_),
    .A1(_2800_),
    .A2(_2801_));
 sg13g2_a221oi_1 _7188_ (.B2(net2051),
    .C1(_2574_),
    .B1(_2803_),
    .A1(net1900),
    .Y(_2804_),
    .A2(_2797_));
 sg13g2_nand3_1 _7189_ (.B(net2141),
    .C(net1867),
    .A(net2042),
    .Y(_2805_));
 sg13g2_nand4_1 _7190_ (.B(_1513_),
    .C(_1796_),
    .A(net2197),
    .Y(_2806_),
    .D(_2048_));
 sg13g2_o21ai_1 _7191_ (.B1(_2806_),
    .Y(_2807_),
    .A1(_2629_),
    .A2(_2805_));
 sg13g2_a21oi_1 _7192_ (.A1(_1546_),
    .A2(_2089_),
    .Y(_2808_),
    .B1(_2566_));
 sg13g2_a221oi_1 _7193_ (.B2(net2049),
    .C1(_2808_),
    .B1(_2807_),
    .A1(net1880),
    .Y(_2809_),
    .A2(_2024_));
 sg13g2_nor2_1 _7194_ (.A(net1896),
    .B(_2809_),
    .Y(_2810_));
 sg13g2_a21oi_1 _7195_ (.A1(_1901_),
    .A2(_2156_),
    .Y(_2811_),
    .B1(_2730_));
 sg13g2_nand3_1 _7196_ (.B(net1849),
    .C(_1799_),
    .A(net1790),
    .Y(_2812_));
 sg13g2_nor2_1 _7197_ (.A(_1725_),
    .B(_2119_),
    .Y(_2813_));
 sg13g2_a21oi_1 _7198_ (.A1(_2812_),
    .A2(_2813_),
    .Y(_2814_),
    .B1(net1935));
 sg13g2_a21oi_1 _7199_ (.A1(_2368_),
    .A2(_2615_),
    .Y(_2815_),
    .B1(net2181));
 sg13g2_o21ai_1 _7200_ (.B1(net1910),
    .Y(_2816_),
    .A1(net2241),
    .A2(_2033_));
 sg13g2_o21ai_1 _7201_ (.B1(_2816_),
    .Y(_2817_),
    .A1(_1481_),
    .A2(_2811_));
 sg13g2_nor4_2 _7202_ (.A(net1940),
    .B(_2814_),
    .C(_2815_),
    .Y(_2818_),
    .D(_2817_));
 sg13g2_o21ai_1 _7203_ (.B1(_1747_),
    .Y(_2819_),
    .A1(_2810_),
    .A2(_2818_));
 sg13g2_a21o_1 _7204_ (.A2(net1958),
    .A1(net2247),
    .B1(_1931_),
    .X(_2820_));
 sg13g2_a21oi_1 _7205_ (.A1(net2220),
    .A2(_2820_),
    .Y(_2821_),
    .B1(_2704_));
 sg13g2_a221oi_1 _7206_ (.B2(_1778_),
    .C1(_2821_),
    .B1(net1928),
    .A1(net1913),
    .Y(_2822_),
    .A2(net1952));
 sg13g2_a21oi_1 _7207_ (.A1(_1912_),
    .A2(_1942_),
    .Y(_2823_),
    .B1(net1844));
 sg13g2_nor2_1 _7208_ (.A(net2196),
    .B(_2271_),
    .Y(_2824_));
 sg13g2_nor3_1 _7209_ (.A(net1930),
    .B(_1731_),
    .C(_1779_),
    .Y(_2825_));
 sg13g2_nor3_1 _7210_ (.A(_2823_),
    .B(_2824_),
    .C(_2825_),
    .Y(_2826_));
 sg13g2_o21ai_1 _7211_ (.B1(net1901),
    .Y(_2827_),
    .A1(net2179),
    .A2(_2826_));
 sg13g2_a21oi_1 _7212_ (.A1(net2179),
    .A2(_2822_),
    .Y(_2828_),
    .B1(_2827_));
 sg13g2_or2_1 _7213_ (.X(_2829_),
    .B(net1795),
    .A(net2044));
 sg13g2_nand2_1 _7214_ (.Y(_2830_),
    .A(_1984_),
    .B(_2829_));
 sg13g2_a22oi_1 _7215_ (.Y(_2831_),
    .B1(_2676_),
    .B2(net1967),
    .A2(_1653_),
    .A1(net2220));
 sg13g2_a221oi_1 _7216_ (.B2(_2049_),
    .C1(net2180),
    .B1(_2831_),
    .A1(_2778_),
    .Y(_2832_),
    .A2(_2830_));
 sg13g2_nand2_1 _7217_ (.Y(_2833_),
    .A(net1958),
    .B(_1610_));
 sg13g2_o21ai_1 _7218_ (.B1(net1962),
    .Y(_2834_),
    .A1(net2137),
    .A2(_2694_));
 sg13g2_a221oi_1 _7219_ (.B2(_2714_),
    .C1(net1936),
    .B1(_2834_),
    .A1(_2716_),
    .Y(_2835_),
    .A2(_2833_));
 sg13g2_o21ai_1 _7220_ (.B1(_1554_),
    .Y(_2836_),
    .A1(net2221),
    .A2(_2280_));
 sg13g2_o21ai_1 _7221_ (.B1(net1944),
    .Y(_2837_),
    .A1(net1905),
    .A2(_2836_));
 sg13g2_nor3_1 _7222_ (.A(_2832_),
    .B(_2835_),
    .C(_2837_),
    .Y(_2838_));
 sg13g2_nor3_1 _7223_ (.A(_1522_),
    .B(_1653_),
    .C(_1927_),
    .Y(_2839_));
 sg13g2_nor3_1 _7224_ (.A(_2828_),
    .B(_2838_),
    .C(_2839_),
    .Y(_2840_));
 sg13g2_nor2_1 _7225_ (.A(_1899_),
    .B(_2840_),
    .Y(_2841_));
 sg13g2_nor2_1 _7226_ (.A(net1945),
    .B(_2735_),
    .Y(_2842_));
 sg13g2_mux2_1 _7227_ (.A0(_2495_),
    .A1(net2189),
    .S(_2842_),
    .X(_2843_));
 sg13g2_a21oi_1 _7228_ (.A1(net2231),
    .A2(_1828_),
    .Y(_2844_),
    .B1(_2012_));
 sg13g2_nor2_1 _7229_ (.A(net2188),
    .B(_2730_),
    .Y(_2845_));
 sg13g2_a221oi_1 _7230_ (.B2(_2593_),
    .C1(_2729_),
    .B1(_2845_),
    .A1(net1928),
    .Y(_2846_),
    .A2(_2844_));
 sg13g2_nand3_1 _7231_ (.B(_1538_),
    .C(net1794),
    .A(net1983),
    .Y(_2847_));
 sg13g2_nand3_1 _7232_ (.B(net1834),
    .C(_2391_),
    .A(net1991),
    .Y(_2848_));
 sg13g2_o21ai_1 _7233_ (.B1(_2848_),
    .Y(_2849_),
    .A1(_1569_),
    .A2(_1643_));
 sg13g2_nand2b_1 _7234_ (.Y(_2850_),
    .B(_2847_),
    .A_N(_2849_));
 sg13g2_nand4_1 _7235_ (.B(_1796_),
    .C(_1880_),
    .A(net2042),
    .Y(_2851_),
    .D(_1912_));
 sg13g2_o21ai_1 _7236_ (.B1(_2851_),
    .Y(_2852_),
    .A1(net2215),
    .A2(_2824_));
 sg13g2_a21oi_1 _7237_ (.A1(net2194),
    .A2(net1837),
    .Y(_2853_),
    .B1(_1811_));
 sg13g2_a22oi_1 _7238_ (.Y(_2854_),
    .B1(_2852_),
    .B2(_2853_),
    .A2(_2850_),
    .A1(net1900));
 sg13g2_nor2b_1 _7239_ (.A(_2854_),
    .B_N(net1742),
    .Y(_2855_));
 sg13g2_a21oi_1 _7240_ (.A1(_1480_),
    .A2(net1885),
    .Y(_2856_),
    .B1(net1991));
 sg13g2_a22oi_1 _7241_ (.Y(_2857_),
    .B1(_1769_),
    .B2(net2031),
    .A2(_1583_),
    .A1(net1801));
 sg13g2_a21o_1 _7242_ (.A2(_2857_),
    .A1(net2040),
    .B1(_2856_),
    .X(_2858_));
 sg13g2_o21ai_1 _7243_ (.B1(_2858_),
    .Y(_2859_),
    .A1(net1797),
    .A2(_2026_));
 sg13g2_o21ai_1 _7244_ (.B1(_2340_),
    .Y(_2860_),
    .A1(_1585_),
    .A2(_2147_));
 sg13g2_a21oi_1 _7245_ (.A1(net2187),
    .A2(_2474_),
    .Y(_2861_),
    .B1(_1811_));
 sg13g2_a22oi_1 _7246_ (.Y(_2862_),
    .B1(_2860_),
    .B2(_2861_),
    .A2(_2859_),
    .A1(net1899));
 sg13g2_inv_1 _7247_ (.Y(_2863_),
    .A(_2862_));
 sg13g2_a21oi_1 _7248_ (.A1(_1790_),
    .A2(_2863_),
    .Y(_2864_),
    .B1(_2855_));
 sg13g2_nand3_1 _7249_ (.B(_1540_),
    .C(_2474_),
    .A(net1993),
    .Y(_2865_));
 sg13g2_a21oi_1 _7250_ (.A1(_1670_),
    .A2(net1834),
    .Y(_2866_),
    .B1(_2643_));
 sg13g2_a21oi_1 _7251_ (.A1(_2586_),
    .A2(_2750_),
    .Y(_2867_),
    .B1(_2866_));
 sg13g2_a21oi_1 _7252_ (.A1(_2865_),
    .A2(_2867_),
    .Y(_2868_),
    .B1(net1895));
 sg13g2_nand2_1 _7253_ (.Y(_2869_),
    .A(net1993),
    .B(_2254_));
 sg13g2_o21ai_1 _7254_ (.B1(net1859),
    .Y(_2870_),
    .A1(net2143),
    .A2(_1515_));
 sg13g2_a21oi_1 _7255_ (.A1(net2034),
    .A2(net1835),
    .Y(_2871_),
    .B1(_2870_));
 sg13g2_nor4_1 _7256_ (.A(net2160),
    .B(_1940_),
    .C(_2743_),
    .D(_2871_),
    .Y(_2872_));
 sg13g2_a21oi_1 _7257_ (.A1(_2869_),
    .A2(_2872_),
    .Y(_2873_),
    .B1(net2158));
 sg13g2_a21oi_1 _7258_ (.A1(net1814),
    .A2(net1835),
    .Y(_2874_),
    .B1(net1948));
 sg13g2_nor3_1 _7259_ (.A(_2868_),
    .B(_2873_),
    .C(_2874_),
    .Y(_2875_));
 sg13g2_nand2_1 _7260_ (.Y(_2876_),
    .A(_1862_),
    .B(_2290_));
 sg13g2_nand2_1 _7261_ (.Y(_2877_),
    .A(_2348_),
    .B(_2876_));
 sg13g2_a221oi_1 _7262_ (.B2(net2040),
    .C1(_2416_),
    .B1(_2877_),
    .A1(_1401_),
    .Y(_2878_),
    .A2(_1528_));
 sg13g2_o21ai_1 _7263_ (.B1(_1843_),
    .Y(_2879_),
    .A1(net2235),
    .A2(_2565_));
 sg13g2_mux2_1 _7264_ (.A0(_1889_),
    .A1(_2879_),
    .S(net2209),
    .X(_2880_));
 sg13g2_nor3_1 _7265_ (.A(net2173),
    .B(_1759_),
    .C(_2880_),
    .Y(_2881_));
 sg13g2_a21o_1 _7266_ (.A2(_2606_),
    .A1(_1580_),
    .B1(net1902),
    .X(_2882_));
 sg13g2_nor3_1 _7267_ (.A(net1885),
    .B(_1497_),
    .C(_1574_),
    .Y(_2883_));
 sg13g2_a21oi_1 _7268_ (.A1(net2207),
    .A2(_1723_),
    .Y(_2884_),
    .B1(_1615_));
 sg13g2_o21ai_1 _7269_ (.B1(net1901),
    .Y(_2885_),
    .A1(net1932),
    .A2(_2883_));
 sg13g2_a221oi_1 _7270_ (.B2(net1992),
    .C1(_2885_),
    .B1(_2884_),
    .A1(net1860),
    .Y(_2886_),
    .A2(_1685_));
 sg13g2_a21oi_1 _7271_ (.A1(_2882_),
    .A2(_2886_),
    .Y(_2887_),
    .B1(_2881_));
 sg13g2_o21ai_1 _7272_ (.B1(_2887_),
    .Y(_2888_),
    .A1(net1840),
    .A2(_2878_));
 sg13g2_o21ai_1 _7273_ (.B1(net2216),
    .Y(_2889_),
    .A1(net1958),
    .A2(_1651_));
 sg13g2_inv_1 _7274_ (.Y(_2890_),
    .A(_2889_));
 sg13g2_nand2_1 _7275_ (.Y(_2891_),
    .A(_1524_),
    .B(_2889_));
 sg13g2_nand2_1 _7276_ (.Y(_2892_),
    .A(net1955),
    .B(_1824_));
 sg13g2_a22oi_1 _7277_ (.Y(_2893_),
    .B1(net1985),
    .B2(_2102_),
    .A2(_0096_),
    .A1(net2205));
 sg13g2_nand2_1 _7278_ (.Y(_2894_),
    .A(_2892_),
    .B(_2893_));
 sg13g2_a22oi_1 _7279_ (.Y(_2895_),
    .B1(_2894_),
    .B2(net1855),
    .A2(_2891_),
    .A1(net1910));
 sg13g2_o21ai_1 _7280_ (.B1(_1480_),
    .Y(_2896_),
    .A1(_1704_),
    .A2(_2730_));
 sg13g2_nor3_1 _7281_ (.A(net2241),
    .B(_1516_),
    .C(_2565_),
    .Y(_2897_));
 sg13g2_o21ai_1 _7282_ (.B1(_1758_),
    .Y(_2898_),
    .A1(net1880),
    .A2(net1963));
 sg13g2_o21ai_1 _7283_ (.B1(net1840),
    .Y(_2899_),
    .A1(_2897_),
    .A2(_2898_));
 sg13g2_nand3_1 _7284_ (.B(_2896_),
    .C(_2899_),
    .A(_2895_),
    .Y(_2900_));
 sg13g2_a21oi_1 _7285_ (.A1(_1668_),
    .A2(_2875_),
    .Y(_2901_),
    .B1(net1732));
 sg13g2_nand3_1 _7286_ (.B(_2864_),
    .C(_2901_),
    .A(_2793_),
    .Y(_2902_));
 sg13g2_nor3_2 _7287_ (.A(_2773_),
    .B(_2804_),
    .C(_2902_),
    .Y(_2903_));
 sg13g2_a21oi_1 _7288_ (.A1(_1698_),
    .A2(_2888_),
    .Y(_2904_),
    .B1(_2841_));
 sg13g2_nor2_1 _7289_ (.A(net1894),
    .B(_2846_),
    .Y(_2905_));
 sg13g2_o21ai_1 _7290_ (.B1(_2905_),
    .Y(_2906_),
    .A1(net2172),
    .A2(_2843_));
 sg13g2_a21o_1 _7291_ (.A2(_2906_),
    .A1(_2900_),
    .B1(_1857_),
    .X(_2907_));
 sg13g2_nand4_1 _7292_ (.B(_2903_),
    .C(_2904_),
    .A(_2819_),
    .Y(_2908_),
    .D(_2907_));
 sg13g2_nor2_1 _7293_ (.A(net2045),
    .B(_2752_),
    .Y(_2909_));
 sg13g2_a221oi_1 _7294_ (.B2(_2751_),
    .C1(net2045),
    .B1(_2750_),
    .A1(net2038),
    .Y(_2910_),
    .A2(_1685_));
 sg13g2_o21ai_1 _7295_ (.B1(_3995_),
    .Y(_2911_),
    .A1(_2323_),
    .A2(_2525_));
 sg13g2_o21ai_1 _7296_ (.B1(_2747_),
    .Y(_2912_),
    .A1(_2910_),
    .A2(_2911_));
 sg13g2_o21ai_1 _7297_ (.B1(_2744_),
    .Y(_2913_),
    .A1(_2366_),
    .A2(_2800_));
 sg13g2_nand3_1 _7298_ (.B(_2912_),
    .C(_2913_),
    .A(net1732),
    .Y(_2914_));
 sg13g2_a21oi_1 _7299_ (.A1(_2908_),
    .A2(_2914_),
    .Y(_2915_),
    .B1(_2758_));
 sg13g2_nand2_1 _7300_ (.Y(_2916_),
    .A(\draw_game_inst.board_x[0] ),
    .B(\draw_game_inst.board_x[1] ));
 sg13g2_o21ai_1 _7301_ (.B1(net2197),
    .Y(_2917_),
    .A1(_2048_),
    .A2(_2565_));
 sg13g2_a21oi_1 _7302_ (.A1(_1754_),
    .A2(_2890_),
    .Y(_2918_),
    .B1(_2917_));
 sg13g2_nand2_1 _7303_ (.Y(_2919_),
    .A(_1654_),
    .B(_1730_));
 sg13g2_nand3_1 _7304_ (.B(net1811),
    .C(net1947),
    .A(net2241),
    .Y(_2920_));
 sg13g2_nand2_1 _7305_ (.Y(_2921_),
    .A(_2919_),
    .B(_2920_));
 sg13g2_inv_1 _7306_ (.Y(_2922_),
    .A(_2921_));
 sg13g2_and3_1 _7307_ (.X(_2923_),
    .A(net1985),
    .B(_1500_),
    .C(net1789));
 sg13g2_nand3_1 _7308_ (.B(_1592_),
    .C(net1842),
    .A(net1956),
    .Y(_2924_));
 sg13g2_o21ai_1 _7309_ (.B1(_2924_),
    .Y(_2925_),
    .A1(_1514_),
    .A2(_1594_));
 sg13g2_o21ai_1 _7310_ (.B1(net1794),
    .Y(_2926_),
    .A1(_2923_),
    .A2(_2925_));
 sg13g2_a221oi_1 _7311_ (.B2(net1928),
    .C1(_2918_),
    .B1(_2922_),
    .A1(net1913),
    .Y(_2927_),
    .A2(_2567_));
 sg13g2_o21ai_1 _7312_ (.B1(_2926_),
    .Y(_2928_),
    .A1(net2181),
    .A2(_2927_));
 sg13g2_and3_1 _7313_ (.X(_2929_),
    .A(net1813),
    .B(_1765_),
    .C(_2919_));
 sg13g2_a22oi_1 _7314_ (.Y(_2930_),
    .B1(net1811),
    .B2(net2024),
    .A2(_1399_),
    .A1(net2242));
 sg13g2_a21oi_1 _7315_ (.A1(net2035),
    .A2(_1635_),
    .Y(_2931_),
    .B1(net1856));
 sg13g2_a22oi_1 _7316_ (.Y(_2932_),
    .B1(_2774_),
    .B2(net1967),
    .A2(net1849),
    .A1(_1603_));
 sg13g2_a221oi_1 _7317_ (.B2(_2932_),
    .C1(_2929_),
    .B1(_2931_),
    .A1(_1732_),
    .Y(_2933_),
    .A2(_2930_));
 sg13g2_o21ai_1 _7318_ (.B1(_2933_),
    .Y(_2934_),
    .A1(_1662_),
    .A2(_1792_));
 sg13g2_a22oi_1 _7319_ (.Y(_2935_),
    .B1(_2934_),
    .B2(net1729),
    .A2(_2928_),
    .A1(net1742));
 sg13g2_nor2_1 _7320_ (.A(net1895),
    .B(_2935_),
    .Y(_2936_));
 sg13g2_nand2_1 _7321_ (.Y(_2937_),
    .A(_1909_),
    .B(_2533_));
 sg13g2_o21ai_1 _7322_ (.B1(net1994),
    .Y(_2938_),
    .A1(_1525_),
    .A2(_2937_));
 sg13g2_o21ai_1 _7323_ (.B1(net1953),
    .Y(_2939_),
    .A1(net2239),
    .A2(net2143));
 sg13g2_a221oi_1 _7324_ (.B2(_2939_),
    .C1(net2164),
    .B1(_1647_),
    .A1(net1909),
    .Y(_2940_),
    .A2(net1803));
 sg13g2_a21oi_2 _7325_ (.B1(_1709_),
    .Y(_2941_),
    .A2(net1812),
    .A1(net1882));
 sg13g2_a22oi_1 _7326_ (.Y(_2942_),
    .B1(_2575_),
    .B2(net2213),
    .A2(_2280_),
    .A1(_1935_));
 sg13g2_o21ai_1 _7327_ (.B1(_2940_),
    .Y(_2943_),
    .A1(_1630_),
    .A2(_2941_));
 sg13g2_o21ai_1 _7328_ (.B1(_2938_),
    .Y(_2944_),
    .A1(net1856),
    .A2(_2942_));
 sg13g2_or3_1 _7329_ (.A(_1656_),
    .B(_2044_),
    .C(_2045_),
    .X(_2945_));
 sg13g2_o21ai_1 _7330_ (.B1(_2945_),
    .Y(_2946_),
    .A1(_2943_),
    .A2(_2944_));
 sg13g2_nor2_1 _7331_ (.A(net2213),
    .B(_1610_),
    .Y(_2947_));
 sg13g2_nand2_1 _7332_ (.Y(_2948_),
    .A(net2033),
    .B(_1611_));
 sg13g2_a21oi_1 _7333_ (.A1(net2239),
    .A2(net1795),
    .Y(_2949_),
    .B1(_1929_));
 sg13g2_nor2_1 _7334_ (.A(net2213),
    .B(_2949_),
    .Y(_2950_));
 sg13g2_nor3_1 _7335_ (.A(net2044),
    .B(_1713_),
    .C(_2950_),
    .Y(_2951_));
 sg13g2_a21o_1 _7336_ (.A2(_2948_),
    .A1(_2263_),
    .B1(_2951_),
    .X(_2952_));
 sg13g2_a21oi_1 _7337_ (.A1(net2212),
    .A2(_1917_),
    .Y(_2953_),
    .B1(_1564_));
 sg13g2_a221oi_1 _7338_ (.B2(net1957),
    .C1(_2236_),
    .B1(net1872),
    .A1(net1988),
    .Y(_2954_),
    .A2(net1953));
 sg13g2_nor3_1 _7339_ (.A(net1840),
    .B(_2953_),
    .C(_2954_),
    .Y(_2955_));
 sg13g2_a221oi_1 _7340_ (.B2(_2636_),
    .C1(_2955_),
    .B1(_2952_),
    .A1(net2158),
    .Y(_2956_),
    .A2(_2946_));
 sg13g2_nand2b_1 _7341_ (.Y(_2957_),
    .B(net1743),
    .A_N(_2956_));
 sg13g2_nand2b_1 _7342_ (.Y(_2958_),
    .B(_1754_),
    .A_N(_2378_));
 sg13g2_o21ai_1 _7343_ (.B1(_2652_),
    .Y(_2959_),
    .A1(net2236),
    .A2(_1729_));
 sg13g2_nor2_1 _7344_ (.A(net1960),
    .B(_1702_),
    .Y(_2960_));
 sg13g2_a21oi_1 _7345_ (.A1(net1848),
    .A2(_1727_),
    .Y(_2961_),
    .B1(_2960_));
 sg13g2_o21ai_1 _7346_ (.B1(_2961_),
    .Y(_2962_),
    .A1(net2029),
    .A2(_1500_));
 sg13g2_a21oi_1 _7347_ (.A1(net2029),
    .A2(_2959_),
    .Y(_2963_),
    .B1(_2962_));
 sg13g2_o21ai_1 _7348_ (.B1(_2958_),
    .Y(_2964_),
    .A1(net2189),
    .A2(_2963_));
 sg13g2_a21oi_2 _7349_ (.B1(_1687_),
    .Y(_2965_),
    .A2(_1556_),
    .A1(net2236));
 sg13g2_nand2_1 _7350_ (.Y(_2966_),
    .A(net1846),
    .B(_2965_));
 sg13g2_nand2_1 _7351_ (.Y(_2967_),
    .A(_2964_),
    .B(_2966_));
 sg13g2_a221oi_1 _7352_ (.B2(net2218),
    .C1(net2042),
    .B1(_2699_),
    .A1(net1864),
    .Y(_2968_),
    .A2(_1715_));
 sg13g2_nand2_1 _7353_ (.Y(_2969_),
    .A(_1912_),
    .B(_2705_));
 sg13g2_a221oi_1 _7354_ (.B2(_1669_),
    .C1(_2968_),
    .B1(_2969_),
    .A1(net1913),
    .Y(_2970_),
    .A2(_2965_));
 sg13g2_a22oi_1 _7355_ (.Y(_2971_),
    .B1(_2970_),
    .B2(net1729),
    .A2(_2967_),
    .A1(net1742));
 sg13g2_o21ai_1 _7356_ (.B1(_2957_),
    .Y(_2972_),
    .A1(_1811_),
    .A2(_2971_));
 sg13g2_o21ai_1 _7357_ (.B1(net2174),
    .Y(_2973_),
    .A1(net2183),
    .A2(_2113_));
 sg13g2_o21ai_1 _7358_ (.B1(_2973_),
    .Y(_2974_),
    .A1(net2174),
    .A2(_1564_));
 sg13g2_nor3_1 _7359_ (.A(net2160),
    .B(_2380_),
    .C(_2974_),
    .Y(_2975_));
 sg13g2_nand2b_1 _7360_ (.Y(_2976_),
    .B(_2185_),
    .A_N(_1957_));
 sg13g2_nand3_1 _7361_ (.B(_1965_),
    .C(_2976_),
    .A(net1900),
    .Y(_2977_));
 sg13g2_o21ai_1 _7362_ (.B1(_2977_),
    .Y(_2978_),
    .A1(net2158),
    .A2(_2975_));
 sg13g2_o21ai_1 _7363_ (.B1(net2234),
    .Y(_2979_),
    .A1(net1996),
    .A2(net1809));
 sg13g2_nand3_1 _7364_ (.B(_1932_),
    .C(_2979_),
    .A(net2207),
    .Y(_2980_));
 sg13g2_nor2_1 _7365_ (.A(net2215),
    .B(_1558_),
    .Y(_2981_));
 sg13g2_a21oi_1 _7366_ (.A1(_1581_),
    .A2(_2981_),
    .Y(_2982_),
    .B1(net1934));
 sg13g2_a221oi_1 _7367_ (.B2(_2434_),
    .C1(net1904),
    .B1(_2045_),
    .A1(net1984),
    .Y(_2983_),
    .A2(_1873_));
 sg13g2_a21o_1 _7368_ (.A2(net1974),
    .A1(net2209),
    .B1(_1869_),
    .X(_2984_));
 sg13g2_a221oi_1 _7369_ (.B2(net1839),
    .C1(_2983_),
    .B1(_2984_),
    .A1(_2980_),
    .Y(_2985_),
    .A2(_2982_));
 sg13g2_nand3_1 _7370_ (.B(_2594_),
    .C(_2979_),
    .A(net1928),
    .Y(_2986_));
 sg13g2_a22oi_1 _7371_ (.Y(_2987_),
    .B1(_1577_),
    .B2(_1963_),
    .A2(net1867),
    .A1(net1892));
 sg13g2_a21oi_1 _7372_ (.A1(_1527_),
    .A2(_2987_),
    .Y(_2988_),
    .B1(net2047));
 sg13g2_o21ai_1 _7373_ (.B1(net1858),
    .Y(_2989_),
    .A1(net2204),
    .A2(_1754_));
 sg13g2_inv_1 _7374_ (.Y(_2990_),
    .A(_2989_));
 sg13g2_a21oi_1 _7375_ (.A1(net2130),
    .A2(net1955),
    .Y(_2991_),
    .B1(_1496_));
 sg13g2_a21oi_1 _7376_ (.A1(_1732_),
    .A2(_1754_),
    .Y(_2992_),
    .B1(net1894));
 sg13g2_o21ai_1 _7377_ (.B1(_2992_),
    .Y(_2993_),
    .A1(net1888),
    .A2(_2991_));
 sg13g2_a221oi_1 _7378_ (.B2(_1879_),
    .C1(_2993_),
    .B1(_2990_),
    .A1(_2986_),
    .Y(_2994_),
    .A2(_2988_));
 sg13g2_nor2_1 _7379_ (.A(_2985_),
    .B(_2994_),
    .Y(_2995_));
 sg13g2_nor2_1 _7380_ (.A(_1857_),
    .B(_2995_),
    .Y(_2996_));
 sg13g2_a221oi_1 _7381_ (.B2(net1993),
    .C1(net1853),
    .B1(_2070_),
    .A1(net2027),
    .Y(_2997_),
    .A2(_1537_));
 sg13g2_a21oi_1 _7382_ (.A1(_1525_),
    .A2(net1853),
    .Y(_2998_),
    .B1(_2997_));
 sg13g2_nand2_1 _7383_ (.Y(_2999_),
    .A(_1612_),
    .B(_2998_));
 sg13g2_a21o_1 _7384_ (.A2(_2948_),
    .A1(_1621_),
    .B1(net2192),
    .X(_3000_));
 sg13g2_a21oi_1 _7385_ (.A1(net1909),
    .A2(net1988),
    .Y(_3001_),
    .B1(_1623_));
 sg13g2_o21ai_1 _7386_ (.B1(_3001_),
    .Y(_3002_),
    .A1(net1906),
    .A2(_2472_));
 sg13g2_a221oi_1 _7387_ (.B2(_3002_),
    .C1(_1659_),
    .B1(net1790),
    .A1(_1393_),
    .Y(_3003_),
    .A2(net1799));
 sg13g2_o21ai_1 _7388_ (.B1(_3003_),
    .Y(_3004_),
    .A1(net2177),
    .A2(_3000_));
 sg13g2_a221oi_1 _7389_ (.B2(net2052),
    .C1(_1607_),
    .B1(_3004_),
    .A1(net1900),
    .Y(_3005_),
    .A2(_2999_));
 sg13g2_nor3_1 _7390_ (.A(net1732),
    .B(_2996_),
    .C(_3005_),
    .Y(_3006_));
 sg13g2_o21ai_1 _7391_ (.B1(_3006_),
    .Y(_3007_),
    .A1(_1954_),
    .A2(_2978_));
 sg13g2_nand2_1 _7392_ (.Y(_3008_),
    .A(net1962),
    .B(net1795));
 sg13g2_a21oi_1 _7393_ (.A1(_1909_),
    .A2(_3008_),
    .Y(_3009_),
    .B1(net2195));
 sg13g2_a221oi_1 _7394_ (.B2(net1850),
    .C1(_3009_),
    .B1(_1933_),
    .A1(net1845),
    .Y(_3010_),
    .A2(net1787));
 sg13g2_a21oi_1 _7395_ (.A1(_1647_),
    .A2(net1795),
    .Y(_3011_),
    .B1(_1946_));
 sg13g2_o21ai_1 _7396_ (.B1(_3011_),
    .Y(_3012_),
    .A1(net2176),
    .A2(_3010_));
 sg13g2_nand2_1 _7397_ (.Y(_3013_),
    .A(net1900),
    .B(_3012_));
 sg13g2_nor4_1 _7398_ (.A(net2195),
    .B(_1918_),
    .C(_1943_),
    .D(_2534_),
    .Y(_3014_));
 sg13g2_a21oi_1 _7399_ (.A1(net1844),
    .A2(_2829_),
    .Y(_3015_),
    .B1(_2950_));
 sg13g2_nor2_1 _7400_ (.A(_3014_),
    .B(_3015_),
    .Y(_3016_));
 sg13g2_a22oi_1 _7401_ (.Y(_3017_),
    .B1(_2290_),
    .B2(_2432_),
    .A2(net1788),
    .A1(net2210));
 sg13g2_a21oi_1 _7402_ (.A1(_1400_),
    .A2(net1807),
    .Y(_3018_),
    .B1(_1984_));
 sg13g2_o21ai_1 _7403_ (.B1(_1631_),
    .Y(_3019_),
    .A1(net1812),
    .A2(net1973));
 sg13g2_a21oi_1 _7404_ (.A1(net2178),
    .A2(_3018_),
    .Y(_3020_),
    .B1(net2160));
 sg13g2_nand2_1 _7405_ (.Y(_3021_),
    .A(_3019_),
    .B(_3020_));
 sg13g2_a221oi_1 _7406_ (.B2(net1909),
    .C1(_3021_),
    .B1(_3017_),
    .A1(net2048),
    .Y(_3022_),
    .A2(_3016_));
 sg13g2_o21ai_1 _7407_ (.B1(_3013_),
    .Y(_3023_),
    .A1(net1948),
    .A2(_1924_));
 sg13g2_nor2_1 _7408_ (.A(_1899_),
    .B(_3023_),
    .Y(_3024_));
 sg13g2_o21ai_1 _7409_ (.B1(_3024_),
    .Y(_3025_),
    .A1(net2159),
    .A2(_3022_));
 sg13g2_o21ai_1 _7410_ (.B1(_2644_),
    .Y(_3026_),
    .A1(_1759_),
    .A2(_2108_));
 sg13g2_a21oi_1 _7411_ (.A1(net2041),
    .A2(net2198),
    .Y(_3027_),
    .B1(net2168));
 sg13g2_nand2_1 _7412_ (.Y(_3028_),
    .A(net1865),
    .B(_3027_));
 sg13g2_nor3_1 _7413_ (.A(net1938),
    .B(_1993_),
    .C(_3028_),
    .Y(_3029_));
 sg13g2_nor3_1 _7414_ (.A(net2225),
    .B(net2038),
    .C(net2198),
    .Y(_3030_));
 sg13g2_a22oi_1 _7415_ (.Y(_3031_),
    .B1(_3030_),
    .B2(_1863_),
    .A2(_1963_),
    .A1(net1873));
 sg13g2_nor2_1 _7416_ (.A(_2644_),
    .B(_3031_),
    .Y(_3032_));
 sg13g2_a21o_1 _7417_ (.A2(_3026_),
    .A1(net2168),
    .B1(_3032_),
    .X(_3033_));
 sg13g2_o21ai_1 _7418_ (.B1(_1668_),
    .Y(_3034_),
    .A1(_3029_),
    .A2(_3033_));
 sg13g2_o21ai_1 _7419_ (.B1(_2979_),
    .Y(_3035_),
    .A1(net2234),
    .A2(_1890_));
 sg13g2_a21oi_1 _7420_ (.A1(net2208),
    .A2(_3035_),
    .Y(_3036_),
    .B1(_1759_));
 sg13g2_o21ai_1 _7421_ (.B1(_3036_),
    .Y(_3037_),
    .A1(net1801),
    .A2(_1716_));
 sg13g2_a221oi_1 _7422_ (.B2(_3998_),
    .C1(net1932),
    .B1(_1753_),
    .A1(_1401_),
    .Y(_3038_),
    .A2(_1651_));
 sg13g2_or2_1 _7423_ (.X(_3039_),
    .B(_3038_),
    .A(_2088_));
 sg13g2_a21oi_1 _7424_ (.A1(net1892),
    .A2(net1812),
    .Y(_3040_),
    .B1(_2025_));
 sg13g2_a221oi_1 _7425_ (.B2(_1499_),
    .C1(_3040_),
    .B1(_3039_),
    .A1(net1839),
    .Y(_3041_),
    .A2(_3037_));
 sg13g2_a21o_1 _7426_ (.A2(_2112_),
    .A1(net1994),
    .B1(_2630_),
    .X(_3042_));
 sg13g2_a221oi_1 _7427_ (.B2(_1684_),
    .C1(_2627_),
    .B1(_3042_),
    .A1(_2173_),
    .Y(_3043_),
    .A2(_2439_));
 sg13g2_o21ai_1 _7428_ (.B1(_1747_),
    .Y(_3044_),
    .A1(_3041_),
    .A2(_3043_));
 sg13g2_a21oi_1 _7429_ (.A1(net2235),
    .A2(_1891_),
    .Y(_3045_),
    .B1(_1721_));
 sg13g2_nor2_1 _7430_ (.A(_1483_),
    .B(_3045_),
    .Y(_3046_));
 sg13g2_a21oi_1 _7431_ (.A1(net2234),
    .A2(net1838),
    .Y(_3047_),
    .B1(_1892_));
 sg13g2_nand3_1 _7432_ (.B(net1870),
    .C(_1545_),
    .A(net1882),
    .Y(_3048_));
 sg13g2_o21ai_1 _7433_ (.B1(_3048_),
    .Y(_3049_),
    .A1(net1876),
    .A2(_2025_));
 sg13g2_nand3_1 _7434_ (.B(net1858),
    .C(net1837),
    .A(_1544_),
    .Y(_3050_));
 sg13g2_o21ai_1 _7435_ (.B1(_3050_),
    .Y(_3051_),
    .A1(_1733_),
    .A2(_3047_));
 sg13g2_nor4_1 _7436_ (.A(_2609_),
    .B(_3046_),
    .C(_3049_),
    .D(_3051_),
    .Y(_3052_));
 sg13g2_nand2_1 _7437_ (.Y(_3053_),
    .A(net1847),
    .B(_2665_));
 sg13g2_a21oi_1 _7438_ (.A1(_2601_),
    .A2(_3053_),
    .Y(_3054_),
    .B1(net2173));
 sg13g2_a221oi_1 _7439_ (.B2(net2205),
    .C1(_1496_),
    .B1(net1838),
    .A1(net2130),
    .Y(_3055_),
    .A2(net1955));
 sg13g2_o21ai_1 _7440_ (.B1(net1852),
    .Y(_3056_),
    .A1(net2208),
    .A2(net1837));
 sg13g2_a21oi_1 _7441_ (.A1(net2208),
    .A2(net1976),
    .Y(_3057_),
    .B1(_3056_));
 sg13g2_a21oi_1 _7442_ (.A1(_2275_),
    .A2(_2512_),
    .Y(_3058_),
    .B1(_1481_));
 sg13g2_o21ai_1 _7443_ (.B1(net1942),
    .Y(_3059_),
    .A1(net1902),
    .A2(_3055_));
 sg13g2_nor4_1 _7444_ (.A(_3054_),
    .B(_3057_),
    .C(_3058_),
    .D(_3059_),
    .Y(_3060_));
 sg13g2_o21ai_1 _7445_ (.B1(_1698_),
    .Y(_3061_),
    .A1(_3052_),
    .A2(_3060_));
 sg13g2_nand4_1 _7446_ (.B(_3034_),
    .C(_3044_),
    .A(_3025_),
    .Y(_3062_),
    .D(_3061_));
 sg13g2_or4_2 _7447_ (.A(_2936_),
    .B(_2972_),
    .C(_3007_),
    .D(_3062_),
    .X(_3063_));
 sg13g2_nand4_1 _7448_ (.B(net1929),
    .C(_2587_),
    .A(_1563_),
    .Y(_3064_),
    .D(_2636_));
 sg13g2_nand2b_1 _7449_ (.Y(_3065_),
    .B(_2909_),
    .A_N(_2450_));
 sg13g2_nand2b_1 _7450_ (.Y(_3066_),
    .B(_2526_),
    .A_N(_2128_));
 sg13g2_nand2_1 _7451_ (.Y(_3067_),
    .A(_3065_),
    .B(_3066_));
 sg13g2_o21ai_1 _7452_ (.B1(_2747_),
    .Y(_3068_),
    .A1(net2162),
    .A2(_3067_));
 sg13g2_nand3_1 _7453_ (.B(_3064_),
    .C(_3068_),
    .A(net1731),
    .Y(_3069_));
 sg13g2_a21oi_1 _7454_ (.A1(_3063_),
    .A2(_3069_),
    .Y(_3070_),
    .B1(_2916_));
 sg13g2_o21ai_1 _7455_ (.B1(_3000_),
    .Y(_3071_),
    .A1(_1527_),
    .A2(net1953));
 sg13g2_a21oi_1 _7456_ (.A1(net1969),
    .A2(net1953),
    .Y(_3072_),
    .B1(net2175));
 sg13g2_nor3_1 _7457_ (.A(net1939),
    .B(_2683_),
    .C(_2751_),
    .Y(_3073_));
 sg13g2_nor2_1 _7458_ (.A(_2636_),
    .B(_3073_),
    .Y(_3074_));
 sg13g2_a221oi_1 _7459_ (.B2(_3072_),
    .C1(_3074_),
    .B1(_3071_),
    .A1(_1642_),
    .Y(_3075_),
    .A2(_2000_));
 sg13g2_nor3_1 _7460_ (.A(_1913_),
    .B(_1927_),
    .C(_2247_),
    .Y(_3076_));
 sg13g2_nor3_1 _7461_ (.A(net2192),
    .B(_1525_),
    .C(_2688_),
    .Y(_3077_));
 sg13g2_nor2_1 _7462_ (.A(_1641_),
    .B(net1787),
    .Y(_3078_));
 sg13g2_nor4_1 _7463_ (.A(net2175),
    .B(_2195_),
    .C(_3077_),
    .D(_3078_),
    .Y(_3079_));
 sg13g2_a21oi_1 _7464_ (.A1(_2273_),
    .A2(_2947_),
    .Y(_3080_),
    .B1(_2014_));
 sg13g2_and2_1 _7465_ (.A(net1853),
    .B(_3080_),
    .X(_3081_));
 sg13g2_a22oi_1 _7466_ (.Y(_3082_),
    .B1(_2271_),
    .B2(net1969),
    .A2(_1547_),
    .A1(_1546_));
 sg13g2_nor4_1 _7467_ (.A(net1895),
    .B(_3079_),
    .C(_3081_),
    .D(_3082_),
    .Y(_3083_));
 sg13g2_nor3_1 _7468_ (.A(_3075_),
    .B(_3076_),
    .C(_3083_),
    .Y(_3084_));
 sg13g2_nor2b_2 _7469_ (.A(_3084_),
    .B_N(net1743),
    .Y(_3085_));
 sg13g2_o21ai_1 _7470_ (.B1(_3008_),
    .Y(_3086_),
    .A1(net2036),
    .A2(_1803_));
 sg13g2_a221oi_1 _7471_ (.B2(net1910),
    .C1(net2164),
    .B1(_2217_),
    .A1(net1913),
    .Y(_3087_),
    .A2(net1795));
 sg13g2_a22oi_1 _7472_ (.Y(_3088_),
    .B1(_3086_),
    .B2(net1859),
    .A2(_1999_),
    .A1(net1813));
 sg13g2_a21oi_1 _7473_ (.A1(_1944_),
    .A2(_3008_),
    .Y(_3089_),
    .B1(net1936));
 sg13g2_nand3b_1 _7474_ (.B(_3088_),
    .C(_3087_),
    .Y(_3090_),
    .A_N(_3089_));
 sg13g2_o21ai_1 _7475_ (.B1(_3090_),
    .Y(_3091_),
    .A1(_1512_),
    .A2(_2044_));
 sg13g2_nor3_1 _7476_ (.A(net2195),
    .B(_1918_),
    .C(_2719_),
    .Y(_3092_));
 sg13g2_nand2_1 _7477_ (.Y(_3093_),
    .A(net2049),
    .B(_2829_));
 sg13g2_nor2_1 _7478_ (.A(_3092_),
    .B(_3093_),
    .Y(_3094_));
 sg13g2_a21oi_1 _7479_ (.A1(net1808),
    .A2(net1962),
    .Y(_3095_),
    .B1(net1935));
 sg13g2_o21ai_1 _7480_ (.B1(_3095_),
    .Y(_3096_),
    .A1(net1962),
    .A2(_1999_));
 sg13g2_nor2_1 _7481_ (.A(net1905),
    .B(_2508_),
    .Y(_3097_));
 sg13g2_o21ai_1 _7482_ (.B1(net1944),
    .Y(_3098_),
    .A1(_1394_),
    .A2(_1596_));
 sg13g2_nor3_1 _7483_ (.A(_3094_),
    .B(_3097_),
    .C(_3098_),
    .Y(_3099_));
 sg13g2_a22oi_1 _7484_ (.Y(_3100_),
    .B1(_3096_),
    .B2(_3099_),
    .A2(_3091_),
    .A1(net2159));
 sg13g2_nor2_2 _7485_ (.A(_1899_),
    .B(_3100_),
    .Y(_3101_));
 sg13g2_a21oi_1 _7486_ (.A1(net2201),
    .A2(_2185_),
    .Y(_3102_),
    .B1(net2046));
 sg13g2_a21oi_1 _7487_ (.A1(net2045),
    .A2(_2740_),
    .Y(_3103_),
    .B1(_3102_));
 sg13g2_nor3_1 _7488_ (.A(net2041),
    .B(_1533_),
    .C(_3103_),
    .Y(_3104_));
 sg13g2_nor4_1 _7489_ (.A(net2160),
    .B(_2148_),
    .C(_2588_),
    .D(_3104_),
    .Y(_3105_));
 sg13g2_nor3_1 _7490_ (.A(net2046),
    .B(_2147_),
    .C(_2584_),
    .Y(_3106_));
 sg13g2_o21ai_1 _7491_ (.B1(_3106_),
    .Y(_3107_),
    .A1(net1844),
    .A2(_2061_));
 sg13g2_o21ai_1 _7492_ (.B1(_1977_),
    .Y(_3108_),
    .A1(net1969),
    .A2(net1864));
 sg13g2_a21oi_1 _7493_ (.A1(_2255_),
    .A2(_3108_),
    .Y(_3109_),
    .B1(net1895));
 sg13g2_a21oi_1 _7494_ (.A1(_3107_),
    .A2(_3109_),
    .Y(_3110_),
    .B1(_1954_));
 sg13g2_o21ai_1 _7495_ (.B1(_3110_),
    .Y(_3111_),
    .A1(net2158),
    .A2(_3105_));
 sg13g2_a22oi_1 _7496_ (.Y(_3112_),
    .B1(net1847),
    .B2(net1797),
    .A2(net2145),
    .A1(net2029));
 sg13g2_nand3_1 _7497_ (.B(_1799_),
    .C(_1964_),
    .A(_1625_),
    .Y(_3113_));
 sg13g2_o21ai_1 _7498_ (.B1(_1810_),
    .Y(_3114_),
    .A1(net2188),
    .A2(_3112_));
 sg13g2_nand2b_1 _7499_ (.Y(_3115_),
    .B(_3113_),
    .A_N(_3114_));
 sg13g2_nand3_1 _7500_ (.B(_1592_),
    .C(net1842),
    .A(net1981),
    .Y(_3116_));
 sg13g2_o21ai_1 _7501_ (.B1(_3116_),
    .Y(_3117_),
    .A1(net1981),
    .A2(net1797));
 sg13g2_nor2_1 _7502_ (.A(_1516_),
    .B(_1753_),
    .Y(_3118_));
 sg13g2_nand2_1 _7503_ (.Y(_3119_),
    .A(net2216),
    .B(_2921_));
 sg13g2_a21oi_1 _7504_ (.A1(_1523_),
    .A2(_1730_),
    .Y(_3120_),
    .B1(net2197));
 sg13g2_nand3_1 _7505_ (.B(net1790),
    .C(_1799_),
    .A(net1988),
    .Y(_3121_));
 sg13g2_nand3_1 _7506_ (.B(_3120_),
    .C(_3121_),
    .A(_3119_),
    .Y(_3122_));
 sg13g2_o21ai_1 _7507_ (.B1(_3122_),
    .Y(_3123_),
    .A1(_2917_),
    .A2(_3118_));
 sg13g2_a22oi_1 _7508_ (.Y(_3124_),
    .B1(_3123_),
    .B2(net2047),
    .A2(_3117_),
    .A1(net1794));
 sg13g2_o21ai_1 _7509_ (.B1(_3115_),
    .Y(_3125_),
    .A1(net1894),
    .A2(_3124_));
 sg13g2_nand2_1 _7510_ (.Y(_3126_),
    .A(net1742),
    .B(_3125_));
 sg13g2_nand2_1 _7511_ (.Y(_3127_),
    .A(_1527_),
    .B(net1871));
 sg13g2_a21oi_1 _7512_ (.A1(_2645_),
    .A2(_3127_),
    .Y(_3128_),
    .B1(_2644_));
 sg13g2_a21oi_1 _7513_ (.A1(net2038),
    .A2(_2394_),
    .Y(_3129_),
    .B1(net2046));
 sg13g2_a221oi_1 _7514_ (.B2(net2038),
    .C1(net2045),
    .B1(_2394_),
    .A1(net2228),
    .Y(_3130_),
    .A2(_2195_));
 sg13g2_nor3_1 _7515_ (.A(net1938),
    .B(_2748_),
    .C(_3130_),
    .Y(_3131_));
 sg13g2_o21ai_1 _7516_ (.B1(_1668_),
    .Y(_3132_),
    .A1(_3128_),
    .A2(_3131_));
 sg13g2_a221oi_1 _7517_ (.B2(_1797_),
    .C1(_2308_),
    .B1(net1849),
    .A1(net2035),
    .Y(_3133_),
    .A2(net2145));
 sg13g2_nor2b_1 _7518_ (.A(_2451_),
    .B_N(_1847_),
    .Y(_3134_));
 sg13g2_nor3_1 _7519_ (.A(_1811_),
    .B(_3018_),
    .C(_3134_),
    .Y(_3135_));
 sg13g2_o21ai_1 _7520_ (.B1(_3135_),
    .Y(_3136_),
    .A1(net2197),
    .A2(_3133_));
 sg13g2_a21oi_1 _7521_ (.A1(_1559_),
    .A2(_1878_),
    .Y(_3137_),
    .B1(net1809));
 sg13g2_a221oi_1 _7522_ (.B2(net2207),
    .C1(net2173),
    .B1(_3137_),
    .A1(net1986),
    .Y(_3138_),
    .A2(_1847_));
 sg13g2_nor2_1 _7523_ (.A(_1727_),
    .B(_2662_),
    .Y(_3139_));
 sg13g2_a22oi_1 _7524_ (.Y(_3140_),
    .B1(_3139_),
    .B2(_1509_),
    .A2(_1832_),
    .A1(net1985));
 sg13g2_nor2_1 _7525_ (.A(net1903),
    .B(_3140_),
    .Y(_3141_));
 sg13g2_a221oi_1 _7526_ (.B2(_3138_),
    .C1(_3141_),
    .B1(_3120_),
    .A1(_1621_),
    .Y(_3142_),
    .A2(_2931_));
 sg13g2_o21ai_1 _7527_ (.B1(_3136_),
    .Y(_3143_),
    .A1(net1895),
    .A2(_3142_));
 sg13g2_o21ai_1 _7528_ (.B1(_1699_),
    .Y(_3144_),
    .A1(net1880),
    .A2(_1722_));
 sg13g2_o21ai_1 _7529_ (.B1(_2630_),
    .Y(_3145_),
    .A1(net2214),
    .A2(_3144_));
 sg13g2_nand2_1 _7530_ (.Y(_3146_),
    .A(net2027),
    .B(_1691_));
 sg13g2_a221oi_1 _7531_ (.B2(net2048),
    .C1(_2627_),
    .B1(_3146_),
    .A1(net1798),
    .Y(_3147_),
    .A2(_2483_));
 sg13g2_nand2_1 _7532_ (.Y(_3148_),
    .A(_3145_),
    .B(_3147_));
 sg13g2_o21ai_1 _7533_ (.B1(net1942),
    .Y(_3149_),
    .A1(_1546_),
    .A2(_1890_));
 sg13g2_a22oi_1 _7534_ (.Y(_3150_),
    .B1(_1901_),
    .B2(_1725_),
    .A2(_1891_),
    .A1(net2216));
 sg13g2_a21oi_1 _7535_ (.A1(_2512_),
    .A2(_2599_),
    .Y(_3151_),
    .B1(_1481_));
 sg13g2_nor3_1 _7536_ (.A(_3040_),
    .B(_3149_),
    .C(_3151_),
    .Y(_3152_));
 sg13g2_o21ai_1 _7537_ (.B1(_3152_),
    .Y(_3153_),
    .A1(net1935),
    .A2(_3150_));
 sg13g2_o21ai_1 _7538_ (.B1(_3148_),
    .Y(_3154_),
    .A1(_2617_),
    .A2(_3153_));
 sg13g2_nand2_1 _7539_ (.Y(_3155_),
    .A(_1747_),
    .B(_3154_));
 sg13g2_o21ai_1 _7540_ (.B1(net1893),
    .Y(_3156_),
    .A1(_1859_),
    .A2(_1925_));
 sg13g2_a22oi_1 _7541_ (.Y(_3157_),
    .B1(_1723_),
    .B2(net1927),
    .A2(_1675_),
    .A1(net1887));
 sg13g2_nand3_1 _7542_ (.B(net1788),
    .C(_1966_),
    .A(_1519_),
    .Y(_3158_));
 sg13g2_a21oi_1 _7543_ (.A1(_3129_),
    .A2(_3158_),
    .Y(_3159_),
    .B1(_3157_));
 sg13g2_o21ai_1 _7544_ (.B1(_3156_),
    .Y(_3160_),
    .A1(net2165),
    .A2(_3159_));
 sg13g2_a221oi_1 _7545_ (.B2(_1528_),
    .C1(_2416_),
    .B1(_1701_),
    .A1(net1801),
    .Y(_3161_),
    .A2(net1927));
 sg13g2_nor2_1 _7546_ (.A(net1840),
    .B(_3161_),
    .Y(_3162_));
 sg13g2_o21ai_1 _7547_ (.B1(net1845),
    .Y(_3163_),
    .A1(_1522_),
    .A2(_1604_));
 sg13g2_nand3_1 _7548_ (.B(_3000_),
    .C(_3163_),
    .A(_2636_),
    .Y(_3164_));
 sg13g2_o21ai_1 _7549_ (.B1(_3160_),
    .Y(_3165_),
    .A1(_2355_),
    .A2(_3164_));
 sg13g2_o21ai_1 _7550_ (.B1(net1730),
    .Y(_3166_),
    .A1(_3162_),
    .A2(_3165_));
 sg13g2_a221oi_1 _7551_ (.B2(net1812),
    .C1(net2030),
    .B1(_1709_),
    .A1(net2232),
    .Y(_3167_),
    .A2(net1947));
 sg13g2_o21ai_1 _7552_ (.B1(net1907),
    .Y(_3168_),
    .A1(_1496_),
    .A2(_3167_));
 sg13g2_o21ai_1 _7553_ (.B1(net1851),
    .Y(_3169_),
    .A1(_1878_),
    .A2(_1936_));
 sg13g2_o21ai_1 _7554_ (.B1(_2211_),
    .Y(_3170_),
    .A1(net2232),
    .A2(_1753_));
 sg13g2_a22oi_1 _7555_ (.Y(_3171_),
    .B1(net1848),
    .B2(net2130),
    .A2(net1960),
    .A1(net1974));
 sg13g2_o21ai_1 _7556_ (.B1(_3171_),
    .Y(_3172_),
    .A1(net1960),
    .A2(_1753_));
 sg13g2_a22oi_1 _7557_ (.Y(_3173_),
    .B1(_3172_),
    .B2(net1991),
    .A2(_3170_),
    .A1(_2990_));
 sg13g2_nand4_1 _7558_ (.B(_3168_),
    .C(_3169_),
    .A(net1899),
    .Y(_3174_),
    .D(_3173_));
 sg13g2_a21oi_1 _7559_ (.A1(net2204),
    .A2(_1830_),
    .Y(_3175_),
    .B1(net2184));
 sg13g2_or2_1 _7560_ (.X(_3176_),
    .B(_3175_),
    .A(net2172));
 sg13g2_o21ai_1 _7561_ (.B1(net2241),
    .Y(_3177_),
    .A1(_1570_),
    .A2(_1737_));
 sg13g2_a21oi_2 _7562_ (.B1(_1481_),
    .Y(_3178_),
    .A2(_3177_),
    .A1(_1722_));
 sg13g2_o21ai_1 _7563_ (.B1(_3178_),
    .Y(_3179_),
    .A1(net2134),
    .A2(_1652_));
 sg13g2_a22oi_1 _7564_ (.Y(_3180_),
    .B1(_1653_),
    .B2(net1863),
    .A2(_1558_),
    .A1(net1870));
 sg13g2_nand2b_1 _7565_ (.Y(_3181_),
    .B(_2493_),
    .A_N(net2232));
 sg13g2_a221oi_1 _7566_ (.B2(_2211_),
    .C1(net1932),
    .B1(_3181_),
    .A1(net2030),
    .Y(_3182_),
    .A2(_3180_));
 sg13g2_nor2_1 _7567_ (.A(_1506_),
    .B(_1546_),
    .Y(_3183_));
 sg13g2_a21oi_1 _7568_ (.A1(_1700_),
    .A2(net1833),
    .Y(_3184_),
    .B1(_2025_));
 sg13g2_nor4_1 _7569_ (.A(net1940),
    .B(_3182_),
    .C(_3183_),
    .D(_3184_),
    .Y(_3185_));
 sg13g2_nand3_1 _7570_ (.B(_3179_),
    .C(_3185_),
    .A(_3176_),
    .Y(_3186_));
 sg13g2_a21oi_2 _7571_ (.B1(_1857_),
    .Y(_3187_),
    .A2(_3186_),
    .A1(_3174_));
 sg13g2_a21oi_1 _7572_ (.A1(_1559_),
    .A2(_2593_),
    .Y(_3188_),
    .B1(_3056_));
 sg13g2_o21ai_1 _7573_ (.B1(net1943),
    .Y(_3189_),
    .A1(net1903),
    .A2(net1876));
 sg13g2_nor4_1 _7574_ (.A(_3054_),
    .B(_3178_),
    .C(_3188_),
    .D(_3189_),
    .Y(_3190_));
 sg13g2_a22oi_1 _7575_ (.Y(_3191_),
    .B1(_2493_),
    .B2(_1545_),
    .A2(net1794),
    .A1(net1975));
 sg13g2_a22oi_1 _7576_ (.Y(_3192_),
    .B1(_1891_),
    .B2(_1732_),
    .A2(net1837),
    .A1(net1858));
 sg13g2_nand2_1 _7577_ (.Y(_3193_),
    .A(_3191_),
    .B(_3192_));
 sg13g2_nor3_1 _7578_ (.A(_2609_),
    .B(_3046_),
    .C(_3193_),
    .Y(_3194_));
 sg13g2_o21ai_1 _7579_ (.B1(_1698_),
    .Y(_3195_),
    .A1(_3190_),
    .A2(_3194_));
 sg13g2_a21oi_1 _7580_ (.A1(net1729),
    .A2(_3143_),
    .Y(_3196_),
    .B1(net1732));
 sg13g2_nand3_1 _7581_ (.B(_3166_),
    .C(_3196_),
    .A(_3155_),
    .Y(_3197_));
 sg13g2_nor4_2 _7582_ (.A(_3085_),
    .B(_3101_),
    .C(_3187_),
    .Y(_3198_),
    .D(_3197_));
 sg13g2_and4_1 _7583_ (.A(_3111_),
    .B(_3126_),
    .C(_3132_),
    .D(_3195_),
    .X(_3199_));
 sg13g2_a221oi_1 _7584_ (.B2(net1854),
    .C1(net1938),
    .B1(_2474_),
    .A1(net1802),
    .Y(_3200_),
    .A2(_1623_));
 sg13g2_a221oi_1 _7585_ (.B2(net1907),
    .C1(_2588_),
    .B1(_2581_),
    .A1(net1798),
    .Y(_3201_),
    .A2(_2575_));
 sg13g2_a21oi_1 _7586_ (.A1(_2236_),
    .A2(_2909_),
    .Y(_3202_),
    .B1(net2162));
 sg13g2_nand2_1 _7587_ (.Y(_3203_),
    .A(_3028_),
    .B(_3202_));
 sg13g2_a22oi_1 _7588_ (.Y(_3204_),
    .B1(_3203_),
    .B2(_2747_),
    .A2(_3201_),
    .A1(_3200_));
 sg13g2_a22oi_1 _7589_ (.Y(_3205_),
    .B1(_3204_),
    .B2(net1732),
    .A2(_3199_),
    .A1(_3198_));
 sg13g2_nor2_1 _7590_ (.A(_2507_),
    .B(_3205_),
    .Y(_3206_));
 sg13g2_o21ai_1 _7591_ (.B1(\draw_game_inst.board_x[2] ),
    .Y(_3207_),
    .A1(_2400_),
    .A2(_2556_));
 sg13g2_nor4_1 _7592_ (.A(_2757_),
    .B(_2915_),
    .C(_3070_),
    .D(_3206_),
    .Y(_3208_));
 sg13g2_o21ai_1 _7593_ (.B1(_1478_),
    .Y(_3209_),
    .A1(\draw_game_inst.board_x[2] ),
    .A2(_3208_));
 sg13g2_nand2b_2 _7594_ (.Y(_3210_),
    .B(_3207_),
    .A_N(_3209_));
 sg13g2_and2_1 _7595_ (.A(_1424_),
    .B(_3210_),
    .X(_3211_));
 sg13g2_inv_1 _7596_ (.Y(_3212_),
    .A(_3211_));
 sg13g2_a21oi_2 _7597_ (.B1(_3959_),
    .Y(_3213_),
    .A2(net5),
    .A1(net6));
 sg13g2_nor2_1 _7598_ (.A(net1949),
    .B(_1632_),
    .Y(_3214_));
 sg13g2_nand3_1 _7599_ (.B(net995),
    .C(net829),
    .A(net998),
    .Y(_3215_));
 sg13g2_or2_2 _7600_ (.X(_3216_),
    .B(_3215_),
    .A(net2028));
 sg13g2_nor2_2 _7601_ (.A(_1402_),
    .B(_3216_),
    .Y(_3217_));
 sg13g2_nor3_1 _7602_ (.A(\draw_game_inst.board_x[2] ),
    .B(_1500_),
    .C(_2758_),
    .Y(_3218_));
 sg13g2_or4_2 _7603_ (.A(_1415_),
    .B(_3214_),
    .C(_3217_),
    .D(_3218_),
    .X(_3219_));
 sg13g2_and2_1 _7604_ (.A(_3213_),
    .B(_3219_),
    .X(_3220_));
 sg13g2_nand2_1 _7605_ (.Y(_3221_),
    .A(_3211_),
    .B(_3220_));
 sg13g2_inv_1 _7606_ (.Y(_3222_),
    .A(_3221_));
 sg13g2_nor2_1 _7607_ (.A(_1425_),
    .B(_3210_),
    .Y(_3223_));
 sg13g2_mux2_1 _7608_ (.A0(\draw_game_inst.new_tiles[15] ),
    .A1(\draw_game_inst.new_tiles[14] ),
    .S(net2129),
    .X(_3224_));
 sg13g2_a21oi_1 _7609_ (.A1(\draw_game_inst.new_tiles[13] ),
    .A2(net1978),
    .Y(_3225_),
    .B1(_3993_));
 sg13g2_a22oi_1 _7610_ (.Y(_3226_),
    .B1(_1427_),
    .B2(_3224_),
    .A2(net1980),
    .A1(\draw_game_inst.new_tiles[12] ));
 sg13g2_mux2_1 _7611_ (.A0(\draw_game_inst.new_tiles[11] ),
    .A1(\draw_game_inst.new_tiles[10] ),
    .S(net2129),
    .X(_3227_));
 sg13g2_a21oi_1 _7612_ (.A1(\draw_game_inst.new_tiles[9] ),
    .A2(net1978),
    .Y(_3228_),
    .B1(net2154));
 sg13g2_a22oi_1 _7613_ (.Y(_3229_),
    .B1(_1427_),
    .B2(_3227_),
    .A2(net1979),
    .A1(\draw_game_inst.new_tiles[8] ));
 sg13g2_a221oi_1 _7614_ (.B2(_3229_),
    .C1(net2153),
    .B1(_3228_),
    .A1(_3225_),
    .Y(_3230_),
    .A2(_3226_));
 sg13g2_mux4_1 _7615_ (.S0(net2129),
    .A0(\draw_game_inst.new_tiles[1] ),
    .A1(\draw_game_inst.new_tiles[2] ),
    .A2(\draw_game_inst.new_tiles[3] ),
    .A3(\draw_game_inst.new_tiles[0] ),
    .S1(net2125),
    .X(_3231_));
 sg13g2_mux4_1 _7616_ (.S0(net2129),
    .A0(\draw_game_inst.new_tiles[5] ),
    .A1(\draw_game_inst.new_tiles[6] ),
    .A2(\draw_game_inst.new_tiles[7] ),
    .A3(\draw_game_inst.new_tiles[4] ),
    .S1(net2125),
    .X(_3232_));
 sg13g2_a221oi_1 _7617_ (.B2(_1398_),
    .C1(_3230_),
    .B1(_3232_),
    .A1(_1409_),
    .Y(_3233_),
    .A2(_3231_));
 sg13g2_nor3_1 _7618_ (.A(\draw_game_inst.new_tiles_counter[0] ),
    .B(\draw_game_inst.new_tiles_counter[1] ),
    .C(_4008_),
    .Y(_3234_));
 sg13g2_nor2_1 _7619_ (.A(_3233_),
    .B(_3234_),
    .Y(_3235_));
 sg13g2_mux2_1 _7620_ (.A0(_3213_),
    .A1(net1044),
    .S(_3235_),
    .X(_3236_));
 sg13g2_nor4_1 _7621_ (.A(_3976_),
    .B(\draw_game_inst.x[9] ),
    .C(net2157),
    .D(_3995_),
    .Y(_3237_));
 sg13g2_o21ai_1 _7622_ (.B1(_3237_),
    .Y(_3238_),
    .A1(net2122),
    .A2(net2123));
 sg13g2_nor4_2 _7623_ (.A(net2153),
    .B(net2154),
    .C(_1416_),
    .Y(_3239_),
    .D(_3238_));
 sg13g2_nor2b_2 _7624_ (.A(_1424_),
    .B_N(_3239_),
    .Y(_3240_));
 sg13g2_a221oi_1 _7625_ (.B2(net2147),
    .C1(_3222_),
    .B1(_3240_),
    .A1(_3223_),
    .Y(_3241_),
    .A2(_3236_));
 sg13g2_nor2_1 _7626_ (.A(_1408_),
    .B(_3241_),
    .Y(_0177_));
 sg13g2_nand2b_1 _7627_ (.Y(_3242_),
    .B(net837),
    .A_N(_3233_));
 sg13g2_a22oi_1 _7628_ (.Y(_3243_),
    .B1(_3242_),
    .B2(_3223_),
    .A2(_3240_),
    .A1(net2144));
 sg13g2_a21oi_1 _7629_ (.A1(_3221_),
    .A2(_3243_),
    .Y(_0178_),
    .B1(_1408_));
 sg13g2_nor3_1 _7630_ (.A(_3963_),
    .B(_3213_),
    .C(_3219_),
    .Y(_3244_));
 sg13g2_o21ai_1 _7631_ (.B1(_3211_),
    .Y(_3245_),
    .A1(_3220_),
    .A2(_3244_));
 sg13g2_nand2_1 _7632_ (.Y(_3246_),
    .A(net1037),
    .B(_3235_));
 sg13g2_a22oi_1 _7633_ (.Y(_3247_),
    .B1(_3246_),
    .B2(_3223_),
    .A2(_3240_),
    .A1(net2135));
 sg13g2_a21oi_1 _7634_ (.A1(_3245_),
    .A2(_3247_),
    .Y(_0179_),
    .B1(_1408_));
 sg13g2_nor2_1 _7635_ (.A(_3212_),
    .B(_3219_),
    .Y(_3248_));
 sg13g2_a21oi_1 _7636_ (.A1(net2129),
    .A2(_3239_),
    .Y(_3249_),
    .B1(_1424_));
 sg13g2_nor3_2 _7637_ (.A(_1408_),
    .B(_3248_),
    .C(net1043),
    .Y(_0180_));
 sg13g2_nand2_1 _7638_ (.Y(_3250_),
    .A(net2123),
    .B(_3240_));
 sg13g2_a21oi_1 _7639_ (.A1(_3221_),
    .A2(_3250_),
    .Y(_0181_),
    .B1(_1408_));
 sg13g2_or4_1 _7640_ (.A(_1425_),
    .B(_3210_),
    .C(_3213_),
    .D(_3235_),
    .X(_3251_));
 sg13g2_a21oi_1 _7641_ (.A1(net2122),
    .A2(_3240_),
    .Y(_3252_),
    .B1(_3222_));
 sg13g2_a21oi_1 _7642_ (.A1(_3251_),
    .A2(_3252_),
    .Y(_0182_),
    .B1(_1408_));
 sg13g2_nand2_1 _7643_ (.Y(_3253_),
    .A(net2061),
    .B(\debug_controller_inst.grid_in[0] ));
 sg13g2_nor2b_2 _7644_ (.A(vsync_prev),
    .B_N(\vga_sync_gen.vsync ),
    .Y(_3254_));
 sg13g2_nand2b_2 _7645_ (.Y(_3255_),
    .B(\vga_sync_gen.vsync ),
    .A_N(vsync_prev));
 sg13g2_a21oi_2 _7646_ (.B1(net1926),
    .Y(_3256_),
    .A2(\welcome_screen_grid[0] ),
    .A1(net2255));
 sg13g2_nor2_1 _7647_ (.A(net2257),
    .B(net1926),
    .Y(_3257_));
 sg13g2_nand2_1 _7648_ (.Y(_3258_),
    .A(net2289),
    .B(_3254_));
 sg13g2_nand2_1 _7649_ (.Y(_3259_),
    .A(net521),
    .B(net2272));
 sg13g2_a22oi_1 _7650_ (.Y(_0183_),
    .B1(net1824),
    .B2(_3259_),
    .A2(_3256_),
    .A1(_3253_));
 sg13g2_nand2_1 _7651_ (.Y(_3260_),
    .A(net2066),
    .B(\debug_controller_inst.grid_in[1] ));
 sg13g2_nand2_1 _7652_ (.Y(_3261_),
    .A(net513),
    .B(net2272));
 sg13g2_a22oi_1 _7653_ (.Y(_0184_),
    .B1(_3261_),
    .B2(net1825),
    .A2(_3260_),
    .A1(_3256_));
 sg13g2_nor2_2 _7654_ (.A(net2260),
    .B(_3254_),
    .Y(_3262_));
 sg13g2_nor2_2 _7655_ (.A(net2255),
    .B(net1824),
    .Y(_3263_));
 sg13g2_a22oi_1 _7656_ (.Y(_3264_),
    .B1(net1792),
    .B2(\debug_controller_inst.grid_in[2] ),
    .A2(net1823),
    .A1(net482));
 sg13g2_inv_1 _7657_ (.Y(_0185_),
    .A(net483));
 sg13g2_nand2_1 _7658_ (.Y(_3265_),
    .A(net2061),
    .B(\debug_controller_inst.grid_in[3] ));
 sg13g2_nand2_1 _7659_ (.Y(_3266_),
    .A(net597),
    .B(net2273));
 sg13g2_a22oi_1 _7660_ (.Y(_0186_),
    .B1(_3266_),
    .B2(net1824),
    .A2(_3265_),
    .A1(_3256_));
 sg13g2_nand2_1 _7661_ (.Y(_3267_),
    .A(net2061),
    .B(\debug_controller_inst.grid_in[4] ));
 sg13g2_a21oi_2 _7662_ (.B1(net1926),
    .Y(_3268_),
    .A2(\welcome_screen_grid[4] ),
    .A1(net2255));
 sg13g2_nand2_1 _7663_ (.Y(_3269_),
    .A(net681),
    .B(net2272));
 sg13g2_a22oi_1 _7664_ (.Y(_0187_),
    .B1(_3269_),
    .B2(net1824),
    .A2(_3268_),
    .A1(_3267_));
 sg13g2_nand2_1 _7665_ (.Y(_3270_),
    .A(net2061),
    .B(\debug_controller_inst.grid_in[5] ));
 sg13g2_nand2_1 _7666_ (.Y(_3271_),
    .A(net697),
    .B(net2273));
 sg13g2_a22oi_1 _7667_ (.Y(_0188_),
    .B1(_3271_),
    .B2(net1824),
    .A2(_3270_),
    .A1(_3268_));
 sg13g2_a22oi_1 _7668_ (.Y(_3272_),
    .B1(net1792),
    .B2(\debug_controller_inst.grid_in[6] ),
    .A2(net1823),
    .A1(net495));
 sg13g2_inv_1 _7669_ (.Y(_0189_),
    .A(net496));
 sg13g2_nand2_1 _7670_ (.Y(_3273_),
    .A(net2061),
    .B(\debug_controller_inst.grid_in[7] ));
 sg13g2_nand2_1 _7671_ (.Y(_3274_),
    .A(net691),
    .B(net2272));
 sg13g2_a22oi_1 _7672_ (.Y(_0190_),
    .B1(_3274_),
    .B2(net1824),
    .A2(_3273_),
    .A1(_3268_));
 sg13g2_a21oi_2 _7673_ (.B1(net1926),
    .Y(_3275_),
    .A2(\welcome_screen_grid[11] ),
    .A1(net2255));
 sg13g2_nand2_1 _7674_ (.Y(_3276_),
    .A(net2066),
    .B(\debug_controller_inst.grid_in[8] ));
 sg13g2_nand2_1 _7675_ (.Y(_3277_),
    .A(net632),
    .B(net2272));
 sg13g2_a22oi_1 _7676_ (.Y(_0191_),
    .B1(_3277_),
    .B2(net1825),
    .A2(_3276_),
    .A1(_3275_));
 sg13g2_nand2_1 _7677_ (.Y(_3278_),
    .A(net2066),
    .B(\debug_controller_inst.grid_in[9] ));
 sg13g2_nand2_1 _7678_ (.Y(_3279_),
    .A(net586),
    .B(net2273));
 sg13g2_a22oi_1 _7679_ (.Y(_0192_),
    .B1(_3279_),
    .B2(net1825),
    .A2(_3278_),
    .A1(_3275_));
 sg13g2_a22oi_1 _7680_ (.Y(_3280_),
    .B1(net1792),
    .B2(\debug_controller_inst.grid_in[10] ),
    .A2(net1822),
    .A1(net507));
 sg13g2_inv_1 _7681_ (.Y(_0193_),
    .A(net508));
 sg13g2_nand2_1 _7682_ (.Y(_3281_),
    .A(net2066),
    .B(\debug_controller_inst.grid_in[11] ));
 sg13g2_nand2_1 _7683_ (.Y(_3282_),
    .A(net675),
    .B(net2273));
 sg13g2_a22oi_1 _7684_ (.Y(_0194_),
    .B1(_3282_),
    .B2(net1824),
    .A2(_3281_),
    .A1(_3275_));
 sg13g2_nand2_1 _7685_ (.Y(_3283_),
    .A(net2064),
    .B(\debug_controller_inst.grid_in[12] ));
 sg13g2_a21oi_2 _7686_ (.B1(net1926),
    .Y(_3284_),
    .A2(\welcome_screen_grid[12] ),
    .A1(net2255));
 sg13g2_nand2_1 _7687_ (.Y(_3285_),
    .A(net560),
    .B(net2272));
 sg13g2_a22oi_1 _7688_ (.Y(_0195_),
    .B1(_3285_),
    .B2(net1824),
    .A2(_3284_),
    .A1(_3283_));
 sg13g2_nand2_1 _7689_ (.Y(_3286_),
    .A(net2061),
    .B(\debug_controller_inst.grid_in[13] ));
 sg13g2_nand2_1 _7690_ (.Y(_3287_),
    .A(net577),
    .B(net2272));
 sg13g2_a22oi_1 _7691_ (.Y(_0196_),
    .B1(_3287_),
    .B2(net1825),
    .A2(_3286_),
    .A1(_3284_));
 sg13g2_a22oi_1 _7692_ (.Y(_3288_),
    .B1(net1792),
    .B2(\debug_controller_inst.grid_in[14] ),
    .A2(net1822),
    .A1(net543));
 sg13g2_inv_1 _7693_ (.Y(_0197_),
    .A(net544));
 sg13g2_nand2_1 _7694_ (.Y(_3289_),
    .A(net2066),
    .B(net449));
 sg13g2_nand2_1 _7695_ (.Y(_3290_),
    .A(\draw_game_inst.grid[15] ),
    .B(net2272));
 sg13g2_a22oi_1 _7696_ (.Y(_0198_),
    .B1(_3290_),
    .B2(net1825),
    .A2(_3289_),
    .A1(_3284_));
 sg13g2_nand2_1 _7697_ (.Y(_3291_),
    .A(net2062),
    .B(\debug_controller_inst.grid_in[16] ));
 sg13g2_a21oi_2 _7698_ (.B1(net1925),
    .Y(_3292_),
    .A2(\welcome_screen_grid[16] ),
    .A1(net2254));
 sg13g2_nand2_1 _7699_ (.Y(_3293_),
    .A(net552),
    .B(net2282));
 sg13g2_a22oi_1 _7700_ (.Y(_0199_),
    .B1(_3293_),
    .B2(net1826),
    .A2(_3292_),
    .A1(_3291_));
 sg13g2_nand2_1 _7701_ (.Y(_3294_),
    .A(net2062),
    .B(\debug_controller_inst.grid_in[17] ));
 sg13g2_nand2_1 _7702_ (.Y(_3295_),
    .A(net660),
    .B(net2282));
 sg13g2_a22oi_1 _7703_ (.Y(_0200_),
    .B1(_3295_),
    .B2(net1826),
    .A2(_3294_),
    .A1(_3292_));
 sg13g2_a22oi_1 _7704_ (.Y(_3296_),
    .B1(net1793),
    .B2(\debug_controller_inst.grid_in[18] ),
    .A2(net1823),
    .A1(net554));
 sg13g2_inv_1 _7705_ (.Y(_0201_),
    .A(net555));
 sg13g2_nand2_1 _7706_ (.Y(_3297_),
    .A(net2062),
    .B(\debug_controller_inst.grid_in[19] ));
 sg13g2_nand2_1 _7707_ (.Y(_3298_),
    .A(net604),
    .B(net2280));
 sg13g2_a22oi_1 _7708_ (.Y(_0202_),
    .B1(_3298_),
    .B2(net1826),
    .A2(_3297_),
    .A1(_3292_));
 sg13g2_nand2_1 _7709_ (.Y(_3299_),
    .A(net2062),
    .B(\debug_controller_inst.grid_in[20] ));
 sg13g2_a21oi_2 _7710_ (.B1(net1925),
    .Y(_3300_),
    .A2(\welcome_screen_grid[20] ),
    .A1(net2254));
 sg13g2_nand2_1 _7711_ (.Y(_3301_),
    .A(net615),
    .B(net2282));
 sg13g2_a22oi_1 _7712_ (.Y(_0203_),
    .B1(_3301_),
    .B2(net1826),
    .A2(_3300_),
    .A1(_3299_));
 sg13g2_nand2_1 _7713_ (.Y(_3302_),
    .A(net2061),
    .B(\debug_controller_inst.grid_in[21] ));
 sg13g2_nand2_1 _7714_ (.Y(_3303_),
    .A(net564),
    .B(net2280));
 sg13g2_a22oi_1 _7715_ (.Y(_0204_),
    .B1(_3303_),
    .B2(net1827),
    .A2(_3302_),
    .A1(_3300_));
 sg13g2_a22oi_1 _7716_ (.Y(_3304_),
    .B1(net1792),
    .B2(\debug_controller_inst.grid_in[22] ),
    .A2(net1822),
    .A1(net623));
 sg13g2_inv_1 _7717_ (.Y(_0205_),
    .A(net624));
 sg13g2_nand2_1 _7718_ (.Y(_3305_),
    .A(net2062),
    .B(\debug_controller_inst.grid_in[23] ));
 sg13g2_nand2_1 _7719_ (.Y(_3306_),
    .A(net646),
    .B(net2280));
 sg13g2_a22oi_1 _7720_ (.Y(_0206_),
    .B1(_3306_),
    .B2(net1826),
    .A2(_3305_),
    .A1(_3300_));
 sg13g2_nand2_1 _7721_ (.Y(_3307_),
    .A(net2062),
    .B(\debug_controller_inst.grid_in[24] ));
 sg13g2_a21oi_2 _7722_ (.B1(net1924),
    .Y(_3308_),
    .A2(\welcome_screen_grid[24] ),
    .A1(net2254));
 sg13g2_nand2_1 _7723_ (.Y(_3309_),
    .A(net621),
    .B(net2282));
 sg13g2_a22oi_1 _7724_ (.Y(_0207_),
    .B1(_3309_),
    .B2(net1827),
    .A2(_3308_),
    .A1(_3307_));
 sg13g2_nand2_1 _7725_ (.Y(_3310_),
    .A(net2062),
    .B(\debug_controller_inst.grid_in[25] ));
 sg13g2_nand2_1 _7726_ (.Y(_3311_),
    .A(net591),
    .B(net2280));
 sg13g2_a22oi_1 _7727_ (.Y(_0208_),
    .B1(_3311_),
    .B2(net1827),
    .A2(_3310_),
    .A1(_3308_));
 sg13g2_a22oi_1 _7728_ (.Y(_3312_),
    .B1(net1793),
    .B2(\debug_controller_inst.grid_in[26] ),
    .A2(_3262_),
    .A1(net630));
 sg13g2_inv_1 _7729_ (.Y(_0209_),
    .A(net631));
 sg13g2_nand2_1 _7730_ (.Y(_3313_),
    .A(net2067),
    .B(\debug_controller_inst.grid_in[27] ));
 sg13g2_nand2_1 _7731_ (.Y(_3314_),
    .A(net638),
    .B(net2280));
 sg13g2_a22oi_1 _7732_ (.Y(_0210_),
    .B1(_3314_),
    .B2(net1827),
    .A2(_3313_),
    .A1(_3308_));
 sg13g2_nand2_1 _7733_ (.Y(_3315_),
    .A(net2063),
    .B(\debug_controller_inst.grid_in[28] ));
 sg13g2_a21oi_2 _7734_ (.B1(net1925),
    .Y(_3316_),
    .A2(\welcome_screen_grid[28] ),
    .A1(net2254));
 sg13g2_nand2_1 _7735_ (.Y(_3317_),
    .A(net599),
    .B(net2282));
 sg13g2_a22oi_1 _7736_ (.Y(_0211_),
    .B1(_3317_),
    .B2(net1826),
    .A2(_3316_),
    .A1(_3315_));
 sg13g2_nand2_1 _7737_ (.Y(_3318_),
    .A(net2062),
    .B(\debug_controller_inst.grid_in[29] ));
 sg13g2_nand2_1 _7738_ (.Y(_3319_),
    .A(net617),
    .B(net2280));
 sg13g2_a22oi_1 _7739_ (.Y(_0212_),
    .B1(_3319_),
    .B2(net1826),
    .A2(_3318_),
    .A1(_3316_));
 sg13g2_a22oi_1 _7740_ (.Y(_3320_),
    .B1(net1792),
    .B2(\debug_controller_inst.grid_in[30] ),
    .A2(net1822),
    .A1(net658));
 sg13g2_inv_1 _7741_ (.Y(_0213_),
    .A(net659));
 sg13g2_nand2_1 _7742_ (.Y(_3321_),
    .A(net2063),
    .B(\debug_controller_inst.grid_in[31] ));
 sg13g2_nand2_1 _7743_ (.Y(_3322_),
    .A(net613),
    .B(net2280));
 sg13g2_a22oi_1 _7744_ (.Y(_0214_),
    .B1(_3322_),
    .B2(net1826),
    .A2(_3321_),
    .A1(_3316_));
 sg13g2_nand2_1 _7745_ (.Y(_3323_),
    .A(net2066),
    .B(\debug_controller_inst.grid_in[32] ));
 sg13g2_a21oi_2 _7746_ (.B1(net1924),
    .Y(_3324_),
    .A2(\welcome_screen_grid[32] ),
    .A1(net2255));
 sg13g2_nand2_1 _7747_ (.Y(_3325_),
    .A(net541),
    .B(net2281));
 sg13g2_a22oi_1 _7748_ (.Y(_0215_),
    .B1(_3325_),
    .B2(net1829),
    .A2(_3324_),
    .A1(_3323_));
 sg13g2_nand2_1 _7749_ (.Y(_3326_),
    .A(net2065),
    .B(\debug_controller_inst.grid_in[33] ));
 sg13g2_nand2_1 _7750_ (.Y(_3327_),
    .A(net490),
    .B(net2288));
 sg13g2_a22oi_1 _7751_ (.Y(_0216_),
    .B1(_3327_),
    .B2(net1829),
    .A2(_3326_),
    .A1(_3324_));
 sg13g2_a22oi_1 _7752_ (.Y(_3328_),
    .B1(net1793),
    .B2(\debug_controller_inst.grid_in[34] ),
    .A2(net1823),
    .A1(net480));
 sg13g2_inv_1 _7753_ (.Y(_0217_),
    .A(net481));
 sg13g2_nand2_1 _7754_ (.Y(_3329_),
    .A(net2065),
    .B(\debug_controller_inst.grid_in[35] ));
 sg13g2_nand2_1 _7755_ (.Y(_3330_),
    .A(net484),
    .B(net2288));
 sg13g2_a22oi_1 _7756_ (.Y(_0218_),
    .B1(_3330_),
    .B2(net1829),
    .A2(_3329_),
    .A1(_3324_));
 sg13g2_nand2_1 _7757_ (.Y(_3331_),
    .A(net2066),
    .B(\debug_controller_inst.grid_in[36] ));
 sg13g2_a21oi_2 _7758_ (.B1(net1924),
    .Y(_3332_),
    .A2(\welcome_screen_grid[36] ),
    .A1(net2254));
 sg13g2_nand2_1 _7759_ (.Y(_3333_),
    .A(net562),
    .B(net2281));
 sg13g2_a22oi_1 _7760_ (.Y(_0219_),
    .B1(_3333_),
    .B2(net1829),
    .A2(_3332_),
    .A1(_3331_));
 sg13g2_nand2_1 _7761_ (.Y(_3334_),
    .A(net2068),
    .B(\debug_controller_inst.grid_in[37] ));
 sg13g2_nand2_1 _7762_ (.Y(_3335_),
    .A(net519),
    .B(net2288));
 sg13g2_a22oi_1 _7763_ (.Y(_0220_),
    .B1(_3335_),
    .B2(net1831),
    .A2(_3334_),
    .A1(_3332_));
 sg13g2_a22oi_1 _7764_ (.Y(_3336_),
    .B1(net1793),
    .B2(\debug_controller_inst.grid_in[38] ),
    .A2(net1823),
    .A1(net535));
 sg13g2_inv_1 _7765_ (.Y(_0221_),
    .A(net536));
 sg13g2_nand2_1 _7766_ (.Y(_3337_),
    .A(net2068),
    .B(\debug_controller_inst.grid_in[39] ));
 sg13g2_nand2_1 _7767_ (.Y(_3338_),
    .A(net523),
    .B(net2288));
 sg13g2_a22oi_1 _7768_ (.Y(_0222_),
    .B1(_3338_),
    .B2(net1830),
    .A2(_3337_),
    .A1(_3332_));
 sg13g2_nand2_1 _7769_ (.Y(_3339_),
    .A(net2065),
    .B(\debug_controller_inst.grid_in[40] ));
 sg13g2_a21oi_2 _7770_ (.B1(net1926),
    .Y(_3340_),
    .A2(\welcome_screen_grid[40] ),
    .A1(net2255));
 sg13g2_nand2_1 _7771_ (.Y(_3341_),
    .A(net668),
    .B(net2273));
 sg13g2_a22oi_1 _7772_ (.Y(_0223_),
    .B1(_3341_),
    .B2(net1829),
    .A2(_3340_),
    .A1(_3339_));
 sg13g2_nand2_1 _7773_ (.Y(_3342_),
    .A(net2068),
    .B(\debug_controller_inst.grid_in[41] ));
 sg13g2_nand2_1 _7774_ (.Y(_3343_),
    .A(net515),
    .B(net2288));
 sg13g2_a22oi_1 _7775_ (.Y(_0224_),
    .B1(_3343_),
    .B2(net1829),
    .A2(_3342_),
    .A1(_3340_));
 sg13g2_a22oi_1 _7776_ (.Y(_3344_),
    .B1(net1793),
    .B2(\debug_controller_inst.grid_in[42] ),
    .A2(net1822),
    .A1(net527));
 sg13g2_inv_1 _7777_ (.Y(_0225_),
    .A(net528));
 sg13g2_nand2_1 _7778_ (.Y(_3345_),
    .A(net2065),
    .B(\debug_controller_inst.grid_in[43] ));
 sg13g2_nand2_1 _7779_ (.Y(_3346_),
    .A(net537),
    .B(net2278));
 sg13g2_a22oi_1 _7780_ (.Y(_0226_),
    .B1(_3346_),
    .B2(net1831),
    .A2(_3345_),
    .A1(_3340_));
 sg13g2_nand2_1 _7781_ (.Y(_3347_),
    .A(net2065),
    .B(\debug_controller_inst.grid_in[44] ));
 sg13g2_a21oi_2 _7782_ (.B1(net1924),
    .Y(_3348_),
    .A2(\welcome_screen_grid[44] ),
    .A1(net2255));
 sg13g2_nand2_1 _7783_ (.Y(_3349_),
    .A(net619),
    .B(net2281));
 sg13g2_a22oi_1 _7784_ (.Y(_0227_),
    .B1(_3349_),
    .B2(net1829),
    .A2(_3348_),
    .A1(_3347_));
 sg13g2_nand2_1 _7785_ (.Y(_3350_),
    .A(net2065),
    .B(\debug_controller_inst.grid_in[45] ));
 sg13g2_nand2_1 _7786_ (.Y(_3351_),
    .A(net463),
    .B(net2288));
 sg13g2_a22oi_1 _7787_ (.Y(_0228_),
    .B1(_3351_),
    .B2(net1831),
    .A2(_3350_),
    .A1(_3348_));
 sg13g2_a22oi_1 _7788_ (.Y(_3352_),
    .B1(net1793),
    .B2(\debug_controller_inst.grid_in[46] ),
    .A2(net1822),
    .A1(net488));
 sg13g2_inv_1 _7789_ (.Y(_0229_),
    .A(net489));
 sg13g2_nand2_1 _7790_ (.Y(_3353_),
    .A(net2065),
    .B(\debug_controller_inst.grid_in[47] ));
 sg13g2_nand2_1 _7791_ (.Y(_3354_),
    .A(net529),
    .B(net2278));
 sg13g2_a22oi_1 _7792_ (.Y(_0230_),
    .B1(_3354_),
    .B2(net1829),
    .A2(_3353_),
    .A1(_3348_));
 sg13g2_nand2_1 _7793_ (.Y(_3355_),
    .A(net2067),
    .B(\debug_controller_inst.grid_in[48] ));
 sg13g2_a21oi_2 _7794_ (.B1(net1924),
    .Y(_3356_),
    .A2(\welcome_screen_grid[48] ),
    .A1(net2256));
 sg13g2_nand2_1 _7795_ (.Y(_3357_),
    .A(net693),
    .B(net2283));
 sg13g2_a22oi_1 _7796_ (.Y(_0231_),
    .B1(_3357_),
    .B2(net1827),
    .A2(_3356_),
    .A1(_3355_));
 sg13g2_nand2_1 _7797_ (.Y(_3358_),
    .A(net2067),
    .B(\debug_controller_inst.grid_in[49] ));
 sg13g2_nand2_1 _7798_ (.Y(_3359_),
    .A(net679),
    .B(net2283));
 sg13g2_a22oi_1 _7799_ (.Y(_0232_),
    .B1(_3359_),
    .B2(net1830),
    .A2(_3358_),
    .A1(_3356_));
 sg13g2_a22oi_1 _7800_ (.Y(_3360_),
    .B1(_3263_),
    .B2(\debug_controller_inst.grid_in[50] ),
    .A2(net1823),
    .A1(net569));
 sg13g2_inv_1 _7801_ (.Y(_0233_),
    .A(net570));
 sg13g2_nand2_1 _7802_ (.Y(_3361_),
    .A(net2067),
    .B(\debug_controller_inst.grid_in[51] ));
 sg13g2_nand2_1 _7803_ (.Y(_3362_),
    .A(net573),
    .B(net2280));
 sg13g2_a22oi_1 _7804_ (.Y(_0234_),
    .B1(_3362_),
    .B2(net1830),
    .A2(_3361_),
    .A1(_3356_));
 sg13g2_nand2_1 _7805_ (.Y(_3363_),
    .A(net2067),
    .B(\debug_controller_inst.grid_in[52] ));
 sg13g2_a21oi_2 _7806_ (.B1(net1924),
    .Y(_3364_),
    .A2(\welcome_screen_grid[52] ),
    .A1(net2254));
 sg13g2_nand2_1 _7807_ (.Y(_3365_),
    .A(net545),
    .B(net2283));
 sg13g2_a22oi_1 _7808_ (.Y(_0235_),
    .B1(_3365_),
    .B2(net1827),
    .A2(_3364_),
    .A1(_3363_));
 sg13g2_nand2_1 _7809_ (.Y(_3366_),
    .A(net2065),
    .B(\debug_controller_inst.grid_in[53] ));
 sg13g2_nand2_1 _7810_ (.Y(_3367_),
    .A(net558),
    .B(net2291));
 sg13g2_a22oi_1 _7811_ (.Y(_0236_),
    .B1(_3367_),
    .B2(net1830),
    .A2(_3366_),
    .A1(_3364_));
 sg13g2_a22oi_1 _7812_ (.Y(_3368_),
    .B1(net1793),
    .B2(\debug_controller_inst.grid_in[54] ),
    .A2(net1823),
    .A1(net517));
 sg13g2_inv_1 _7813_ (.Y(_0237_),
    .A(net518));
 sg13g2_nand2_1 _7814_ (.Y(_3369_),
    .A(net2066),
    .B(\debug_controller_inst.grid_in[55] ));
 sg13g2_nand2_1 _7815_ (.Y(_3370_),
    .A(net533),
    .B(net2288));
 sg13g2_a22oi_1 _7816_ (.Y(_0238_),
    .B1(_3370_),
    .B2(net1830),
    .A2(_3369_),
    .A1(_3364_));
 sg13g2_nand2_1 _7817_ (.Y(_3371_),
    .A(net2067),
    .B(\debug_controller_inst.grid_in[56] ));
 sg13g2_a21oi_2 _7818_ (.B1(net1924),
    .Y(_3372_),
    .A2(\welcome_screen_grid[56] ),
    .A1(net2254));
 sg13g2_nand2_1 _7819_ (.Y(_3373_),
    .A(net636),
    .B(net2283));
 sg13g2_a22oi_1 _7820_ (.Y(_0239_),
    .B1(_3373_),
    .B2(net1830),
    .A2(_3372_),
    .A1(_3371_));
 sg13g2_nand2_1 _7821_ (.Y(_3374_),
    .A(net2067),
    .B(\debug_controller_inst.grid_in[57] ));
 sg13g2_nand2_1 _7822_ (.Y(_3375_),
    .A(net644),
    .B(net2281));
 sg13g2_a22oi_1 _7823_ (.Y(_0240_),
    .B1(_3375_),
    .B2(net1830),
    .A2(_3374_),
    .A1(_3372_));
 sg13g2_a22oi_1 _7824_ (.Y(_3376_),
    .B1(net1792),
    .B2(\debug_controller_inst.grid_in[58] ),
    .A2(net1822),
    .A1(net579));
 sg13g2_inv_1 _7825_ (.Y(_0241_),
    .A(net580));
 sg13g2_nand2_1 _7826_ (.Y(_3377_),
    .A(net2067),
    .B(\debug_controller_inst.grid_in[59] ));
 sg13g2_nand2_1 _7827_ (.Y(_3378_),
    .A(net539),
    .B(net2281));
 sg13g2_a22oi_1 _7828_ (.Y(_0242_),
    .B1(_3378_),
    .B2(net1830),
    .A2(_3377_),
    .A1(_3372_));
 sg13g2_nand2_1 _7829_ (.Y(_3379_),
    .A(net2063),
    .B(\debug_controller_inst.grid_in[60] ));
 sg13g2_a21oi_2 _7830_ (.B1(net1924),
    .Y(_3380_),
    .A2(\welcome_screen_grid[60] ),
    .A1(net2254));
 sg13g2_nand2_1 _7831_ (.Y(_3381_),
    .A(net706),
    .B(net2283));
 sg13g2_a22oi_1 _7832_ (.Y(_0243_),
    .B1(_3381_),
    .B2(net1828),
    .A2(_3380_),
    .A1(_3379_));
 sg13g2_nand2_1 _7833_ (.Y(_3382_),
    .A(net2063),
    .B(\debug_controller_inst.grid_in[61] ));
 sg13g2_nand2_1 _7834_ (.Y(_3383_),
    .A(net556),
    .B(net2281));
 sg13g2_a22oi_1 _7835_ (.Y(_0244_),
    .B1(_3383_),
    .B2(net1827),
    .A2(_3382_),
    .A1(_3380_));
 sg13g2_a22oi_1 _7836_ (.Y(_3384_),
    .B1(net1792),
    .B2(\debug_controller_inst.grid_in[62] ),
    .A2(net1822),
    .A1(net471));
 sg13g2_inv_1 _7837_ (.Y(_0245_),
    .A(net472));
 sg13g2_nand2_1 _7838_ (.Y(_3385_),
    .A(net2063),
    .B(\debug_controller_inst.grid_in[63] ));
 sg13g2_nand2_1 _7839_ (.Y(_3386_),
    .A(net548),
    .B(net2281));
 sg13g2_a22oi_1 _7840_ (.Y(_0246_),
    .B1(_3386_),
    .B2(net1828),
    .A2(_3385_),
    .A1(_3380_));
 sg13g2_nand2_2 _7841_ (.Y(_3387_),
    .A(net758),
    .B(_0509_));
 sg13g2_nor3_1 _7842_ (.A(_0512_),
    .B(_0514_),
    .C(_0516_),
    .Y(_3388_));
 sg13g2_nand3b_1 _7843_ (.B(_3387_),
    .C(_3388_),
    .Y(_3389_),
    .A_N(_0510_));
 sg13g2_a22oi_1 _7844_ (.Y(_0247_),
    .B1(_3257_),
    .B2(_3389_),
    .A2(net2271),
    .A1(net2061));
 sg13g2_nand2_1 _7845_ (.Y(_3390_),
    .A(net703),
    .B(_0509_));
 sg13g2_nor2_1 _7846_ (.A(net2259),
    .B(_3390_),
    .Y(_0248_));
 sg13g2_nor2_1 _7847_ (.A(net798),
    .B(\new_tiles_counter[0] ),
    .Y(_3391_));
 sg13g2_nand2b_1 _7848_ (.Y(_3392_),
    .B(_3391_),
    .A_N(\draw_game_inst.new_tiles_counter[1] ));
 sg13g2_nand3b_1 _7849_ (.B(_4006_),
    .C(_4005_),
    .Y(_3393_),
    .A_N(_3392_));
 sg13g2_o21ai_1 _7850_ (.B1(net451),
    .Y(_3394_),
    .A1(net1832),
    .A2(_3393_));
 sg13g2_inv_1 _7851_ (.Y(_0249_),
    .A(net452));
 sg13g2_nand2_1 _7852_ (.Y(_3395_),
    .A(net2261),
    .B(net473));
 sg13g2_nand2b_1 _7853_ (.Y(_3396_),
    .B(\game_logic_inst.added_tile_index[0] ),
    .A_N(\game_logic_inst.added_tile_index[1] ));
 sg13g2_nor3_1 _7854_ (.A(net2100),
    .B(net2101),
    .C(_3396_),
    .Y(_3397_));
 sg13g2_nor2b_1 _7855_ (.A(_3397_),
    .B_N(_0070_),
    .Y(_3398_));
 sg13g2_o21ai_1 _7856_ (.B1(net2289),
    .Y(_3399_),
    .A1(_3255_),
    .A2(_3393_));
 sg13g2_o21ai_1 _7857_ (.B1(_3395_),
    .Y(_0250_),
    .A1(_3398_),
    .A2(net1786));
 sg13g2_nand2_1 _7858_ (.Y(_3400_),
    .A(net2262),
    .B(net606));
 sg13g2_nand2b_1 _7859_ (.Y(_3401_),
    .B(\game_logic_inst.added_tile_index[1] ),
    .A_N(\game_logic_inst.added_tile_index[0] ));
 sg13g2_nor3_1 _7860_ (.A(net2100),
    .B(net2101),
    .C(_3401_),
    .Y(_3402_));
 sg13g2_nor2b_1 _7861_ (.A(_3402_),
    .B_N(_0071_),
    .Y(_3403_));
 sg13g2_o21ai_1 _7862_ (.B1(_3400_),
    .Y(_0251_),
    .A1(net1786),
    .A2(_3403_));
 sg13g2_nand2_1 _7863_ (.Y(_3404_),
    .A(net2262),
    .B(net611));
 sg13g2_nand2_1 _7864_ (.Y(_3405_),
    .A(\game_logic_inst.added_tile_index[1] ),
    .B(\game_logic_inst.added_tile_index[0] ));
 sg13g2_nor3_1 _7865_ (.A(net2100),
    .B(net2101),
    .C(_3405_),
    .Y(_3406_));
 sg13g2_nor2b_1 _7866_ (.A(_3406_),
    .B_N(_0072_),
    .Y(_3407_));
 sg13g2_o21ai_1 _7867_ (.B1(_3404_),
    .Y(_0252_),
    .A1(net1786),
    .A2(_3407_));
 sg13g2_nor2_1 _7868_ (.A(\game_logic_inst.added_tile_index[1] ),
    .B(\game_logic_inst.added_tile_index[0] ),
    .Y(_3408_));
 sg13g2_nand3_1 _7869_ (.B(net2101),
    .C(_3408_),
    .A(_4003_),
    .Y(_3409_));
 sg13g2_a21oi_1 _7870_ (.A1(net640),
    .A2(_3409_),
    .Y(_3410_),
    .B1(net1785));
 sg13g2_a21o_1 _7871_ (.A2(\draw_game_inst.new_tiles[4] ),
    .A1(net2262),
    .B1(_3410_),
    .X(_0253_));
 sg13g2_nand3b_1 _7872_ (.B(\game_logic_inst.added_tile_index[0] ),
    .C(net2101),
    .Y(_3411_),
    .A_N(\game_logic_inst.added_tile_index[1] ));
 sg13g2_o21ai_1 _7873_ (.B1(_0074_),
    .Y(_3412_),
    .A1(net2100),
    .A2(_3411_));
 sg13g2_nor2b_1 _7874_ (.A(net1785),
    .B_N(_3412_),
    .Y(_3413_));
 sg13g2_a21o_1 _7875_ (.A2(net792),
    .A1(net2262),
    .B1(_3413_),
    .X(_0254_));
 sg13g2_nand3b_1 _7876_ (.B(\game_logic_inst.added_tile_index[1] ),
    .C(net2102),
    .Y(_3414_),
    .A_N(\game_logic_inst.added_tile_index[0] ));
 sg13g2_o21ai_1 _7877_ (.B1(_0075_),
    .Y(_3415_),
    .A1(net2100),
    .A2(_3414_));
 sg13g2_nor2b_1 _7878_ (.A(net1785),
    .B_N(_3415_),
    .Y(_3416_));
 sg13g2_a21o_1 _7879_ (.A2(net718),
    .A1(net2263),
    .B1(_3416_),
    .X(_0255_));
 sg13g2_nand3_1 _7880_ (.B(\game_logic_inst.added_tile_index[1] ),
    .C(\game_logic_inst.added_tile_index[0] ),
    .A(net2102),
    .Y(_3417_));
 sg13g2_o21ai_1 _7881_ (.B1(_0076_),
    .Y(_3418_),
    .A1(net2100),
    .A2(_3417_));
 sg13g2_nand2b_1 _7882_ (.Y(_3419_),
    .B(_3418_),
    .A_N(net1785));
 sg13g2_o21ai_1 _7883_ (.B1(_3419_),
    .Y(_0256_),
    .A1(net2278),
    .A2(_4007_));
 sg13g2_nor3_1 _7884_ (.A(net2101),
    .B(\game_logic_inst.added_tile_index[1] ),
    .C(\game_logic_inst.added_tile_index[0] ),
    .Y(_3420_));
 sg13g2_nand2_1 _7885_ (.Y(_3421_),
    .A(net2100),
    .B(_3420_));
 sg13g2_a21oi_1 _7886_ (.A1(net666),
    .A2(_3421_),
    .Y(_3422_),
    .B1(net1786));
 sg13g2_a21o_1 _7887_ (.A2(\draw_game_inst.new_tiles[8] ),
    .A1(net2261),
    .B1(_3422_),
    .X(_0257_));
 sg13g2_nand2_1 _7888_ (.Y(_3423_),
    .A(net2261),
    .B(net642));
 sg13g2_nor3_1 _7889_ (.A(_4003_),
    .B(net2101),
    .C(_3396_),
    .Y(_3424_));
 sg13g2_nor2b_1 _7890_ (.A(_3424_),
    .B_N(_0078_),
    .Y(_3425_));
 sg13g2_o21ai_1 _7891_ (.B1(_3423_),
    .Y(_0258_),
    .A1(net1786),
    .A2(_3425_));
 sg13g2_nand2_1 _7892_ (.Y(_3426_),
    .A(net2262),
    .B(net525));
 sg13g2_nor3_1 _7893_ (.A(_4003_),
    .B(net2102),
    .C(_3401_),
    .Y(_3427_));
 sg13g2_nor2b_1 _7894_ (.A(_3427_),
    .B_N(_0079_),
    .Y(_3428_));
 sg13g2_o21ai_1 _7895_ (.B1(_3426_),
    .Y(_0259_),
    .A1(net1786),
    .A2(_3428_));
 sg13g2_or3_1 _7896_ (.A(_4003_),
    .B(net2102),
    .C(_3405_),
    .X(_3429_));
 sg13g2_a21oi_1 _7897_ (.A1(net575),
    .A2(_3429_),
    .Y(_3430_),
    .B1(net1786));
 sg13g2_a21o_1 _7898_ (.A2(\draw_game_inst.new_tiles[11] ),
    .A1(net2261),
    .B1(_3430_),
    .X(_0260_));
 sg13g2_nand3_1 _7899_ (.B(net2101),
    .C(_3408_),
    .A(\game_logic_inst.added_tile_index[3] ),
    .Y(_3431_));
 sg13g2_a21oi_1 _7900_ (.A1(net655),
    .A2(_3431_),
    .Y(_3432_),
    .B1(net1785));
 sg13g2_a21o_1 _7901_ (.A2(\draw_game_inst.new_tiles[12] ),
    .A1(net2261),
    .B1(net656),
    .X(_0261_));
 sg13g2_nand2_1 _7902_ (.Y(_3433_),
    .A(net2261),
    .B(net571));
 sg13g2_nor2_1 _7903_ (.A(_4003_),
    .B(_3411_),
    .Y(_3434_));
 sg13g2_nor2b_1 _7904_ (.A(_3434_),
    .B_N(_0082_),
    .Y(_3435_));
 sg13g2_o21ai_1 _7905_ (.B1(_3433_),
    .Y(_0262_),
    .A1(net1785),
    .A2(_3435_));
 sg13g2_o21ai_1 _7906_ (.B1(_0083_),
    .Y(_3436_),
    .A1(_4003_),
    .A2(_3414_));
 sg13g2_nor2b_1 _7907_ (.A(net1785),
    .B_N(_3436_),
    .Y(_3437_));
 sg13g2_a21o_1 _7908_ (.A2(net745),
    .A1(net2263),
    .B1(_3437_),
    .X(_0263_));
 sg13g2_or2_1 _7909_ (.X(_3438_),
    .B(_3417_),
    .A(_4003_));
 sg13g2_a21oi_1 _7910_ (.A1(net650),
    .A2(_3438_),
    .Y(_3439_),
    .B1(net1785));
 sg13g2_a21o_1 _7911_ (.A2(\draw_game_inst.new_tiles[15] ),
    .A1(net2263),
    .B1(_3439_),
    .X(_0264_));
 sg13g2_and2_1 _7912_ (.A(_3254_),
    .B(_3393_),
    .X(_3440_));
 sg13g2_nand2_1 _7913_ (.Y(_3441_),
    .A(_3254_),
    .B(_3393_));
 sg13g2_and2_1 _7914_ (.A(_4003_),
    .B(_3420_),
    .X(_3442_));
 sg13g2_nand2_1 _7915_ (.Y(_3443_),
    .A(_3441_),
    .B(_3442_));
 sg13g2_o21ai_1 _7916_ (.B1(net2289),
    .Y(_3444_),
    .A1(net446),
    .A2(_3440_));
 sg13g2_a21oi_1 _7917_ (.A1(net446),
    .A2(_3443_),
    .Y(_3445_),
    .B1(_3444_));
 sg13g2_a21oi_1 _7918_ (.A1(net2261),
    .A2(_4004_),
    .Y(_0265_),
    .B1(_3445_));
 sg13g2_o21ai_1 _7919_ (.B1(net2289),
    .Y(_3446_),
    .A1(_4004_),
    .A2(_3255_));
 sg13g2_nand2_1 _7920_ (.Y(_3447_),
    .A(_3391_),
    .B(_3440_));
 sg13g2_o21ai_1 _7921_ (.B1(_3447_),
    .Y(_3448_),
    .A1(_0086_),
    .A2(_3443_));
 sg13g2_a22oi_1 _7922_ (.Y(_3449_),
    .B1(_3448_),
    .B2(net2289),
    .A2(_3446_),
    .A1(net798));
 sg13g2_inv_1 _7923_ (.Y(_0266_),
    .A(net799));
 sg13g2_or2_1 _7924_ (.X(_3450_),
    .B(_3392_),
    .A(net2261));
 sg13g2_o21ai_1 _7925_ (.B1(net837),
    .Y(_3451_),
    .A1(net798),
    .A2(\new_tiles_counter[0] ));
 sg13g2_and2_1 _7926_ (.A(_3450_),
    .B(_3451_),
    .X(_3452_));
 sg13g2_nand2b_1 _7927_ (.Y(_3453_),
    .B(net2289),
    .A_N(_3442_));
 sg13g2_nand3_1 _7928_ (.B(net1832),
    .C(_3453_),
    .A(net837),
    .Y(_3454_));
 sg13g2_o21ai_1 _7929_ (.B1(_3454_),
    .Y(_0267_),
    .A1(_3441_),
    .A2(_3452_));
 sg13g2_a21oi_1 _7930_ (.A1(\draw_game_inst.new_tiles_counter[2] ),
    .A2(_3392_),
    .Y(_3455_),
    .B1(_3262_));
 sg13g2_o21ai_1 _7931_ (.B1(_3455_),
    .Y(_3456_),
    .A1(\draw_game_inst.new_tiles_counter[2] ),
    .A2(_3450_));
 sg13g2_o21ai_1 _7932_ (.B1(_3456_),
    .Y(_3457_),
    .A1(_4008_),
    .A2(_3443_));
 sg13g2_o21ai_1 _7933_ (.B1(net844),
    .Y(_0268_),
    .A1(net2289),
    .A2(_4005_));
 sg13g2_o21ai_1 _7934_ (.B1(net689),
    .Y(_3458_),
    .A1(\draw_game_inst.new_tiles_counter[2] ),
    .A2(_3450_));
 sg13g2_a22oi_1 _7935_ (.Y(_0269_),
    .B1(net690),
    .B2(_3440_),
    .A2(_3453_),
    .A1(_4006_));
 sg13g2_nor2_1 _7936_ (.A(btn_select_prev),
    .B(_3390_),
    .Y(_3459_));
 sg13g2_o21ai_1 _7937_ (.B1(net2282),
    .Y(_3460_),
    .A1(retro_colors),
    .A2(_3459_));
 sg13g2_a21oi_1 _7938_ (.A1(_3959_),
    .A2(_3459_),
    .Y(_0270_),
    .B1(_3460_));
 sg13g2_and2_1 _7939_ (.A(net2290),
    .B(net1),
    .X(_0271_));
 sg13g2_xor2_1 _7940_ (.B(\btn_up_debounce.button_sync_1 ),
    .A(\btn_up_debounce.debounced ),
    .X(_3461_));
 sg13g2_nor4_1 _7941_ (.A(\btn_up_debounce.debounce_counter[1] ),
    .B(\btn_up_debounce.debounce_counter[0] ),
    .C(\btn_up_debounce.debounce_counter[3] ),
    .D(\btn_up_debounce.debounce_counter[2] ),
    .Y(_3462_));
 sg13g2_nand3_1 _7942_ (.B(\btn_up_debounce.debounce_counter[16] ),
    .C(_3462_),
    .A(\btn_up_debounce.debounce_counter[15] ),
    .Y(_3463_));
 sg13g2_nand4_1 _7943_ (.B(\btn_up_debounce.debounce_counter[12] ),
    .C(\btn_up_debounce.debounce_counter[14] ),
    .A(_3988_),
    .Y(_3464_),
    .D(\btn_up_debounce.debounce_counter[17] ));
 sg13g2_nor4_1 _7944_ (.A(\btn_up_debounce.debounce_counter[9] ),
    .B(net806),
    .C(\btn_up_debounce.debounce_counter[11] ),
    .D(net593),
    .Y(_3465_));
 sg13g2_nor4_1 _7945_ (.A(\btn_up_debounce.debounce_counter[5] ),
    .B(\btn_up_debounce.debounce_counter[6] ),
    .C(_3463_),
    .D(_3464_),
    .Y(_3466_));
 sg13g2_and4_1 _7946_ (.A(net736),
    .B(net725),
    .C(_3465_),
    .D(_3466_),
    .X(_3467_));
 sg13g2_inv_1 _7947_ (.Y(_3468_),
    .A(_3467_));
 sg13g2_nand3_1 _7948_ (.B(_3461_),
    .C(_3468_),
    .A(net2287),
    .Y(_3469_));
 sg13g2_nor2_1 _7949_ (.A(_0504_),
    .B(net1773),
    .Y(_0272_));
 sg13g2_xnor2_1 _7950_ (.Y(_3470_),
    .A(\btn_up_debounce.debounce_counter[1] ),
    .B(net825));
 sg13g2_nor2_1 _7951_ (.A(net1773),
    .B(net826),
    .Y(_0273_));
 sg13g2_and3_1 _7952_ (.X(_3471_),
    .A(\btn_up_debounce.debounce_counter[1] ),
    .B(\btn_up_debounce.debounce_counter[0] ),
    .C(net501));
 sg13g2_a21oi_1 _7953_ (.A1(\btn_up_debounce.debounce_counter[1] ),
    .A2(\btn_up_debounce.debounce_counter[0] ),
    .Y(_3472_),
    .B1(net501));
 sg13g2_nor3_1 _7954_ (.A(net1773),
    .B(_3471_),
    .C(net502),
    .Y(_0274_));
 sg13g2_and2_1 _7955_ (.A(net781),
    .B(_3471_),
    .X(_3473_));
 sg13g2_nor2_1 _7956_ (.A(net781),
    .B(_3471_),
    .Y(_3474_));
 sg13g2_nor3_1 _7957_ (.A(net1773),
    .B(_3473_),
    .C(net782),
    .Y(_0275_));
 sg13g2_and2_1 _7958_ (.A(net736),
    .B(_3473_),
    .X(_3475_));
 sg13g2_nor2_1 _7959_ (.A(net736),
    .B(_3473_),
    .Y(_3476_));
 sg13g2_nor3_1 _7960_ (.A(net1773),
    .B(_3475_),
    .C(net737),
    .Y(_0276_));
 sg13g2_and2_1 _7961_ (.A(net711),
    .B(_3475_),
    .X(_3477_));
 sg13g2_nor2_1 _7962_ (.A(net711),
    .B(_3475_),
    .Y(_3478_));
 sg13g2_nor3_1 _7963_ (.A(net1772),
    .B(_3477_),
    .C(net712),
    .Y(_0277_));
 sg13g2_nor2_1 _7964_ (.A(net731),
    .B(_3477_),
    .Y(_3479_));
 sg13g2_and2_1 _7965_ (.A(net731),
    .B(_3477_),
    .X(_3480_));
 sg13g2_nor3_1 _7966_ (.A(net1772),
    .B(_3479_),
    .C(_3480_),
    .Y(_0278_));
 sg13g2_nor2_1 _7967_ (.A(net725),
    .B(_3480_),
    .Y(_3481_));
 sg13g2_and2_1 _7968_ (.A(net725),
    .B(_3480_),
    .X(_3482_));
 sg13g2_nor3_1 _7969_ (.A(net1772),
    .B(net726),
    .C(_3482_),
    .Y(_0279_));
 sg13g2_nor2_1 _7970_ (.A(net806),
    .B(_3482_),
    .Y(_3483_));
 sg13g2_and2_1 _7971_ (.A(net806),
    .B(_3482_),
    .X(_3484_));
 sg13g2_nor3_1 _7972_ (.A(net1772),
    .B(_3483_),
    .C(_3484_),
    .Y(_0280_));
 sg13g2_xnor2_1 _7973_ (.Y(_3485_),
    .A(net853),
    .B(_3484_));
 sg13g2_nor2_1 _7974_ (.A(net1772),
    .B(_3485_),
    .Y(_0281_));
 sg13g2_a21oi_1 _7975_ (.A1(\btn_up_debounce.debounce_counter[9] ),
    .A2(_3484_),
    .Y(_3486_),
    .B1(net593));
 sg13g2_and3_1 _7976_ (.X(_3487_),
    .A(net853),
    .B(net593),
    .C(_3484_));
 sg13g2_nor3_1 _7977_ (.A(net1772),
    .B(net594),
    .C(_3487_),
    .Y(_0282_));
 sg13g2_xnor2_1 _7978_ (.Y(_3488_),
    .A(net866),
    .B(_3487_));
 sg13g2_nor2_1 _7979_ (.A(net1774),
    .B(_3488_),
    .Y(_0283_));
 sg13g2_a21oi_1 _7980_ (.A1(\btn_up_debounce.debounce_counter[11] ),
    .A2(_3487_),
    .Y(_3489_),
    .B1(net652));
 sg13g2_and3_1 _7981_ (.X(_3490_),
    .A(\btn_up_debounce.debounce_counter[11] ),
    .B(net652),
    .C(_3487_));
 sg13g2_nor3_1 _7982_ (.A(net1772),
    .B(net653),
    .C(_3490_),
    .Y(_0284_));
 sg13g2_nor2_1 _7983_ (.A(net815),
    .B(_3490_),
    .Y(_3491_));
 sg13g2_and2_1 _7984_ (.A(net815),
    .B(_3490_),
    .X(_3492_));
 sg13g2_nor3_1 _7985_ (.A(net1772),
    .B(net816),
    .C(_3492_),
    .Y(_0285_));
 sg13g2_nor2_1 _7986_ (.A(net800),
    .B(_3492_),
    .Y(_3493_));
 sg13g2_and2_1 _7987_ (.A(net800),
    .B(_3492_),
    .X(_3494_));
 sg13g2_nor3_1 _7988_ (.A(net1773),
    .B(net801),
    .C(_3494_),
    .Y(_0286_));
 sg13g2_nor2_1 _7989_ (.A(net734),
    .B(_3494_),
    .Y(_3495_));
 sg13g2_and2_1 _7990_ (.A(net734),
    .B(_3494_),
    .X(_3496_));
 sg13g2_nor3_1 _7991_ (.A(net1774),
    .B(net735),
    .C(_3496_),
    .Y(_0287_));
 sg13g2_nor2_1 _7992_ (.A(net817),
    .B(_3496_),
    .Y(_3497_));
 sg13g2_and2_1 _7993_ (.A(net817),
    .B(_3496_),
    .X(_3498_));
 sg13g2_nor3_1 _7994_ (.A(net1773),
    .B(_3497_),
    .C(_3498_),
    .Y(_0288_));
 sg13g2_nor2_1 _7995_ (.A(net720),
    .B(_3498_),
    .Y(_3499_));
 sg13g2_a21oi_1 _7996_ (.A1(net720),
    .A2(_3498_),
    .Y(_3500_),
    .B1(net1773));
 sg13g2_nor2b_1 _7997_ (.A(net721),
    .B_N(_3500_),
    .Y(_0289_));
 sg13g2_and2_1 _7998_ (.A(net2285),
    .B(net1026),
    .X(_0290_));
 sg13g2_o21ai_1 _7999_ (.B1(net2287),
    .Y(_3501_),
    .A1(\btn_up_debounce.button_sync_1 ),
    .A2(_3468_));
 sg13g2_a21oi_1 _8000_ (.A1(_3958_),
    .A2(_3468_),
    .Y(_0291_),
    .B1(_3501_));
 sg13g2_and2_1 _8001_ (.A(net2290),
    .B(net2),
    .X(_0292_));
 sg13g2_xor2_1 _8002_ (.B(net769),
    .A(\btn_down_debounce.debounced ),
    .X(_3502_));
 sg13g2_nor2_1 _8003_ (.A(\btn_down_debounce.debounce_counter[0] ),
    .B(net871),
    .Y(_3503_));
 sg13g2_nor3_1 _8004_ (.A(\btn_down_debounce.debounce_counter[3] ),
    .B(\btn_down_debounce.debounce_counter[2] ),
    .C(net701),
    .Y(_3504_));
 sg13g2_nand4_1 _8005_ (.B(\btn_down_debounce.debounce_counter[14] ),
    .C(net492),
    .A(\btn_down_debounce.debounce_counter[15] ),
    .Y(_3505_),
    .D(\btn_down_debounce.debounce_counter[16] ));
 sg13g2_nor3_1 _8006_ (.A(\btn_down_debounce.debounce_counter[11] ),
    .B(net601),
    .C(net732),
    .Y(_3506_));
 sg13g2_nand2_1 _8007_ (.Y(_3507_),
    .A(net608),
    .B(_3506_));
 sg13g2_nor4_1 _8008_ (.A(\btn_down_debounce.debounce_counter[6] ),
    .B(_3991_),
    .C(\btn_down_debounce.debounce_counter[9] ),
    .D(_3505_),
    .Y(_3508_));
 sg13g2_nand4_1 _8009_ (.B(_3503_),
    .C(_3504_),
    .A(net699),
    .Y(_3509_),
    .D(_3508_));
 sg13g2_nor3_1 _8010_ (.A(net738),
    .B(_3507_),
    .C(_3509_),
    .Y(_3510_));
 sg13g2_inv_1 _8011_ (.Y(_3511_),
    .A(_3510_));
 sg13g2_nand3_1 _8012_ (.B(_3502_),
    .C(_3511_),
    .A(net2286),
    .Y(_3512_));
 sg13g2_inv_1 _8013_ (.Y(_3513_),
    .A(net1771));
 sg13g2_and2_1 _8014_ (.A(net422),
    .B(_3513_),
    .X(_0293_));
 sg13g2_and2_1 _8015_ (.A(\btn_down_debounce.debounce_counter[0] ),
    .B(net871),
    .X(_3514_));
 sg13g2_nor3_1 _8016_ (.A(net872),
    .B(net1771),
    .C(_3514_),
    .Y(_0294_));
 sg13g2_and2_1 _8017_ (.A(net728),
    .B(_3514_),
    .X(_3515_));
 sg13g2_nor2_1 _8018_ (.A(net728),
    .B(_3514_),
    .Y(_3516_));
 sg13g2_nor3_1 _8019_ (.A(net1771),
    .B(_3515_),
    .C(net729),
    .Y(_0295_));
 sg13g2_and2_1 _8020_ (.A(net708),
    .B(_3515_),
    .X(_3517_));
 sg13g2_nor2_1 _8021_ (.A(net708),
    .B(_3515_),
    .Y(_3518_));
 sg13g2_nor3_1 _8022_ (.A(net1771),
    .B(_3517_),
    .C(net709),
    .Y(_0296_));
 sg13g2_and2_1 _8023_ (.A(net699),
    .B(_3517_),
    .X(_3519_));
 sg13g2_nor2_1 _8024_ (.A(net699),
    .B(_3517_),
    .Y(_3520_));
 sg13g2_nor3_1 _8025_ (.A(net1771),
    .B(_3519_),
    .C(net700),
    .Y(_0297_));
 sg13g2_and2_1 _8026_ (.A(net701),
    .B(_3519_),
    .X(_3521_));
 sg13g2_nor2_1 _8027_ (.A(net701),
    .B(_3519_),
    .Y(_3522_));
 sg13g2_nor3_1 _8028_ (.A(net1771),
    .B(_3521_),
    .C(_3522_),
    .Y(_0298_));
 sg13g2_nor2_1 _8029_ (.A(net807),
    .B(_3521_),
    .Y(_3523_));
 sg13g2_and2_1 _8030_ (.A(net807),
    .B(_3521_),
    .X(_3524_));
 sg13g2_nor3_1 _8031_ (.A(net1771),
    .B(_3523_),
    .C(_3524_),
    .Y(_0299_));
 sg13g2_nor2_1 _8032_ (.A(net822),
    .B(_3524_),
    .Y(_3525_));
 sg13g2_and2_1 _8033_ (.A(net822),
    .B(_3524_),
    .X(_3526_));
 sg13g2_nor3_1 _8034_ (.A(net1770),
    .B(_3525_),
    .C(_3526_),
    .Y(_0300_));
 sg13g2_nor2_1 _8035_ (.A(net738),
    .B(_3526_),
    .Y(_3527_));
 sg13g2_and2_1 _8036_ (.A(net738),
    .B(_3526_),
    .X(_3528_));
 sg13g2_nor3_1 _8037_ (.A(net1770),
    .B(net739),
    .C(_3528_),
    .Y(_0301_));
 sg13g2_xnor2_1 _8038_ (.Y(_3529_),
    .A(net868),
    .B(_3528_));
 sg13g2_nor2_1 _8039_ (.A(net1770),
    .B(_3529_),
    .Y(_0302_));
 sg13g2_a21oi_1 _8040_ (.A1(\btn_down_debounce.debounce_counter[9] ),
    .A2(_3528_),
    .Y(_3530_),
    .B1(net601));
 sg13g2_and3_1 _8041_ (.X(_3531_),
    .A(\btn_down_debounce.debounce_counter[9] ),
    .B(net601),
    .C(_3528_));
 sg13g2_nor3_1 _8042_ (.A(net1770),
    .B(net602),
    .C(_3531_),
    .Y(_0303_));
 sg13g2_xnor2_1 _8043_ (.Y(_3532_),
    .A(net854),
    .B(_3531_));
 sg13g2_nor2_1 _8044_ (.A(net1770),
    .B(net855),
    .Y(_0304_));
 sg13g2_a21oi_1 _8045_ (.A1(\btn_down_debounce.debounce_counter[11] ),
    .A2(_3531_),
    .Y(_3533_),
    .B1(net608));
 sg13g2_and3_1 _8046_ (.X(_3534_),
    .A(\btn_down_debounce.debounce_counter[11] ),
    .B(net608),
    .C(_3531_));
 sg13g2_nor3_1 _8047_ (.A(net1770),
    .B(net609),
    .C(_3534_),
    .Y(_0305_));
 sg13g2_nor2_1 _8048_ (.A(net732),
    .B(_3534_),
    .Y(_3535_));
 sg13g2_and2_1 _8049_ (.A(net732),
    .B(_3534_),
    .X(_3536_));
 sg13g2_nor3_1 _8050_ (.A(net1770),
    .B(net733),
    .C(_3536_),
    .Y(_0306_));
 sg13g2_and2_1 _8051_ (.A(net867),
    .B(_3536_),
    .X(_3537_));
 sg13g2_o21ai_1 _8052_ (.B1(_3513_),
    .Y(_3538_),
    .A1(net867),
    .A2(_3536_));
 sg13g2_nor2_1 _8053_ (.A(_3537_),
    .B(_3538_),
    .Y(_0307_));
 sg13g2_and2_1 _8054_ (.A(net874),
    .B(_3537_),
    .X(_3539_));
 sg13g2_o21ai_1 _8055_ (.B1(_3513_),
    .Y(_3540_),
    .A1(net874),
    .A2(_3537_));
 sg13g2_nor2_1 _8056_ (.A(_3539_),
    .B(_3540_),
    .Y(_0308_));
 sg13g2_o21ai_1 _8057_ (.B1(_3513_),
    .Y(_3541_),
    .A1(net584),
    .A2(_3539_));
 sg13g2_a21oi_1 _8058_ (.A1(net584),
    .A2(_3539_),
    .Y(_0309_),
    .B1(_3541_));
 sg13g2_a21oi_1 _8059_ (.A1(\btn_down_debounce.debounce_counter[16] ),
    .A2(_3539_),
    .Y(_3542_),
    .B1(net492));
 sg13g2_nor2b_1 _8060_ (.A(_3505_),
    .B_N(_3536_),
    .Y(_3543_));
 sg13g2_nor3_1 _8061_ (.A(net1770),
    .B(net493),
    .C(_3543_),
    .Y(_0310_));
 sg13g2_o21ai_1 _8062_ (.B1(net2286),
    .Y(_3544_),
    .A1(net769),
    .A2(_3511_));
 sg13g2_a21oi_1 _8063_ (.A1(_3957_),
    .A2(_3511_),
    .Y(_0311_),
    .B1(_3544_));
 sg13g2_and2_1 _8064_ (.A(net2289),
    .B(net3),
    .X(_0312_));
 sg13g2_xor2_1 _8065_ (.B(\btn_left_debounce.button_sync_1 ),
    .A(\btn_left_debounce.debounced ),
    .X(_3545_));
 sg13g2_nor4_1 _8066_ (.A(\btn_left_debounce.debounce_counter[1] ),
    .B(\btn_left_debounce.debounce_counter[0] ),
    .C(\btn_left_debounce.debounce_counter[3] ),
    .D(net504),
    .Y(_3546_));
 sg13g2_nand2_1 _8067_ (.Y(_3547_),
    .A(\btn_left_debounce.debounce_counter[12] ),
    .B(\btn_left_debounce.debounce_counter[17] ));
 sg13g2_or4_1 _8068_ (.A(\btn_left_debounce.debounce_counter[9] ),
    .B(net821),
    .C(\btn_left_debounce.debounce_counter[11] ),
    .D(net510),
    .X(_3548_));
 sg13g2_nand2_1 _8069_ (.Y(_3549_),
    .A(\btn_left_debounce.debounce_counter[4] ),
    .B(\btn_left_debounce.debounce_counter[7] ));
 sg13g2_nor4_1 _8070_ (.A(net764),
    .B(_3990_),
    .C(_3547_),
    .D(_3549_),
    .Y(_3550_));
 sg13g2_nand4_1 _8071_ (.B(net818),
    .C(_3546_),
    .A(net810),
    .Y(_3551_),
    .D(_3550_));
 sg13g2_nor4_1 _8072_ (.A(net790),
    .B(net762),
    .C(_3548_),
    .D(_3551_),
    .Y(_3552_));
 sg13g2_inv_1 _8073_ (.Y(_3553_),
    .A(_3552_));
 sg13g2_nand3_1 _8074_ (.B(_3545_),
    .C(_3553_),
    .A(net2286),
    .Y(_3554_));
 sg13g2_nor2_1 _8075_ (.A(_0505_),
    .B(net1767),
    .Y(_0313_));
 sg13g2_xnor2_1 _8076_ (.Y(_3555_),
    .A(net862),
    .B(\btn_left_debounce.debounce_counter[0] ));
 sg13g2_nor2_1 _8077_ (.A(net1767),
    .B(net863),
    .Y(_0314_));
 sg13g2_and3_1 _8078_ (.X(_3556_),
    .A(\btn_left_debounce.debounce_counter[1] ),
    .B(\btn_left_debounce.debounce_counter[0] ),
    .C(net504));
 sg13g2_a21oi_1 _8079_ (.A1(\btn_left_debounce.debounce_counter[1] ),
    .A2(\btn_left_debounce.debounce_counter[0] ),
    .Y(_3557_),
    .B1(net504));
 sg13g2_nor3_1 _8080_ (.A(net1767),
    .B(_3556_),
    .C(net505),
    .Y(_0315_));
 sg13g2_and2_1 _8081_ (.A(net740),
    .B(_3556_),
    .X(_3558_));
 sg13g2_nor2_1 _8082_ (.A(net740),
    .B(_3556_),
    .Y(_3559_));
 sg13g2_nor3_1 _8083_ (.A(net1767),
    .B(_3558_),
    .C(net741),
    .Y(_0316_));
 sg13g2_and2_1 _8084_ (.A(net754),
    .B(_3558_),
    .X(_3560_));
 sg13g2_nor2_1 _8085_ (.A(net754),
    .B(_3558_),
    .Y(_3561_));
 sg13g2_nor3_1 _8086_ (.A(net1767),
    .B(_3560_),
    .C(_3561_),
    .Y(_0317_));
 sg13g2_and2_1 _8087_ (.A(net790),
    .B(_3560_),
    .X(_3562_));
 sg13g2_nor2_1 _8088_ (.A(net790),
    .B(_3560_),
    .Y(_3563_));
 sg13g2_nor3_1 _8089_ (.A(net1769),
    .B(_3562_),
    .C(_3563_),
    .Y(_0318_));
 sg13g2_nor2_1 _8090_ (.A(net762),
    .B(_3562_),
    .Y(_3564_));
 sg13g2_and2_1 _8091_ (.A(net762),
    .B(_3562_),
    .X(_3565_));
 sg13g2_nor3_1 _8092_ (.A(net1767),
    .B(net763),
    .C(_3565_),
    .Y(_0319_));
 sg13g2_nor2_1 _8093_ (.A(net780),
    .B(_3565_),
    .Y(_3566_));
 sg13g2_and2_1 _8094_ (.A(net780),
    .B(_3565_),
    .X(_3567_));
 sg13g2_nor3_1 _8095_ (.A(net1767),
    .B(_3566_),
    .C(_3567_),
    .Y(_0320_));
 sg13g2_nor2_1 _8096_ (.A(net821),
    .B(_3567_),
    .Y(_3568_));
 sg13g2_and2_1 _8097_ (.A(net821),
    .B(_3567_),
    .X(_3569_));
 sg13g2_nor3_1 _8098_ (.A(net1767),
    .B(_3568_),
    .C(_3569_),
    .Y(_0321_));
 sg13g2_xnor2_1 _8099_ (.Y(_3570_),
    .A(net846),
    .B(_3569_));
 sg13g2_nor2_1 _8100_ (.A(net1769),
    .B(_3570_),
    .Y(_0322_));
 sg13g2_a21oi_1 _8101_ (.A1(\btn_left_debounce.debounce_counter[9] ),
    .A2(_3569_),
    .Y(_3571_),
    .B1(net510));
 sg13g2_and3_1 _8102_ (.X(_3572_),
    .A(\btn_left_debounce.debounce_counter[9] ),
    .B(net510),
    .C(_3569_));
 sg13g2_nor3_1 _8103_ (.A(net1768),
    .B(net511),
    .C(_3572_),
    .Y(_0323_));
 sg13g2_xnor2_1 _8104_ (.Y(_3573_),
    .A(net839),
    .B(_3572_));
 sg13g2_nor2_1 _8105_ (.A(net1768),
    .B(net840),
    .Y(_0324_));
 sg13g2_a21oi_1 _8106_ (.A1(\btn_left_debounce.debounce_counter[11] ),
    .A2(_3572_),
    .Y(_3574_),
    .B1(net627));
 sg13g2_and3_1 _8107_ (.X(_3575_),
    .A(\btn_left_debounce.debounce_counter[11] ),
    .B(net627),
    .C(_3572_));
 sg13g2_nor3_1 _8108_ (.A(net1768),
    .B(net628),
    .C(_3575_),
    .Y(_0325_));
 sg13g2_nor2_1 _8109_ (.A(net764),
    .B(_3575_),
    .Y(_3576_));
 sg13g2_and2_1 _8110_ (.A(net764),
    .B(_3575_),
    .X(_3577_));
 sg13g2_nor3_1 _8111_ (.A(net1768),
    .B(net765),
    .C(_3577_),
    .Y(_0326_));
 sg13g2_nor2_1 _8112_ (.A(net784),
    .B(_3577_),
    .Y(_3578_));
 sg13g2_and2_1 _8113_ (.A(net784),
    .B(_3577_),
    .X(_3579_));
 sg13g2_nor3_1 _8114_ (.A(net1768),
    .B(_3578_),
    .C(_3579_),
    .Y(_0327_));
 sg13g2_nor2_1 _8115_ (.A(net810),
    .B(_3579_),
    .Y(_3580_));
 sg13g2_and2_1 _8116_ (.A(net810),
    .B(_3579_),
    .X(_3581_));
 sg13g2_nor3_1 _8117_ (.A(net1768),
    .B(_3580_),
    .C(_3581_),
    .Y(_0328_));
 sg13g2_nor2_1 _8118_ (.A(net818),
    .B(_3581_),
    .Y(_3582_));
 sg13g2_and2_1 _8119_ (.A(net818),
    .B(_3581_),
    .X(_3583_));
 sg13g2_nor3_1 _8120_ (.A(net1768),
    .B(_3582_),
    .C(_3583_),
    .Y(_0329_));
 sg13g2_nor2_1 _8121_ (.A(net742),
    .B(_3583_),
    .Y(_3584_));
 sg13g2_a21oi_1 _8122_ (.A1(net742),
    .A2(_3583_),
    .Y(_3585_),
    .B1(net1768));
 sg13g2_nor2b_1 _8123_ (.A(net743),
    .B_N(_3585_),
    .Y(_0330_));
 sg13g2_and2_1 _8124_ (.A(net2287),
    .B(net509),
    .X(_0331_));
 sg13g2_o21ai_1 _8125_ (.B1(net2286),
    .Y(_3586_),
    .A1(\btn_left_debounce.button_sync_1 ),
    .A2(_3553_));
 sg13g2_a21oi_1 _8126_ (.A1(_3956_),
    .A2(_3553_),
    .Y(_0332_),
    .B1(_3586_));
 sg13g2_and2_1 _8127_ (.A(net2277),
    .B(net4),
    .X(_0333_));
 sg13g2_xor2_1 _8128_ (.B(\btn_right_debounce.button_sync_1 ),
    .A(net685),
    .X(_3587_));
 sg13g2_nor4_1 _8129_ (.A(\btn_right_debounce.debounce_counter[1] ),
    .B(\btn_right_debounce.debounce_counter[0] ),
    .C(\btn_right_debounce.debounce_counter[3] ),
    .D(\btn_right_debounce.debounce_counter[2] ),
    .Y(_3588_));
 sg13g2_nand3_1 _8130_ (.B(\btn_right_debounce.debounce_counter[16] ),
    .C(_3588_),
    .A(\btn_right_debounce.debounce_counter[15] ),
    .Y(_3589_));
 sg13g2_nand4_1 _8131_ (.B(\btn_right_debounce.debounce_counter[12] ),
    .C(\btn_right_debounce.debounce_counter[14] ),
    .A(_3989_),
    .Y(_3590_),
    .D(\btn_right_debounce.debounce_counter[17] ));
 sg13g2_nor4_1 _8132_ (.A(\btn_right_debounce.debounce_counter[9] ),
    .B(\btn_right_debounce.debounce_counter[8] ),
    .C(\btn_right_debounce.debounce_counter[11] ),
    .D(net566),
    .Y(_3591_));
 sg13g2_nor4_1 _8133_ (.A(\btn_right_debounce.debounce_counter[5] ),
    .B(\btn_right_debounce.debounce_counter[6] ),
    .C(_3589_),
    .D(_3590_),
    .Y(_3592_));
 sg13g2_and4_1 _8134_ (.A(\btn_right_debounce.debounce_counter[4] ),
    .B(\btn_right_debounce.debounce_counter[7] ),
    .C(_3591_),
    .D(_3592_),
    .X(_3593_));
 sg13g2_inv_1 _8135_ (.Y(_3594_),
    .A(_3593_));
 sg13g2_nand3_1 _8136_ (.B(_3587_),
    .C(_3594_),
    .A(net2286),
    .Y(_3595_));
 sg13g2_inv_1 _8137_ (.Y(_3596_),
    .A(net1766));
 sg13g2_and2_1 _8138_ (.A(net423),
    .B(_3596_),
    .X(_0334_));
 sg13g2_xnor2_1 _8139_ (.Y(_3597_),
    .A(\btn_right_debounce.debounce_counter[1] ),
    .B(net831));
 sg13g2_nor2_1 _8140_ (.A(net1766),
    .B(net832),
    .Y(_0335_));
 sg13g2_and3_1 _8141_ (.X(_3598_),
    .A(\btn_right_debounce.debounce_counter[1] ),
    .B(\btn_right_debounce.debounce_counter[0] ),
    .C(net581));
 sg13g2_a21oi_1 _8142_ (.A1(\btn_right_debounce.debounce_counter[1] ),
    .A2(\btn_right_debounce.debounce_counter[0] ),
    .Y(_3599_),
    .B1(net581));
 sg13g2_nor3_1 _8143_ (.A(net1766),
    .B(_3598_),
    .C(net582),
    .Y(_0336_));
 sg13g2_and2_1 _8144_ (.A(net787),
    .B(_3598_),
    .X(_3600_));
 sg13g2_nor2_1 _8145_ (.A(net787),
    .B(_3598_),
    .Y(_3601_));
 sg13g2_nor3_1 _8146_ (.A(net1766),
    .B(_3600_),
    .C(net788),
    .Y(_0337_));
 sg13g2_and2_1 _8147_ (.A(net750),
    .B(_3600_),
    .X(_3602_));
 sg13g2_nor2_1 _8148_ (.A(net750),
    .B(_3600_),
    .Y(_3603_));
 sg13g2_nor3_1 _8149_ (.A(net1766),
    .B(_3602_),
    .C(net751),
    .Y(_0338_));
 sg13g2_and2_1 _8150_ (.A(net760),
    .B(_3602_),
    .X(_3604_));
 sg13g2_nor2_1 _8151_ (.A(net760),
    .B(_3602_),
    .Y(_3605_));
 sg13g2_nor3_1 _8152_ (.A(net1766),
    .B(_3604_),
    .C(_3605_),
    .Y(_0339_));
 sg13g2_nor2_1 _8153_ (.A(net747),
    .B(_3604_),
    .Y(_3606_));
 sg13g2_and2_1 _8154_ (.A(net747),
    .B(_3604_),
    .X(_3607_));
 sg13g2_nor3_1 _8155_ (.A(net1766),
    .B(net748),
    .C(_3607_),
    .Y(_0340_));
 sg13g2_nor2_1 _8156_ (.A(net811),
    .B(_3607_),
    .Y(_3608_));
 sg13g2_and2_1 _8157_ (.A(net811),
    .B(_3607_),
    .X(_3609_));
 sg13g2_nor3_1 _8158_ (.A(net1765),
    .B(_3608_),
    .C(_3609_),
    .Y(_0341_));
 sg13g2_nor2_1 _8159_ (.A(net808),
    .B(_3609_),
    .Y(_3610_));
 sg13g2_and2_1 _8160_ (.A(net808),
    .B(_3609_),
    .X(_3611_));
 sg13g2_nor3_1 _8161_ (.A(net1765),
    .B(net809),
    .C(_3611_),
    .Y(_0342_));
 sg13g2_xnor2_1 _8162_ (.Y(_3612_),
    .A(net875),
    .B(_3611_));
 sg13g2_nor2_1 _8163_ (.A(net1765),
    .B(_3612_),
    .Y(_0343_));
 sg13g2_a21oi_1 _8164_ (.A1(\btn_right_debounce.debounce_counter[9] ),
    .A2(_3611_),
    .Y(_3613_),
    .B1(net566));
 sg13g2_and3_1 _8165_ (.X(_3614_),
    .A(\btn_right_debounce.debounce_counter[9] ),
    .B(net566),
    .C(_3611_));
 sg13g2_nor3_1 _8166_ (.A(net1765),
    .B(net567),
    .C(_3614_),
    .Y(_0344_));
 sg13g2_xnor2_1 _8167_ (.Y(_3615_),
    .A(net849),
    .B(_3614_));
 sg13g2_nor2_1 _8168_ (.A(net1765),
    .B(net850),
    .Y(_0345_));
 sg13g2_a21oi_1 _8169_ (.A1(\btn_right_debounce.debounce_counter[11] ),
    .A2(_3614_),
    .Y(_3616_),
    .B1(net670));
 sg13g2_and3_1 _8170_ (.X(_3617_),
    .A(\btn_right_debounce.debounce_counter[11] ),
    .B(net670),
    .C(_3614_));
 sg13g2_nor3_1 _8171_ (.A(net1765),
    .B(net671),
    .C(_3617_),
    .Y(_0346_));
 sg13g2_nor2_1 _8172_ (.A(net775),
    .B(_3617_),
    .Y(_3618_));
 sg13g2_and2_1 _8173_ (.A(net775),
    .B(_3617_),
    .X(_3619_));
 sg13g2_nor3_1 _8174_ (.A(net1765),
    .B(net776),
    .C(_3619_),
    .Y(_0347_));
 sg13g2_and2_1 _8175_ (.A(net889),
    .B(_3619_),
    .X(_3620_));
 sg13g2_o21ai_1 _8176_ (.B1(_3596_),
    .Y(_3621_),
    .A1(net889),
    .A2(_3619_));
 sg13g2_nor2_1 _8177_ (.A(_3620_),
    .B(_3621_),
    .Y(_0348_));
 sg13g2_o21ai_1 _8178_ (.B1(_3596_),
    .Y(_3622_),
    .A1(net687),
    .A2(_3620_));
 sg13g2_a21oi_1 _8179_ (.A1(net687),
    .A2(_3620_),
    .Y(_0349_),
    .B1(_3622_));
 sg13g2_a21oi_1 _8180_ (.A1(\btn_right_debounce.debounce_counter[15] ),
    .A2(_3620_),
    .Y(_3623_),
    .B1(net588));
 sg13g2_and3_1 _8181_ (.X(_3624_),
    .A(\btn_right_debounce.debounce_counter[15] ),
    .B(net588),
    .C(_3620_));
 sg13g2_nor3_1 _8182_ (.A(net1765),
    .B(net589),
    .C(_3624_),
    .Y(_0350_));
 sg13g2_o21ai_1 _8183_ (.B1(_3596_),
    .Y(_3625_),
    .A1(net460),
    .A2(_3624_));
 sg13g2_a21oi_1 _8184_ (.A1(net460),
    .A2(_3624_),
    .Y(_0351_),
    .B1(_3625_));
 sg13g2_and2_1 _8185_ (.A(net2286),
    .B(net1013),
    .X(_0352_));
 sg13g2_o21ai_1 _8186_ (.B1(net2286),
    .Y(_3626_),
    .A1(\btn_right_debounce.button_sync_1 ),
    .A2(_3594_));
 sg13g2_a21oi_1 _8187_ (.A1(_3955_),
    .A2(_3594_),
    .Y(_0353_),
    .B1(_3626_));
 sg13g2_and2_1 _8188_ (.A(net2268),
    .B(_0519_),
    .X(_0354_));
 sg13g2_nor2b_1 _8189_ (.A(net783),
    .B_N(net416),
    .Y(_3627_));
 sg13g2_nor2_1 _8190_ (.A(net2259),
    .B(net1923),
    .Y(_3628_));
 sg13g2_a22oi_1 _8191_ (.Y(_0355_),
    .B1(net1820),
    .B2(_3953_),
    .A2(net1923),
    .A1(_3954_));
 sg13g2_a22oi_1 _8192_ (.Y(_0356_),
    .B1(net1820),
    .B2(_3952_),
    .A2(net1922),
    .A1(_3953_));
 sg13g2_a22oi_1 _8193_ (.Y(_0357_),
    .B1(net1820),
    .B2(_3951_),
    .A2(net1922),
    .A1(_3952_));
 sg13g2_a22oi_1 _8194_ (.Y(_0358_),
    .B1(net1820),
    .B2(_3950_),
    .A2(net1922),
    .A1(_3951_));
 sg13g2_a22oi_1 _8195_ (.Y(_0359_),
    .B1(net1820),
    .B2(_3949_),
    .A2(net1922),
    .A1(_3950_));
 sg13g2_a22oi_1 _8196_ (.Y(_0360_),
    .B1(net1820),
    .B2(_3948_),
    .A2(net1922),
    .A1(_3949_));
 sg13g2_a22oi_1 _8197_ (.Y(_0361_),
    .B1(net1820),
    .B2(_3947_),
    .A2(net1922),
    .A1(_3948_));
 sg13g2_a22oi_1 _8198_ (.Y(_0362_),
    .B1(net1820),
    .B2(_3946_),
    .A2(net1922),
    .A1(_3947_));
 sg13g2_a22oi_1 _8199_ (.Y(_0363_),
    .B1(net1821),
    .B2(_3945_),
    .A2(net1923),
    .A1(_3946_));
 sg13g2_a22oi_1 _8200_ (.Y(_0364_),
    .B1(net1821),
    .B2(_3944_),
    .A2(net1923),
    .A1(_3945_));
 sg13g2_a22oi_1 _8201_ (.Y(_0365_),
    .B1(net1821),
    .B2(_3943_),
    .A2(net1922),
    .A1(_3944_));
 sg13g2_a22oi_1 _8202_ (.Y(_0366_),
    .B1(net1821),
    .B2(_3942_),
    .A2(net1923),
    .A1(_3943_));
 sg13g2_and2_1 _8203_ (.A(net2277),
    .B(net7),
    .X(_0367_));
 sg13g2_and2_1 _8204_ (.A(net2286),
    .B(net988),
    .X(_0368_));
 sg13g2_and2_1 _8205_ (.A(net2283),
    .B(net6),
    .X(_0369_));
 sg13g2_and2_1 _8206_ (.A(net2282),
    .B(net421),
    .X(_0370_));
 sg13g2_xor2_1 _8207_ (.B(net459),
    .A(net757),
    .X(_3629_));
 sg13g2_xor2_1 _8208_ (.B(net684),
    .A(net927),
    .X(_3630_));
 sg13g2_o21ai_1 _8209_ (.B1(net2270),
    .Y(_3631_),
    .A1(_3629_),
    .A2(_3630_));
 sg13g2_a21oi_1 _8210_ (.A1(_3629_),
    .A2(_3630_),
    .Y(_0371_),
    .B1(_3631_));
 sg13g2_nand2b_1 _8211_ (.Y(_0372_),
    .B(net2268),
    .A_N(net684));
 sg13g2_and2_1 _8212_ (.A(net2265),
    .B(net757),
    .X(_0373_));
 sg13g2_nand2b_1 _8213_ (.Y(_0374_),
    .B(net2264),
    .A_N(net444));
 sg13g2_nand2b_1 _8214_ (.Y(_0375_),
    .B(net2267),
    .A_N(net453));
 sg13g2_nand2b_1 _8215_ (.Y(_0376_),
    .B(net2267),
    .A_N(net448));
 sg13g2_nand2b_1 _8216_ (.Y(_0377_),
    .B(net2264),
    .A_N(net475));
 sg13g2_nand2b_1 _8217_ (.Y(_0378_),
    .B(net2265),
    .A_N(net455));
 sg13g2_and2_1 _8218_ (.A(net2265),
    .B(net458),
    .X(_0379_));
 sg13g2_nand2b_1 _8219_ (.Y(_0380_),
    .B(net2267),
    .A_N(net454));
 sg13g2_and2_1 _8220_ (.A(net2267),
    .B(net456),
    .X(_0381_));
 sg13g2_nand2b_1 _8221_ (.Y(_0382_),
    .B(net2264),
    .A_N(net437));
 sg13g2_nand2b_1 _8222_ (.Y(_0383_),
    .B(net2267),
    .A_N(net476));
 sg13g2_nand2b_1 _8223_ (.Y(_0384_),
    .B(net2267),
    .A_N(net462));
 sg13g2_nand2b_1 _8224_ (.Y(_0385_),
    .B(net2267),
    .A_N(net547));
 sg13g2_nand2b_1 _8225_ (.Y(_0386_),
    .B(net2264),
    .A_N(net457));
 sg13g2_and2_1 _8226_ (.A(net2264),
    .B(net479),
    .X(_0387_));
 sg13g2_and2_1 _8227_ (.A(net2264),
    .B(net428),
    .X(_0388_));
 sg13g2_and2_1 _8228_ (.A(net2264),
    .B(net445),
    .X(_0389_));
 sg13g2_nand2b_1 _8229_ (.Y(_0390_),
    .B(net2265),
    .A_N(net435));
 sg13g2_and2_1 _8230_ (.A(net2267),
    .B(net429),
    .X(_0391_));
 sg13g2_and2_1 _8231_ (.A(net2268),
    .B(net426),
    .X(_0392_));
 sg13g2_nand2b_1 _8232_ (.Y(_0393_),
    .B(net2270),
    .A_N(net459));
 sg13g2_and2_1 _8233_ (.A(net2270),
    .B(net427),
    .X(_0394_));
 sg13g2_and2_1 _8234_ (.A(net2270),
    .B(net431),
    .X(_0395_));
 sg13g2_and2_1 _8235_ (.A(net2270),
    .B(net443),
    .X(_0396_));
 sg13g2_and2_1 _8236_ (.A(net2270),
    .B(net430),
    .X(_0397_));
 sg13g2_and2_1 _8237_ (.A(net2270),
    .B(net425),
    .X(_0398_));
 sg13g2_and2_1 _8238_ (.A(net2271),
    .B(net436),
    .X(_0399_));
 sg13g2_nand2b_1 _8239_ (.Y(_0400_),
    .B(net2271),
    .A_N(net2253));
 sg13g2_and2_1 _8240_ (.A(net2252),
    .B(net2271),
    .X(_0401_));
 sg13g2_nor2_1 _8241_ (.A(_3961_),
    .B(net2259),
    .Y(_0402_));
 sg13g2_nand3_1 _8242_ (.B(net945),
    .C(_1426_),
    .A(net2122),
    .Y(_3632_));
 sg13g2_nor3_2 _8243_ (.A(net1958),
    .B(_3216_),
    .C(_3632_),
    .Y(_3633_));
 sg13g2_nor2_2 _8244_ (.A(net2263),
    .B(_3633_),
    .Y(_3634_));
 sg13g2_nand2b_2 _8245_ (.Y(_3635_),
    .B(net2290),
    .A_N(_3633_));
 sg13g2_nor4_1 _8246_ (.A(_3992_),
    .B(\draw_game_inst.y[8] ),
    .C(net2152),
    .D(net2154),
    .Y(_3636_));
 sg13g2_nand3_1 _8247_ (.B(net1852),
    .C(_3636_),
    .A(_1414_),
    .Y(_3637_));
 sg13g2_nand2_1 _8248_ (.Y(_3638_),
    .A(net2288),
    .B(_3637_));
 sg13g2_inv_1 _8249_ (.Y(_3639_),
    .A(_3638_));
 sg13g2_nand2_2 _8250_ (.Y(_3640_),
    .A(_3633_),
    .B(_3639_));
 sg13g2_inv_1 _8251_ (.Y(_3641_),
    .A(_3640_));
 sg13g2_a22oi_1 _8252_ (.Y(_3642_),
    .B1(_3641_),
    .B2(net2225),
    .A2(_3634_),
    .A1(net2228));
 sg13g2_inv_1 _8253_ (.Y(_0403_),
    .A(_3642_));
 sg13g2_nand2_1 _8254_ (.Y(_3643_),
    .A(net2200),
    .B(_3634_));
 sg13g2_o21ai_1 _8255_ (.B1(_3643_),
    .Y(_0404_),
    .A1(_2662_),
    .A2(_3640_));
 sg13g2_a22oi_1 _8256_ (.Y(_3644_),
    .B1(_3641_),
    .B2(_2451_),
    .A2(_3634_),
    .A1(net2190));
 sg13g2_nor2_1 _8257_ (.A(_1963_),
    .B(_3644_),
    .Y(_0405_));
 sg13g2_nand2_1 _8258_ (.Y(_3645_),
    .A(net2166),
    .B(net1784));
 sg13g2_nor2_1 _8259_ (.A(net2183),
    .B(net1959),
    .Y(_3646_));
 sg13g2_xnor2_1 _8260_ (.Y(_3647_),
    .A(net2166),
    .B(_3646_));
 sg13g2_o21ai_1 _8261_ (.B1(_3645_),
    .Y(_0406_),
    .A1(_3640_),
    .A2(_3647_));
 sg13g2_nor2_1 _8262_ (.A(_1632_),
    .B(net1784),
    .Y(_3648_));
 sg13g2_nor2_1 _8263_ (.A(net1784),
    .B(_3639_),
    .Y(_3649_));
 sg13g2_xnor2_1 _8264_ (.Y(_3650_),
    .A(net2162),
    .B(_3648_));
 sg13g2_nor2_1 _8265_ (.A(_3649_),
    .B(_3650_),
    .Y(_0407_));
 sg13g2_nand2_1 _8266_ (.Y(_3651_),
    .A(net2155),
    .B(net1784));
 sg13g2_nor2_1 _8267_ (.A(net2161),
    .B(_1632_),
    .Y(_3652_));
 sg13g2_xnor2_1 _8268_ (.Y(_3653_),
    .A(net2155),
    .B(_3652_));
 sg13g2_o21ai_1 _8269_ (.B1(_3651_),
    .Y(_0408_),
    .A1(_3640_),
    .A2(_3653_));
 sg13g2_a21oi_1 _8270_ (.A1(_3214_),
    .A2(_3635_),
    .Y(_3654_),
    .B1(net753));
 sg13g2_nor4_2 _8271_ (.A(_3993_),
    .B(net1949),
    .C(_1632_),
    .Y(_3655_),
    .D(net1784));
 sg13g2_nor3_1 _8272_ (.A(_3649_),
    .B(_3654_),
    .C(_3655_),
    .Y(_0409_));
 sg13g2_nand2_1 _8273_ (.Y(_3656_),
    .A(net2152),
    .B(net1784));
 sg13g2_nor3_1 _8274_ (.A(net848),
    .B(net1949),
    .C(_1632_),
    .Y(_3657_));
 sg13g2_xnor2_1 _8275_ (.Y(_3658_),
    .A(net2152),
    .B(_3657_));
 sg13g2_o21ai_1 _8276_ (.B1(_3656_),
    .Y(_0410_),
    .A1(_3640_),
    .A2(_3658_));
 sg13g2_nand3_1 _8277_ (.B(net2152),
    .C(_3655_),
    .A(net883),
    .Y(_3659_));
 sg13g2_nand2b_1 _8278_ (.Y(_3660_),
    .B(_3659_),
    .A_N(_3649_));
 sg13g2_a21oi_1 _8279_ (.A1(net2152),
    .A2(_3655_),
    .Y(_3661_),
    .B1(net883));
 sg13g2_nor2_1 _8280_ (.A(_3660_),
    .B(_3661_),
    .Y(_0411_));
 sg13g2_a22oi_1 _8281_ (.Y(_0412_),
    .B1(_3660_),
    .B2(_1407_),
    .A2(_3659_),
    .A1(_3992_));
 sg13g2_and2_1 _8282_ (.A(net2282),
    .B(net5),
    .X(_0413_));
 sg13g2_and2_1 _8283_ (.A(net2287),
    .B(net434),
    .X(_0414_));
 sg13g2_nor2b_1 _8284_ (.A(\gamepad_pmod.driver.pmod_latch_prev ),
    .B_N(net417),
    .Y(_3662_));
 sg13g2_nor2_1 _8285_ (.A(net2259),
    .B(net1920),
    .Y(_3663_));
 sg13g2_a22oi_1 _8286_ (.Y(_0415_),
    .B1(net1819),
    .B2(_3965_),
    .A2(net1921),
    .A1(_3953_));
 sg13g2_a22oi_1 _8287_ (.Y(_0416_),
    .B1(net1819),
    .B2(_3964_),
    .A2(net1921),
    .A1(_3952_));
 sg13g2_a22oi_1 _8288_ (.Y(_0417_),
    .B1(net1819),
    .B2(_3967_),
    .A2(net1921),
    .A1(_3951_));
 sg13g2_a22oi_1 _8289_ (.Y(_0418_),
    .B1(net1819),
    .B2(_3966_),
    .A2(net1921),
    .A1(_3950_));
 sg13g2_a22oi_1 _8290_ (.Y(_0419_),
    .B1(net1818),
    .B2(_3969_),
    .A2(net1920),
    .A1(_3949_));
 sg13g2_a22oi_1 _8291_ (.Y(_0420_),
    .B1(net1818),
    .B2(_3968_),
    .A2(net1920),
    .A1(_3948_));
 sg13g2_a22oi_1 _8292_ (.Y(_0421_),
    .B1(net1818),
    .B2(_3971_),
    .A2(net1920),
    .A1(_3947_));
 sg13g2_a22oi_1 _8293_ (.Y(_0422_),
    .B1(net1818),
    .B2(_3970_),
    .A2(net1920),
    .A1(_3946_));
 sg13g2_a22oi_1 _8294_ (.Y(_0423_),
    .B1(net1818),
    .B2(_3973_),
    .A2(net1920),
    .A1(_3945_));
 sg13g2_a22oi_1 _8295_ (.Y(_0424_),
    .B1(net1818),
    .B2(_3972_),
    .A2(net1921),
    .A1(_3944_));
 sg13g2_a22oi_1 _8296_ (.Y(_0425_),
    .B1(net1818),
    .B2(_3975_),
    .A2(net1920),
    .A1(_3943_));
 sg13g2_a22oi_1 _8297_ (.Y(_0426_),
    .B1(net1818),
    .B2(_3974_),
    .A2(net1920),
    .A1(_3942_));
 sg13g2_and2_1 _8298_ (.A(net418),
    .B(net1784),
    .X(_0427_));
 sg13g2_a21oi_1 _8299_ (.A1(_2226_),
    .A2(_2507_),
    .Y(_0428_),
    .B1(_3635_));
 sg13g2_nand2_1 _8300_ (.Y(_3664_),
    .A(net2291),
    .B(_3215_));
 sg13g2_a21oi_1 _8301_ (.A1(_4000_),
    .A2(_2916_),
    .Y(_0429_),
    .B1(_3664_));
 sg13g2_nand2_1 _8302_ (.Y(_3665_),
    .A(net2290),
    .B(_3216_));
 sg13g2_a21oi_1 _8303_ (.A1(net2028),
    .A2(net996),
    .Y(_0430_),
    .B1(_3665_));
 sg13g2_xnor2_1 _8304_ (.Y(_3666_),
    .A(net2023),
    .B(_3216_));
 sg13g2_nor2_1 _8305_ (.A(_3635_),
    .B(_3666_),
    .Y(_0431_));
 sg13g2_nor2_1 _8306_ (.A(_2492_),
    .B(_3215_),
    .Y(_3667_));
 sg13g2_xnor2_1 _8307_ (.Y(_3668_),
    .A(net2135),
    .B(_3667_));
 sg13g2_nor2_1 _8308_ (.A(_3635_),
    .B(_3668_),
    .Y(_0432_));
 sg13g2_o21ai_1 _8309_ (.B1(net1784),
    .Y(_3669_),
    .A1(net2128),
    .A2(_3217_));
 sg13g2_a21oi_1 _8310_ (.A1(net2128),
    .A2(_3217_),
    .Y(_0433_),
    .B1(_3669_));
 sg13g2_a21oi_1 _8311_ (.A1(net2129),
    .A2(_3217_),
    .Y(_3670_),
    .B1(net2123));
 sg13g2_and2_1 _8312_ (.A(net1979),
    .B(_3217_),
    .X(_3671_));
 sg13g2_nor3_1 _8313_ (.A(_3635_),
    .B(_3670_),
    .C(_3671_),
    .Y(_0434_));
 sg13g2_a21oi_1 _8314_ (.A1(net1979),
    .A2(_3217_),
    .Y(_3672_),
    .B1(net2122));
 sg13g2_and3_1 _8315_ (.X(_3673_),
    .A(net2122),
    .B(net1979),
    .C(_3217_));
 sg13g2_nor3_1 _8316_ (.A(_3635_),
    .B(_3672_),
    .C(_3673_),
    .Y(_0435_));
 sg13g2_xnor2_1 _8317_ (.Y(_3674_),
    .A(net945),
    .B(_3673_));
 sg13g2_nor2_1 _8318_ (.A(_3635_),
    .B(_3674_),
    .Y(_0436_));
 sg13g2_nand4_1 _8319_ (.B(\welcome_screen_inst.welcome_counter[3] ),
    .C(net804),
    .A(net834),
    .Y(_3675_),
    .D(net802));
 sg13g2_or2_1 _8320_ (.X(_3676_),
    .B(_3675_),
    .A(\welcome_screen_inst.welcome_counter[0] ));
 sg13g2_nand2_1 _8321_ (.Y(_3677_),
    .A(_3254_),
    .B(_3676_));
 sg13g2_nor2b_2 _8322_ (.A(net2252),
    .B_N(\lfsr_inst.lfsr[28] ),
    .Y(_3678_));
 sg13g2_nand2b_1 _8323_ (.Y(_3679_),
    .B(net2253),
    .A_N(\lfsr_inst.lfsr[29] ));
 sg13g2_nor2b_2 _8324_ (.A(net2253),
    .B_N(net2252),
    .Y(_3680_));
 sg13g2_nand2b_1 _8325_ (.Y(_3681_),
    .B(net2252),
    .A_N(net2253));
 sg13g2_nand2_1 _8326_ (.Y(_3682_),
    .A(\welcome_screen_grid[56] ),
    .B(_3680_));
 sg13g2_nor2_2 _8327_ (.A(net2252),
    .B(net2253),
    .Y(_3683_));
 sg13g2_or2_1 _8328_ (.X(_3684_),
    .B(net2253),
    .A(net2252));
 sg13g2_and2_2 _8329_ (.A(net2252),
    .B(net2253),
    .X(_3685_));
 sg13g2_nand2_1 _8330_ (.Y(_3686_),
    .A(net2252),
    .B(net2253));
 sg13g2_a21oi_1 _8331_ (.A1(\welcome_screen_grid[48] ),
    .A2(_3683_),
    .Y(_3687_),
    .B1(_3961_));
 sg13g2_a22oi_1 _8332_ (.Y(_3688_),
    .B1(_3685_),
    .B2(\welcome_screen_grid[60] ),
    .A2(_3678_),
    .A1(\welcome_screen_grid[52] ));
 sg13g2_nand3_1 _8333_ (.B(_3687_),
    .C(_3688_),
    .A(_3682_),
    .Y(_3689_));
 sg13g2_a22oi_1 _8334_ (.Y(_3690_),
    .B1(_3685_),
    .B2(\welcome_screen_grid[44] ),
    .A2(_3683_),
    .A1(\welcome_screen_grid[32] ));
 sg13g2_a221oi_1 _8335_ (.B2(\welcome_screen_grid[40] ),
    .C1(\lfsr_inst.lfsr[30] ),
    .B1(_3680_),
    .A1(\welcome_screen_grid[36] ),
    .Y(_3691_),
    .A2(_3678_));
 sg13g2_a21oi_1 _8336_ (.A1(_3690_),
    .A2(_3691_),
    .Y(_3692_),
    .B1(_3962_));
 sg13g2_nand2_1 _8337_ (.Y(_3693_),
    .A(\welcome_screen_grid[11] ),
    .B(_3680_));
 sg13g2_a21oi_1 _8338_ (.A1(\welcome_screen_grid[12] ),
    .A2(_3685_),
    .Y(_3694_),
    .B1(\lfsr_inst.lfsr[30] ));
 sg13g2_a22oi_1 _8339_ (.Y(_3695_),
    .B1(_3683_),
    .B2(\welcome_screen_grid[0] ),
    .A2(_3678_),
    .A1(\welcome_screen_grid[4] ));
 sg13g2_nand3_1 _8340_ (.B(_3694_),
    .C(_3695_),
    .A(_3693_),
    .Y(_3696_));
 sg13g2_a22oi_1 _8341_ (.Y(_3697_),
    .B1(_3680_),
    .B2(\welcome_screen_grid[24] ),
    .A2(_3678_),
    .A1(\welcome_screen_grid[20] ));
 sg13g2_a221oi_1 _8342_ (.B2(\welcome_screen_grid[28] ),
    .C1(_3961_),
    .B1(_3685_),
    .A1(\welcome_screen_grid[16] ),
    .Y(_3698_),
    .A2(_3683_));
 sg13g2_a21oi_1 _8343_ (.A1(_3697_),
    .A2(_3698_),
    .Y(_3699_),
    .B1(\lfsr_inst.lfsr[31] ));
 sg13g2_a221oi_1 _8344_ (.B2(_3699_),
    .C1(_3676_),
    .B1(_3696_),
    .A1(_3689_),
    .Y(_3700_),
    .A2(_3692_));
 sg13g2_a21o_2 _8345_ (.A2(_3676_),
    .A1(_3254_),
    .B1(_3700_),
    .X(_3701_));
 sg13g2_nor2b_1 _8346_ (.A(_3675_),
    .B_N(_3701_),
    .Y(_3702_));
 sg13g2_nand2_1 _8347_ (.Y(_3703_),
    .A(net1014),
    .B(_3701_));
 sg13g2_nor2b_1 _8348_ (.A(_3702_),
    .B_N(_3703_),
    .Y(_3704_));
 sg13g2_or2_1 _8349_ (.X(_3705_),
    .B(_3701_),
    .A(net1014));
 sg13g2_and3_1 _8350_ (.X(_0437_),
    .A(net2285),
    .B(_3704_),
    .C(_3705_));
 sg13g2_a21oi_1 _8351_ (.A1(net802),
    .A2(_3704_),
    .Y(_3706_),
    .B1(net2259));
 sg13g2_o21ai_1 _8352_ (.B1(_3706_),
    .Y(_0438_),
    .A1(net802),
    .A2(_3703_));
 sg13g2_and3_1 _8353_ (.X(_3707_),
    .A(\welcome_screen_inst.welcome_counter[2] ),
    .B(\welcome_screen_inst.welcome_counter[1] ),
    .C(\welcome_screen_inst.welcome_counter[0] ));
 sg13g2_a21oi_1 _8354_ (.A1(net802),
    .A2(\welcome_screen_inst.welcome_counter[0] ),
    .Y(_3708_),
    .B1(net804));
 sg13g2_nor3_1 _8355_ (.A(_3677_),
    .B(_3707_),
    .C(_3708_),
    .Y(_3709_));
 sg13g2_nor2_1 _8356_ (.A(net2259),
    .B(_3709_),
    .Y(_3710_));
 sg13g2_o21ai_1 _8357_ (.B1(_3710_),
    .Y(_0439_),
    .A1(_3941_),
    .A2(_3701_));
 sg13g2_nand2_1 _8358_ (.Y(_3711_),
    .A(net2285),
    .B(_3700_));
 sg13g2_nand3_1 _8359_ (.B(_3701_),
    .C(_3707_),
    .A(net1005),
    .Y(_3712_));
 sg13g2_a21oi_1 _8360_ (.A1(_3701_),
    .A2(_3707_),
    .Y(_3713_),
    .B1(net1005));
 sg13g2_nor2_1 _8361_ (.A(_3700_),
    .B(_3713_),
    .Y(_3714_));
 sg13g2_a21o_1 _8362_ (.A2(_3714_),
    .A1(net1006),
    .B1(net2259),
    .X(_0440_));
 sg13g2_nor2b_1 _8363_ (.A(net834),
    .B_N(_3712_),
    .Y(_3715_));
 sg13g2_o21ai_1 _8364_ (.B1(net2285),
    .Y(_0441_),
    .A1(_3702_),
    .A2(net835));
 sg13g2_nor2_1 _8365_ (.A(net2103),
    .B(net1775),
    .Y(_3716_));
 sg13g2_nand2b_1 _8366_ (.Y(_3717_),
    .B(net1776),
    .A_N(net2103));
 sg13g2_nor4_1 _8367_ (.A(debug_btn_right),
    .B(debug_btn_up),
    .C(debug_btn_down),
    .D(debug_btn_left),
    .Y(_3718_));
 sg13g2_o21ai_1 _8368_ (.B1(net2266),
    .Y(_3719_),
    .A1(net827),
    .A2(_3716_));
 sg13g2_a21oi_1 _8369_ (.A1(_3716_),
    .A2(_3718_),
    .Y(_0442_),
    .B1(_3719_));
 sg13g2_nor2_1 _8370_ (.A(_0552_),
    .B(_0925_),
    .Y(_3720_));
 sg13g2_or2_1 _8371_ (.X(_3721_),
    .B(_0811_),
    .A(_0580_));
 sg13g2_nand2_1 _8372_ (.Y(_3722_),
    .A(_0562_),
    .B(_0937_));
 sg13g2_nor2_1 _8373_ (.A(_0581_),
    .B(_1007_),
    .Y(_3723_));
 sg13g2_xnor2_1 _8374_ (.Y(_3724_),
    .A(_0549_),
    .B(_0950_));
 sg13g2_and2_1 _8375_ (.A(_0545_),
    .B(_0980_),
    .X(_3725_));
 sg13g2_xnor2_1 _8376_ (.Y(_3726_),
    .A(_0553_),
    .B(_0969_));
 sg13g2_xnor2_1 _8377_ (.Y(_3727_),
    .A(_0560_),
    .B(_0862_));
 sg13g2_and2_1 _8378_ (.A(_0576_),
    .B(_0800_),
    .X(_3728_));
 sg13g2_nor2b_1 _8379_ (.A(_0990_),
    .B_N(_0573_),
    .Y(_3729_));
 sg13g2_and2_1 _8380_ (.A(_0577_),
    .B(_0999_),
    .X(_3730_));
 sg13g2_nor2b_1 _8381_ (.A(_0702_),
    .B_N(_0544_),
    .Y(_3731_));
 sg13g2_and2_1 _8382_ (.A(_0555_),
    .B(_0908_),
    .X(_3732_));
 sg13g2_nor2_1 _8383_ (.A(_0576_),
    .B(_0799_),
    .Y(_3733_));
 sg13g2_nor2b_1 _8384_ (.A(_0575_),
    .B_N(_0783_),
    .Y(_3734_));
 sg13g2_nor2_1 _8385_ (.A(_0579_),
    .B(_0700_),
    .Y(_3735_));
 sg13g2_nor2_1 _8386_ (.A(_0555_),
    .B(_0908_),
    .Y(_3736_));
 sg13g2_nor4_1 _8387_ (.A(_3724_),
    .B(_3731_),
    .C(_3732_),
    .D(_3733_),
    .Y(_3737_));
 sg13g2_xnor2_1 _8388_ (.Y(_3738_),
    .A(_0557_),
    .B(_0960_));
 sg13g2_o21ai_1 _8389_ (.B1(_3722_),
    .Y(_3739_),
    .A1(_0577_),
    .A2(_0998_));
 sg13g2_nor4_1 _8390_ (.A(_3725_),
    .B(_3736_),
    .C(_3738_),
    .D(_3739_),
    .Y(_3740_));
 sg13g2_a221oi_1 _8391_ (.B2(_0580_),
    .C1(_3729_),
    .B1(_0813_),
    .A1(_0574_),
    .Y(_3741_),
    .A2(_0784_));
 sg13g2_a21o_1 _8392_ (.A2(_0925_),
    .A1(_0552_),
    .B1(_3723_),
    .X(_3742_));
 sg13g2_o21ai_1 _8393_ (.B1(_3721_),
    .Y(_3743_),
    .A1(_0562_),
    .A2(_0937_));
 sg13g2_nor4_1 _8394_ (.A(_3726_),
    .B(_3728_),
    .C(_3742_),
    .D(_3743_),
    .Y(_3744_));
 sg13g2_and4_2 _8395_ (.A(_3737_),
    .B(_3740_),
    .C(_3741_),
    .D(_3744_),
    .X(_3745_));
 sg13g2_a21o_1 _8396_ (.A2(_1009_),
    .A1(_0581_),
    .B1(_3727_),
    .X(_3746_));
 sg13g2_xnor2_1 _8397_ (.Y(_3747_),
    .A(_0547_),
    .B(_0890_));
 sg13g2_or4_1 _8398_ (.A(_3720_),
    .B(_3734_),
    .C(_3735_),
    .D(_3747_),
    .X(_3748_));
 sg13g2_nor4_2 _8399_ (.A(\game_logic_inst.valid_move ),
    .B(_3730_),
    .C(_3746_),
    .Y(_3749_),
    .D(_3748_));
 sg13g2_nand3_1 _8400_ (.B(_3745_),
    .C(_3749_),
    .A(net1737),
    .Y(_3750_));
 sg13g2_nor3_2 _8401_ (.A(net2103),
    .B(net1752),
    .C(_0895_),
    .Y(_3751_));
 sg13g2_inv_1 _8402_ (.Y(_3752_),
    .A(_3751_));
 sg13g2_or2_1 _8403_ (.X(_3753_),
    .B(_3751_),
    .A(net1041));
 sg13g2_and4_1 _8404_ (.A(net2266),
    .B(_3717_),
    .C(_3750_),
    .D(_3753_),
    .X(_0443_));
 sg13g2_nand3b_1 _8405_ (.B(net2000),
    .C(net2107),
    .Y(_3754_),
    .A_N(net1752));
 sg13g2_a22oi_1 _8406_ (.Y(_3755_),
    .B1(_3754_),
    .B2(net2119),
    .A2(net1776),
    .A1(net2110));
 sg13g2_nor2_1 _8407_ (.A(net2257),
    .B(_3755_),
    .Y(_0444_));
 sg13g2_and2_1 _8408_ (.A(net2264),
    .B(net424),
    .X(_0445_));
 sg13g2_xor2_1 _8409_ (.B(net993),
    .A(\game_logic_inst.lfsr_shift[0] ),
    .X(_3756_));
 sg13g2_nor2_1 _8410_ (.A(net2257),
    .B(net994),
    .Y(_0446_));
 sg13g2_o21ai_1 _8411_ (.B1(net2103),
    .Y(_3757_),
    .A1(net2256),
    .A2(_3387_));
 sg13g2_o21ai_1 _8412_ (.B1(net2270),
    .Y(_3758_),
    .A1(net1777),
    .A2(_3757_));
 sg13g2_inv_1 _8413_ (.Y(_0447_),
    .A(_3758_));
 sg13g2_nor4_2 _8414_ (.A(net2103),
    .B(_0760_),
    .C(_0761_),
    .Y(_3759_),
    .D(net1917));
 sg13g2_nand2b_1 _8415_ (.Y(_3760_),
    .B(\game_logic_inst.should_transpose ),
    .A_N(net2103));
 sg13g2_nand4_1 _8416_ (.B(net2104),
    .C(_0069_),
    .A(_3940_),
    .Y(_3761_),
    .D(_0760_));
 sg13g2_o21ai_1 _8417_ (.B1(net2055),
    .Y(_3762_),
    .A1(net2256),
    .A2(_3387_));
 sg13g2_nand3_1 _8418_ (.B(_3761_),
    .C(_3762_),
    .A(_3760_),
    .Y(_3763_));
 sg13g2_o21ai_1 _8419_ (.B1(net1775),
    .Y(_3764_),
    .A1(_3759_),
    .A2(_3763_));
 sg13g2_nand3_1 _8420_ (.B(net1998),
    .C(net1737),
    .A(net2104),
    .Y(_3765_));
 sg13g2_nand3_1 _8421_ (.B(_3764_),
    .C(_3765_),
    .A(_3717_),
    .Y(_3766_));
 sg13g2_nand2_1 _8422_ (.Y(_3767_),
    .A(net796),
    .B(_3766_));
 sg13g2_a21oi_1 _8423_ (.A1(_3745_),
    .A2(_3749_),
    .Y(_3768_),
    .B1(\game_logic_inst.debug_move_reg ));
 sg13g2_a21oi_1 _8424_ (.A1(net796),
    .A2(_3940_),
    .Y(_3769_),
    .B1(net2053));
 sg13g2_nor2b_1 _8425_ (.A(_3766_),
    .B_N(_3769_),
    .Y(_3770_));
 sg13g2_o21ai_1 _8426_ (.B1(_3770_),
    .Y(_3771_),
    .A1(_3940_),
    .A2(_3768_));
 sg13g2_a21oi_1 _8427_ (.A1(_3767_),
    .A2(_3771_),
    .Y(_0448_),
    .B1(net2257));
 sg13g2_and2_1 _8428_ (.A(\game_logic_inst.add_new_tiles[1] ),
    .B(\game_logic_inst.add_new_tiles[0] ),
    .X(_3772_));
 sg13g2_o21ai_1 _8429_ (.B1(net440),
    .Y(_3773_),
    .A1(_0760_),
    .A2(_3772_));
 sg13g2_nor2_1 _8430_ (.A(net2103),
    .B(_3766_),
    .Y(_3774_));
 sg13g2_a221oi_1 _8431_ (.B2(_3774_),
    .C1(net2257),
    .B1(net441),
    .A1(_3939_),
    .Y(_0449_),
    .A2(_3766_));
 sg13g2_nand3_1 _8432_ (.B(_0763_),
    .C(_0895_),
    .A(_0524_),
    .Y(_3775_));
 sg13g2_nor2b_2 _8433_ (.A(_3775_),
    .B_N(_0717_),
    .Y(_0450_));
 sg13g2_nor2b_2 _8434_ (.A(_3775_),
    .B_N(_0716_),
    .Y(_0451_));
 sg13g2_nor2_2 _8435_ (.A(_0714_),
    .B(_3775_),
    .Y(_0452_));
 sg13g2_nor2_2 _8436_ (.A(_0708_),
    .B(_3775_),
    .Y(_0453_));
 sg13g2_nand2_1 _8437_ (.Y(_3776_),
    .A(net8),
    .B(net11));
 sg13g2_nand2b_2 _8438_ (.Y(_3777_),
    .B(_3776_),
    .A_N(net12));
 sg13g2_nand2_1 _8439_ (.Y(_3778_),
    .A(net9),
    .B(net8));
 sg13g2_nor3_2 _8440_ (.A(net10),
    .B(_3777_),
    .C(_3778_),
    .Y(_3779_));
 sg13g2_and2_1 _8441_ (.A(net2276),
    .B(net1817),
    .X(_0454_));
 sg13g2_nand3_1 _8442_ (.B(_0513_),
    .C(net1777),
    .A(_0511_),
    .Y(_3780_));
 sg13g2_a21oi_1 _8443_ (.A1(net2107),
    .A2(_3780_),
    .Y(_3781_),
    .B1(net887));
 sg13g2_nor2_1 _8444_ (.A(\game_logic_inst.current_direction[3] ),
    .B(net634),
    .Y(_3782_));
 sg13g2_nor4_1 _8445_ (.A(_3987_),
    .B(net440),
    .C(net1997),
    .D(_3782_),
    .Y(_3783_));
 sg13g2_nor3_1 _8446_ (.A(net2054),
    .B(net1776),
    .C(_3783_),
    .Y(_3784_));
 sg13g2_nor3_1 _8447_ (.A(net2257),
    .B(_3781_),
    .C(_3784_),
    .Y(_0455_));
 sg13g2_nor2_1 _8448_ (.A(net2103),
    .B(net1733),
    .Y(_3785_));
 sg13g2_a22oi_1 _8449_ (.Y(_3786_),
    .B1(_3785_),
    .B2(net673),
    .A2(_3752_),
    .A1(net2099));
 sg13g2_nor2_1 _8450_ (.A(net2257),
    .B(net674),
    .Y(_0456_));
 sg13g2_nand4_1 _8451_ (.B(net2017),
    .C(net1997),
    .A(_0524_),
    .Y(_3787_),
    .D(net1738));
 sg13g2_nand2_1 _8452_ (.Y(_3788_),
    .A(net2096),
    .B(net2269));
 sg13g2_o21ai_1 _8453_ (.B1(_3787_),
    .Y(_0457_),
    .A1(_3751_),
    .A2(_3788_));
 sg13g2_o21ai_1 _8454_ (.B1(net2276),
    .Y(_3789_),
    .A1(net894),
    .A2(net1817));
 sg13g2_mux4_1 _8455_ (.S0(net2081),
    .A0(\debug_controller_inst.grid_in[32] ),
    .A1(\debug_controller_inst.grid_in[36] ),
    .A2(\debug_controller_inst.grid_in[40] ),
    .A3(\debug_controller_inst.grid_in[44] ),
    .S1(net2076),
    .X(_3790_));
 sg13g2_nor2_1 _8456_ (.A(net2072),
    .B(_3790_),
    .Y(_3791_));
 sg13g2_o21ai_1 _8457_ (.B1(net2070),
    .Y(_3792_),
    .A1(net2078),
    .A2(\debug_controller_inst.grid_in[48] ));
 sg13g2_a21oi_1 _8458_ (.A1(net2078),
    .A2(_3980_),
    .Y(_3793_),
    .B1(_3792_));
 sg13g2_nor2_1 _8459_ (.A(net2081),
    .B(\debug_controller_inst.grid_in[56] ),
    .Y(_3794_));
 sg13g2_o21ai_1 _8460_ (.B1(net2075),
    .Y(_3795_),
    .A1(net2069),
    .A2(\debug_controller_inst.grid_in[60] ));
 sg13g2_o21ai_1 _8461_ (.B1(net2071),
    .Y(_3796_),
    .A1(_3794_),
    .A2(_3795_));
 sg13g2_o21ai_1 _8462_ (.B1(\debug_controller_inst.grid_addr[3] ),
    .Y(_3797_),
    .A1(_3793_),
    .A2(_3796_));
 sg13g2_mux4_1 _8463_ (.S0(net2080),
    .A0(\debug_controller_inst.grid_in[0] ),
    .A1(\debug_controller_inst.grid_in[4] ),
    .A2(\debug_controller_inst.grid_in[8] ),
    .A3(\debug_controller_inst.grid_in[12] ),
    .S1(net2075),
    .X(_3798_));
 sg13g2_nor2_1 _8464_ (.A(net2071),
    .B(_3798_),
    .Y(_3799_));
 sg13g2_o21ai_1 _8465_ (.B1(net2070),
    .Y(_3800_),
    .A1(net2078),
    .A2(\debug_controller_inst.grid_in[16] ));
 sg13g2_a21oi_1 _8466_ (.A1(net2078),
    .A2(_3979_),
    .Y(_3801_),
    .B1(_3800_));
 sg13g2_nor2_1 _8467_ (.A(net2069),
    .B(\debug_controller_inst.grid_in[28] ),
    .Y(_3802_));
 sg13g2_o21ai_1 _8468_ (.B1(net2075),
    .Y(_3803_),
    .A1(net2079),
    .A2(\debug_controller_inst.grid_in[24] ));
 sg13g2_o21ai_1 _8469_ (.B1(net2071),
    .Y(_3804_),
    .A1(_3802_),
    .A2(_3803_));
 sg13g2_o21ai_1 _8470_ (.B1(_3929_),
    .Y(_3805_),
    .A1(_3801_),
    .A2(_3804_));
 sg13g2_nor2_1 _8471_ (.A(_3799_),
    .B(_3805_),
    .Y(_3806_));
 sg13g2_o21ai_1 _8472_ (.B1(_3779_),
    .Y(_3807_),
    .A1(_3791_),
    .A2(_3797_));
 sg13g2_nor2_2 _8473_ (.A(_3806_),
    .B(_3807_),
    .Y(_3808_));
 sg13g2_nor2_1 _8474_ (.A(_3789_),
    .B(_3808_),
    .Y(_0458_));
 sg13g2_mux4_1 _8475_ (.S0(net2082),
    .A0(\debug_controller_inst.grid_in[33] ),
    .A1(\debug_controller_inst.grid_in[37] ),
    .A2(\debug_controller_inst.grid_in[41] ),
    .A3(\debug_controller_inst.grid_in[45] ),
    .S1(net2076),
    .X(_3809_));
 sg13g2_nor2_1 _8476_ (.A(net2072),
    .B(_3809_),
    .Y(_3810_));
 sg13g2_o21ai_1 _8477_ (.B1(net2070),
    .Y(_3811_),
    .A1(net2079),
    .A2(\debug_controller_inst.grid_in[49] ));
 sg13g2_a21oi_1 _8478_ (.A1(net2081),
    .A2(_3982_),
    .Y(_3812_),
    .B1(_3811_));
 sg13g2_nor2_1 _8479_ (.A(net2081),
    .B(\debug_controller_inst.grid_in[57] ),
    .Y(_3813_));
 sg13g2_o21ai_1 _8480_ (.B1(net2076),
    .Y(_3814_),
    .A1(net2069),
    .A2(\debug_controller_inst.grid_in[61] ));
 sg13g2_o21ai_1 _8481_ (.B1(net2072),
    .Y(_3815_),
    .A1(_3813_),
    .A2(_3814_));
 sg13g2_o21ai_1 _8482_ (.B1(\debug_controller_inst.grid_addr[3] ),
    .Y(_3816_),
    .A1(_3812_),
    .A2(_3815_));
 sg13g2_mux4_1 _8483_ (.S0(net2080),
    .A0(\debug_controller_inst.grid_in[1] ),
    .A1(\debug_controller_inst.grid_in[5] ),
    .A2(\debug_controller_inst.grid_in[9] ),
    .A3(\debug_controller_inst.grid_in[13] ),
    .S1(net2075),
    .X(_3817_));
 sg13g2_nor2_1 _8484_ (.A(net2071),
    .B(_3817_),
    .Y(_3818_));
 sg13g2_o21ai_1 _8485_ (.B1(net2070),
    .Y(_3819_),
    .A1(net2080),
    .A2(\debug_controller_inst.grid_in[17] ));
 sg13g2_a21oi_1 _8486_ (.A1(net2080),
    .A2(_3981_),
    .Y(_3820_),
    .B1(_3819_));
 sg13g2_nor2_1 _8487_ (.A(net2069),
    .B(\debug_controller_inst.grid_in[29] ),
    .Y(_3821_));
 sg13g2_o21ai_1 _8488_ (.B1(net2075),
    .Y(_3822_),
    .A1(net2081),
    .A2(\debug_controller_inst.grid_in[25] ));
 sg13g2_o21ai_1 _8489_ (.B1(net2071),
    .Y(_3823_),
    .A1(_3821_),
    .A2(_3822_));
 sg13g2_o21ai_1 _8490_ (.B1(_3929_),
    .Y(_3824_),
    .A1(_3820_),
    .A2(_3823_));
 sg13g2_nor2_1 _8491_ (.A(_3818_),
    .B(_3824_),
    .Y(_3825_));
 sg13g2_o21ai_1 _8492_ (.B1(net1817),
    .Y(_3826_),
    .A1(_3810_),
    .A2(_3816_));
 sg13g2_nor2_2 _8493_ (.A(_3825_),
    .B(_3826_),
    .Y(_3827_));
 sg13g2_o21ai_1 _8494_ (.B1(net2275),
    .Y(_3828_),
    .A1(net864),
    .A2(net1817));
 sg13g2_nor2_1 _8495_ (.A(_3827_),
    .B(_3828_),
    .Y(_0459_));
 sg13g2_mux4_1 _8496_ (.S0(net2082),
    .A0(\debug_controller_inst.grid_in[34] ),
    .A1(\debug_controller_inst.grid_in[38] ),
    .A2(\debug_controller_inst.grid_in[42] ),
    .A3(\debug_controller_inst.grid_in[46] ),
    .S1(net2077),
    .X(_3829_));
 sg13g2_nor2_1 _8497_ (.A(net2073),
    .B(_3829_),
    .Y(_3830_));
 sg13g2_o21ai_1 _8498_ (.B1(net2070),
    .Y(_3831_),
    .A1(net2082),
    .A2(\debug_controller_inst.grid_in[50] ));
 sg13g2_a21oi_1 _8499_ (.A1(net2082),
    .A2(_3984_),
    .Y(_3832_),
    .B1(_3831_));
 sg13g2_nor2_1 _8500_ (.A(net2083),
    .B(\debug_controller_inst.grid_in[58] ),
    .Y(_3833_));
 sg13g2_o21ai_1 _8501_ (.B1(net2076),
    .Y(_3834_),
    .A1(_3932_),
    .A2(\debug_controller_inst.grid_in[62] ));
 sg13g2_o21ai_1 _8502_ (.B1(net2073),
    .Y(_3835_),
    .A1(_3833_),
    .A2(_3834_));
 sg13g2_o21ai_1 _8503_ (.B1(\debug_controller_inst.grid_addr[3] ),
    .Y(_3836_),
    .A1(_3832_),
    .A2(_3835_));
 sg13g2_mux4_1 _8504_ (.S0(net2083),
    .A0(\debug_controller_inst.grid_in[2] ),
    .A1(\debug_controller_inst.grid_in[6] ),
    .A2(\debug_controller_inst.grid_in[10] ),
    .A3(\debug_controller_inst.grid_in[14] ),
    .S1(net2077),
    .X(_3837_));
 sg13g2_nor2_1 _8505_ (.A(net2073),
    .B(_3837_),
    .Y(_3838_));
 sg13g2_o21ai_1 _8506_ (.B1(net2070),
    .Y(_3839_),
    .A1(net2082),
    .A2(\debug_controller_inst.grid_in[18] ));
 sg13g2_a21oi_1 _8507_ (.A1(net2082),
    .A2(_3983_),
    .Y(_3840_),
    .B1(_3839_));
 sg13g2_nor2_1 _8508_ (.A(net2069),
    .B(\debug_controller_inst.grid_in[30] ),
    .Y(_3841_));
 sg13g2_o21ai_1 _8509_ (.B1(net2076),
    .Y(_3842_),
    .A1(net2082),
    .A2(\debug_controller_inst.grid_in[26] ));
 sg13g2_o21ai_1 _8510_ (.B1(net2073),
    .Y(_3843_),
    .A1(_3841_),
    .A2(_3842_));
 sg13g2_o21ai_1 _8511_ (.B1(_3929_),
    .Y(_3844_),
    .A1(_3840_),
    .A2(_3843_));
 sg13g2_nor2_1 _8512_ (.A(_3838_),
    .B(_3844_),
    .Y(_3845_));
 sg13g2_o21ai_1 _8513_ (.B1(net1817),
    .Y(_3846_),
    .A1(_3830_),
    .A2(_3836_));
 sg13g2_nor2_2 _8514_ (.A(_3845_),
    .B(_3846_),
    .Y(_3847_));
 sg13g2_o21ai_1 _8515_ (.B1(net2275),
    .Y(_3848_),
    .A1(net865),
    .A2(net1817));
 sg13g2_nor2_1 _8516_ (.A(_3847_),
    .B(_3848_),
    .Y(_0460_));
 sg13g2_o21ai_1 _8517_ (.B1(net2276),
    .Y(_3849_),
    .A1(net897),
    .A2(net1817));
 sg13g2_mux4_1 _8518_ (.S0(net2081),
    .A0(\debug_controller_inst.grid_in[35] ),
    .A1(\debug_controller_inst.grid_in[39] ),
    .A2(\debug_controller_inst.grid_in[43] ),
    .A3(\debug_controller_inst.grid_in[47] ),
    .S1(net2076),
    .X(_3850_));
 sg13g2_nor2_1 _8519_ (.A(net2072),
    .B(_3850_),
    .Y(_3851_));
 sg13g2_o21ai_1 _8520_ (.B1(net2070),
    .Y(_3852_),
    .A1(net2079),
    .A2(\debug_controller_inst.grid_in[51] ));
 sg13g2_a21oi_1 _8521_ (.A1(net2078),
    .A2(_3986_),
    .Y(_3853_),
    .B1(_3852_));
 sg13g2_nor2_1 _8522_ (.A(net2081),
    .B(\debug_controller_inst.grid_in[59] ),
    .Y(_3854_));
 sg13g2_o21ai_1 _8523_ (.B1(net2075),
    .Y(_3855_),
    .A1(net2069),
    .A2(\debug_controller_inst.grid_in[63] ));
 sg13g2_o21ai_1 _8524_ (.B1(net2071),
    .Y(_3856_),
    .A1(_3854_),
    .A2(_3855_));
 sg13g2_o21ai_1 _8525_ (.B1(\debug_controller_inst.grid_addr[3] ),
    .Y(_3857_),
    .A1(_3853_),
    .A2(_3856_));
 sg13g2_mux4_1 _8526_ (.S0(net2078),
    .A0(\debug_controller_inst.grid_in[3] ),
    .A1(\debug_controller_inst.grid_in[7] ),
    .A2(\debug_controller_inst.grid_in[11] ),
    .A3(\debug_controller_inst.grid_in[15] ),
    .S1(net2075),
    .X(_3858_));
 sg13g2_nor2_1 _8527_ (.A(net2071),
    .B(_3858_),
    .Y(_3859_));
 sg13g2_o21ai_1 _8528_ (.B1(net2070),
    .Y(_3860_),
    .A1(net2078),
    .A2(\debug_controller_inst.grid_in[19] ));
 sg13g2_a21oi_1 _8529_ (.A1(net2078),
    .A2(_3985_),
    .Y(_3861_),
    .B1(_3860_));
 sg13g2_nor2_1 _8530_ (.A(net2069),
    .B(\debug_controller_inst.grid_in[31] ),
    .Y(_3862_));
 sg13g2_o21ai_1 _8531_ (.B1(net2075),
    .Y(_3863_),
    .A1(net2079),
    .A2(\debug_controller_inst.grid_in[27] ));
 sg13g2_o21ai_1 _8532_ (.B1(net2071),
    .Y(_3864_),
    .A1(_3862_),
    .A2(_3863_));
 sg13g2_o21ai_1 _8533_ (.B1(_3929_),
    .Y(_3865_),
    .A1(_3861_),
    .A2(_3864_));
 sg13g2_nor2_1 _8534_ (.A(_3859_),
    .B(_3865_),
    .Y(_3866_));
 sg13g2_o21ai_1 _8535_ (.B1(net1817),
    .Y(_3867_),
    .A1(_3851_),
    .A2(_3857_));
 sg13g2_nor2_2 _8536_ (.A(_3866_),
    .B(_3867_),
    .Y(_3868_));
 sg13g2_nor2_1 _8537_ (.A(_3849_),
    .B(_3868_),
    .Y(_0461_));
 sg13g2_nand2_1 _8538_ (.Y(_3869_),
    .A(net8),
    .B(net10));
 sg13g2_nand2_1 _8539_ (.Y(_3870_),
    .A(_3778_),
    .B(_3869_));
 sg13g2_nor4_2 _8540_ (.A(net12),
    .B(net2260),
    .C(_3776_),
    .Y(_3871_),
    .D(_3870_));
 sg13g2_and2_1 _8541_ (.A(net13),
    .B(_3871_),
    .X(_0462_));
 sg13g2_and2_1 _8542_ (.A(net14),
    .B(_3871_),
    .X(_0463_));
 sg13g2_and2_1 _8543_ (.A(net15),
    .B(_3871_),
    .X(_0464_));
 sg13g2_and2_1 _8544_ (.A(net16),
    .B(_3871_),
    .X(_0465_));
 sg13g2_nor3_2 _8545_ (.A(net9),
    .B(_3777_),
    .C(_3869_),
    .Y(_3872_));
 sg13g2_and2_1 _8546_ (.A(net2276),
    .B(net1815),
    .X(_0466_));
 sg13g2_o21ai_1 _8547_ (.B1(net2275),
    .Y(_3873_),
    .A1(net2093),
    .A2(_3872_));
 sg13g2_a21oi_1 _8548_ (.A1(_3937_),
    .A2(_3872_),
    .Y(_0467_),
    .B1(_3873_));
 sg13g2_o21ai_1 _8549_ (.B1(net2277),
    .Y(_3874_),
    .A1(net2091),
    .A2(net1816));
 sg13g2_a21oi_1 _8550_ (.A1(_3935_),
    .A2(net1816),
    .Y(_0468_),
    .B1(_3874_));
 sg13g2_o21ai_1 _8551_ (.B1(net2277),
    .Y(_3875_),
    .A1(net2089),
    .A2(net1816));
 sg13g2_a21oi_1 _8552_ (.A1(_3934_),
    .A2(net1816),
    .Y(_0469_),
    .B1(_3875_));
 sg13g2_o21ai_1 _8553_ (.B1(net2275),
    .Y(_3876_),
    .A1(net2087),
    .A2(net1816));
 sg13g2_a21oi_1 _8554_ (.A1(_3933_),
    .A2(net1816),
    .Y(_0470_),
    .B1(_3876_));
 sg13g2_o21ai_1 _8555_ (.B1(net2278),
    .Y(_3877_),
    .A1(\debug_controller_inst.grid_out_addr[0] ),
    .A2(net1816));
 sg13g2_a21oi_1 _8556_ (.A1(net2069),
    .A2(net1815),
    .Y(_0471_),
    .B1(_3877_));
 sg13g2_o21ai_1 _8557_ (.B1(net2278),
    .Y(_3878_),
    .A1(\debug_controller_inst.grid_out_addr[1] ),
    .A2(net1815));
 sg13g2_a21oi_1 _8558_ (.A1(_3931_),
    .A2(net1815),
    .Y(_0472_),
    .B1(_3878_));
 sg13g2_o21ai_1 _8559_ (.B1(net2277),
    .Y(_3879_),
    .A1(net2085),
    .A2(net1815));
 sg13g2_a21oi_1 _8560_ (.A1(_3930_),
    .A2(net1815),
    .Y(_0473_),
    .B1(_3879_));
 sg13g2_o21ai_1 _8561_ (.B1(net2278),
    .Y(_3880_),
    .A1(net895),
    .A2(net1815));
 sg13g2_a21oi_1 _8562_ (.A1(_3929_),
    .A2(net1815),
    .Y(_0474_),
    .B1(_3880_));
 sg13g2_and2_1 _8563_ (.A(net2287),
    .B(net890),
    .X(_0475_));
 sg13g2_nand3_1 _8564_ (.B(net8),
    .C(net10),
    .A(net9),
    .Y(_3881_));
 sg13g2_inv_1 _8565_ (.Y(_3882_),
    .A(_3881_));
 sg13g2_nand2b_2 _8566_ (.Y(_3883_),
    .B(_3882_),
    .A_N(_3777_));
 sg13g2_nor2b_2 _8567_ (.A(_3777_),
    .B_N(_3870_),
    .Y(_3884_));
 sg13g2_nand2b_1 _8568_ (.Y(_3885_),
    .B(_3870_),
    .A_N(_3777_));
 sg13g2_a22oi_1 _8569_ (.Y(_3886_),
    .B1(_3883_),
    .B2(net438),
    .A2(_3882_),
    .A1(net13));
 sg13g2_o21ai_1 _8570_ (.B1(net2277),
    .Y(_3887_),
    .A1(net2083),
    .A2(_3884_));
 sg13g2_a21oi_1 _8571_ (.A1(_3884_),
    .A2(_3886_),
    .Y(_0476_),
    .B1(_3887_));
 sg13g2_nand2_1 _8572_ (.Y(_3888_),
    .A(net2077),
    .B(net2083));
 sg13g2_a21o_1 _8573_ (.A2(_3888_),
    .A1(_3881_),
    .B1(_3885_),
    .X(_3889_));
 sg13g2_nor2_1 _8574_ (.A(_3935_),
    .B(_3883_),
    .Y(_3890_));
 sg13g2_o21ai_1 _8575_ (.B1(_3884_),
    .Y(_3891_),
    .A1(net2083),
    .A2(_3882_));
 sg13g2_o21ai_1 _8576_ (.B1(net2277),
    .Y(_3892_),
    .A1(_3889_),
    .A2(_3890_));
 sg13g2_a21oi_1 _8577_ (.A1(_3931_),
    .A2(_3891_),
    .Y(_0477_),
    .B1(_3892_));
 sg13g2_o21ai_1 _8578_ (.B1(_3883_),
    .Y(_3893_),
    .A1(net2074),
    .A2(_3888_));
 sg13g2_o21ai_1 _8579_ (.B1(_3884_),
    .Y(_3894_),
    .A1(net15),
    .A2(_3881_));
 sg13g2_inv_1 _8580_ (.Y(_3895_),
    .A(_3894_));
 sg13g2_a22oi_1 _8581_ (.Y(_3896_),
    .B1(_3893_),
    .B2(_3895_),
    .A2(_3889_),
    .A1(net2074));
 sg13g2_nor2_1 _8582_ (.A(net2260),
    .B(_3896_),
    .Y(_0478_));
 sg13g2_nor2_1 _8583_ (.A(net1011),
    .B(_3888_),
    .Y(_3897_));
 sg13g2_xnor2_1 _8584_ (.Y(_3898_),
    .A(\debug_controller_inst.grid_addr[3] ),
    .B(_3897_));
 sg13g2_a221oi_1 _8585_ (.B2(_3898_),
    .C1(_3885_),
    .B1(_3883_),
    .A1(_3933_),
    .Y(_3899_),
    .A2(_3882_));
 sg13g2_a21oi_1 _8586_ (.A1(\debug_controller_inst.grid_addr[3] ),
    .A2(_3885_),
    .Y(_3900_),
    .B1(_3899_));
 sg13g2_nor2_1 _8587_ (.A(net2260),
    .B(net1012),
    .Y(_0479_));
 sg13g2_nor3_2 _8588_ (.A(\lfsr_inst.lfsr[30] ),
    .B(\lfsr_inst.lfsr[31] ),
    .C(_3684_),
    .Y(_3901_));
 sg13g2_o21ai_1 _8589_ (.B1(\lfsr_inst.lfsr[31] ),
    .Y(_3902_),
    .A1(\lfsr_inst.lfsr[30] ),
    .A2(_3684_));
 sg13g2_nor2b_2 _8590_ (.A(_3901_),
    .B_N(_3902_),
    .Y(_3903_));
 sg13g2_nand2b_2 _8591_ (.Y(_3904_),
    .B(_3902_),
    .A_N(_3901_));
 sg13g2_nor4_1 _8592_ (.A(net2251),
    .B(_3679_),
    .C(net1780),
    .D(_3903_),
    .Y(_3905_));
 sg13g2_a21o_1 _8593_ (.A2(net1780),
    .A1(net851),
    .B1(_3905_),
    .X(_0480_));
 sg13g2_nor4_1 _8594_ (.A(net2251),
    .B(_3681_),
    .C(net1780),
    .D(_3903_),
    .Y(_3906_));
 sg13g2_a21o_1 _8595_ (.A2(net1780),
    .A1(net819),
    .B1(_3906_),
    .X(_0481_));
 sg13g2_nor4_1 _8596_ (.A(net2251),
    .B(_3686_),
    .C(net1780),
    .D(_3903_),
    .Y(_3907_));
 sg13g2_a21o_1 _8597_ (.A2(net1780),
    .A1(net858),
    .B1(_3907_),
    .X(_0482_));
 sg13g2_nand3_1 _8598_ (.B(_3685_),
    .C(_3904_),
    .A(net2250),
    .Y(_3908_));
 sg13g2_nand2_1 _8599_ (.Y(_3909_),
    .A(net723),
    .B(net1779));
 sg13g2_o21ai_1 _8600_ (.B1(_3909_),
    .Y(_0483_),
    .A1(net1779),
    .A2(_3908_));
 sg13g2_nand3_1 _8601_ (.B(_3680_),
    .C(_3904_),
    .A(net2250),
    .Y(_3910_));
 sg13g2_nand2_1 _8602_ (.Y(_3911_),
    .A(net716),
    .B(net1778));
 sg13g2_o21ai_1 _8603_ (.B1(_3911_),
    .Y(_0484_),
    .A1(net1778),
    .A2(_3910_));
 sg13g2_nand3_1 _8604_ (.B(_3680_),
    .C(_3903_),
    .A(net2250),
    .Y(_3912_));
 sg13g2_nand2_1 _8605_ (.Y(_3913_),
    .A(net695),
    .B(net1778));
 sg13g2_o21ai_1 _8606_ (.B1(_3913_),
    .Y(_0485_),
    .A1(net1778),
    .A2(_3912_));
 sg13g2_nand3_1 _8607_ (.B(_3683_),
    .C(_3903_),
    .A(net2250),
    .Y(_3914_));
 sg13g2_nand2_1 _8608_ (.Y(_3915_),
    .A(net664),
    .B(net1779));
 sg13g2_o21ai_1 _8609_ (.B1(_3915_),
    .Y(_0486_),
    .A1(net1779),
    .A2(_3914_));
 sg13g2_nand2_1 _8610_ (.Y(_3916_),
    .A(net2250),
    .B(_3901_));
 sg13g2_nand2_1 _8611_ (.Y(_3917_),
    .A(net755),
    .B(net1778));
 sg13g2_o21ai_1 _8612_ (.B1(_3917_),
    .Y(_0487_),
    .A1(net1778),
    .A2(_3916_));
 sg13g2_nor4_1 _8613_ (.A(net2251),
    .B(_3679_),
    .C(net1781),
    .D(_3904_),
    .Y(_3918_));
 sg13g2_a21o_1 _8614_ (.A2(net1780),
    .A1(net841),
    .B1(_3918_),
    .X(_0488_));
 sg13g2_nand3_1 _8615_ (.B(_3678_),
    .C(_3904_),
    .A(net2250),
    .Y(_3919_));
 sg13g2_nand2_1 _8616_ (.Y(_3920_),
    .A(net794),
    .B(net1779));
 sg13g2_o21ai_1 _8617_ (.B1(_3920_),
    .Y(_0489_),
    .A1(_3711_),
    .A2(_3919_));
 sg13g2_nor4_1 _8618_ (.A(net2251),
    .B(_3684_),
    .C(net1782),
    .D(_3904_),
    .Y(_3921_));
 sg13g2_a21o_1 _8619_ (.A2(net1781),
    .A1(net860),
    .B1(_3921_),
    .X(_0490_));
 sg13g2_nor4_1 _8620_ (.A(net2251),
    .B(_3684_),
    .C(net1782),
    .D(_3902_),
    .Y(_3922_));
 sg13g2_a21o_1 _8621_ (.A2(net1782),
    .A1(net884),
    .B1(_3922_),
    .X(_0491_));
 sg13g2_nor4_1 _8622_ (.A(net2251),
    .B(_3686_),
    .C(net1781),
    .D(_3904_),
    .Y(_3923_));
 sg13g2_a21o_1 _8623_ (.A2(net1781),
    .A1(net856),
    .B1(_3923_),
    .X(_0492_));
 sg13g2_nor4_1 _8624_ (.A(net2251),
    .B(_3681_),
    .C(net1780),
    .D(_3904_),
    .Y(_3924_));
 sg13g2_a21o_1 _8625_ (.A2(net1781),
    .A1(net879),
    .B1(_3924_),
    .X(_0493_));
 sg13g2_nand3_1 _8626_ (.B(_3685_),
    .C(_3903_),
    .A(net2250),
    .Y(_3925_));
 sg13g2_nand2_1 _8627_ (.Y(_3926_),
    .A(net813),
    .B(net1778));
 sg13g2_o21ai_1 _8628_ (.B1(_3926_),
    .Y(_0494_),
    .A1(net1779),
    .A2(_3925_));
 sg13g2_nand3_1 _8629_ (.B(_3678_),
    .C(_3903_),
    .A(net2250),
    .Y(_3927_));
 sg13g2_nand2_1 _8630_ (.Y(_3928_),
    .A(net778),
    .B(net1779));
 sg13g2_o21ai_1 _8631_ (.B1(_3928_),
    .Y(_0495_),
    .A1(net1778),
    .A2(_3927_));
 sg13g2_dfrbp_1 _8632_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net204),
    .D(_0176_),
    .Q_N(_4307_),
    .Q(vsync_prev));
 sg13g2_dfrbp_1 _8633_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net201),
    .D(_0177_),
    .Q_N(_4306_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _8634_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net200),
    .D(_0178_),
    .Q_N(_4305_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _8635_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net199),
    .D(net1038),
    .Q_N(_4304_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _8636_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net198),
    .D(_0180_),
    .Q_N(_4303_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _8637_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net197),
    .D(_0181_),
    .Q_N(_4302_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _8638_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net196),
    .D(_0182_),
    .Q_N(_4301_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _8639_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net195),
    .D(net522),
    .Q_N(_4300_),
    .Q(\draw_game_inst.grid[0] ));
 sg13g2_dfrbp_1 _8640_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net193),
    .D(net514),
    .Q_N(_4299_),
    .Q(\draw_game_inst.grid[1] ));
 sg13g2_dfrbp_1 _8641_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net191),
    .D(_0185_),
    .Q_N(_4298_),
    .Q(\draw_game_inst.grid[2] ));
 sg13g2_dfrbp_1 _8642_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net189),
    .D(net598),
    .Q_N(_4297_),
    .Q(\draw_game_inst.grid[3] ));
 sg13g2_dfrbp_1 _8643_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net187),
    .D(net682),
    .Q_N(_4296_),
    .Q(\draw_game_inst.grid[4] ));
 sg13g2_dfrbp_1 _8644_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net185),
    .D(net698),
    .Q_N(_4295_),
    .Q(\draw_game_inst.grid[5] ));
 sg13g2_dfrbp_1 _8645_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net183),
    .D(_0189_),
    .Q_N(_4294_),
    .Q(\draw_game_inst.grid[6] ));
 sg13g2_dfrbp_1 _8646_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net181),
    .D(net692),
    .Q_N(_4293_),
    .Q(\draw_game_inst.grid[7] ));
 sg13g2_dfrbp_1 _8647_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net179),
    .D(net633),
    .Q_N(_4292_),
    .Q(\draw_game_inst.grid[8] ));
 sg13g2_dfrbp_1 _8648_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net177),
    .D(net587),
    .Q_N(_4291_),
    .Q(\draw_game_inst.grid[9] ));
 sg13g2_dfrbp_1 _8649_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net175),
    .D(_0193_),
    .Q_N(_4290_),
    .Q(\draw_game_inst.grid[10] ));
 sg13g2_dfrbp_1 _8650_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net173),
    .D(net676),
    .Q_N(_4289_),
    .Q(\draw_game_inst.grid[11] ));
 sg13g2_dfrbp_1 _8651_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net171),
    .D(net561),
    .Q_N(_4288_),
    .Q(\draw_game_inst.grid[12] ));
 sg13g2_dfrbp_1 _8652_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net169),
    .D(net578),
    .Q_N(_4287_),
    .Q(\draw_game_inst.grid[13] ));
 sg13g2_dfrbp_1 _8653_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net167),
    .D(_0197_),
    .Q_N(_4286_),
    .Q(\draw_game_inst.grid[14] ));
 sg13g2_dfrbp_1 _8654_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net165),
    .D(net450),
    .Q_N(_4285_),
    .Q(\draw_game_inst.grid[15] ));
 sg13g2_dfrbp_1 _8655_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net163),
    .D(net553),
    .Q_N(_4284_),
    .Q(\draw_game_inst.grid[16] ));
 sg13g2_dfrbp_1 _8656_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net161),
    .D(net661),
    .Q_N(_4283_),
    .Q(\draw_game_inst.grid[17] ));
 sg13g2_dfrbp_1 _8657_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net159),
    .D(_0201_),
    .Q_N(_4282_),
    .Q(\draw_game_inst.grid[18] ));
 sg13g2_dfrbp_1 _8658_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net157),
    .D(net605),
    .Q_N(_4281_),
    .Q(\draw_game_inst.grid[19] ));
 sg13g2_dfrbp_1 _8659_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net155),
    .D(net616),
    .Q_N(_4280_),
    .Q(\draw_game_inst.grid[20] ));
 sg13g2_dfrbp_1 _8660_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net153),
    .D(net565),
    .Q_N(_4279_),
    .Q(\draw_game_inst.grid[21] ));
 sg13g2_dfrbp_1 _8661_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net151),
    .D(_0205_),
    .Q_N(_4278_),
    .Q(\draw_game_inst.grid[22] ));
 sg13g2_dfrbp_1 _8662_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net149),
    .D(net647),
    .Q_N(_4277_),
    .Q(\draw_game_inst.grid[23] ));
 sg13g2_dfrbp_1 _8663_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net147),
    .D(net622),
    .Q_N(_4276_),
    .Q(\draw_game_inst.grid[24] ));
 sg13g2_dfrbp_1 _8664_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net145),
    .D(net592),
    .Q_N(_4275_),
    .Q(\draw_game_inst.grid[25] ));
 sg13g2_dfrbp_1 _8665_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net143),
    .D(_0209_),
    .Q_N(_4274_),
    .Q(\draw_game_inst.grid[26] ));
 sg13g2_dfrbp_1 _8666_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net141),
    .D(net639),
    .Q_N(_4273_),
    .Q(\draw_game_inst.grid[27] ));
 sg13g2_dfrbp_1 _8667_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net139),
    .D(net600),
    .Q_N(_4272_),
    .Q(\draw_game_inst.grid[28] ));
 sg13g2_dfrbp_1 _8668_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net137),
    .D(net618),
    .Q_N(_4271_),
    .Q(\draw_game_inst.grid[29] ));
 sg13g2_dfrbp_1 _8669_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net135),
    .D(_0213_),
    .Q_N(_4270_),
    .Q(\draw_game_inst.grid[30] ));
 sg13g2_dfrbp_1 _8670_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net133),
    .D(net614),
    .Q_N(_4269_),
    .Q(\draw_game_inst.grid[31] ));
 sg13g2_dfrbp_1 _8671_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net131),
    .D(net542),
    .Q_N(_4268_),
    .Q(\draw_game_inst.grid[32] ));
 sg13g2_dfrbp_1 _8672_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net129),
    .D(net491),
    .Q_N(_4267_),
    .Q(\draw_game_inst.grid[33] ));
 sg13g2_dfrbp_1 _8673_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net127),
    .D(_0217_),
    .Q_N(_4266_),
    .Q(\draw_game_inst.grid[34] ));
 sg13g2_dfrbp_1 _8674_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net125),
    .D(net485),
    .Q_N(_4265_),
    .Q(\draw_game_inst.grid[35] ));
 sg13g2_dfrbp_1 _8675_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net123),
    .D(net563),
    .Q_N(_4264_),
    .Q(\draw_game_inst.grid[36] ));
 sg13g2_dfrbp_1 _8676_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net121),
    .D(net520),
    .Q_N(_4263_),
    .Q(\draw_game_inst.grid[37] ));
 sg13g2_dfrbp_1 _8677_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net119),
    .D(_0221_),
    .Q_N(_4262_),
    .Q(\draw_game_inst.grid[38] ));
 sg13g2_dfrbp_1 _8678_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net117),
    .D(net524),
    .Q_N(_4261_),
    .Q(\draw_game_inst.grid[39] ));
 sg13g2_dfrbp_1 _8679_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net115),
    .D(net669),
    .Q_N(_4260_),
    .Q(\draw_game_inst.grid[40] ));
 sg13g2_dfrbp_1 _8680_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net113),
    .D(net516),
    .Q_N(_4259_),
    .Q(\draw_game_inst.grid[41] ));
 sg13g2_dfrbp_1 _8681_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net111),
    .D(_0225_),
    .Q_N(_4258_),
    .Q(\draw_game_inst.grid[42] ));
 sg13g2_dfrbp_1 _8682_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net109),
    .D(net538),
    .Q_N(_4257_),
    .Q(\draw_game_inst.grid[43] ));
 sg13g2_dfrbp_1 _8683_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net107),
    .D(net620),
    .Q_N(_4256_),
    .Q(\draw_game_inst.grid[44] ));
 sg13g2_dfrbp_1 _8684_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net105),
    .D(net464),
    .Q_N(_4255_),
    .Q(\draw_game_inst.grid[45] ));
 sg13g2_dfrbp_1 _8685_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net103),
    .D(_0229_),
    .Q_N(_4254_),
    .Q(\draw_game_inst.grid[46] ));
 sg13g2_dfrbp_1 _8686_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net101),
    .D(net530),
    .Q_N(_4253_),
    .Q(\draw_game_inst.grid[47] ));
 sg13g2_dfrbp_1 _8687_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net99),
    .D(net694),
    .Q_N(_4252_),
    .Q(\draw_game_inst.grid[48] ));
 sg13g2_dfrbp_1 _8688_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net97),
    .D(net680),
    .Q_N(_4251_),
    .Q(\draw_game_inst.grid[49] ));
 sg13g2_dfrbp_1 _8689_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net95),
    .D(_0233_),
    .Q_N(_4250_),
    .Q(\draw_game_inst.grid[50] ));
 sg13g2_dfrbp_1 _8690_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net93),
    .D(net574),
    .Q_N(_4249_),
    .Q(\draw_game_inst.grid[51] ));
 sg13g2_dfrbp_1 _8691_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net91),
    .D(net546),
    .Q_N(_4248_),
    .Q(\draw_game_inst.grid[52] ));
 sg13g2_dfrbp_1 _8692_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net89),
    .D(net559),
    .Q_N(_4247_),
    .Q(\draw_game_inst.grid[53] ));
 sg13g2_dfrbp_1 _8693_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net87),
    .D(_0237_),
    .Q_N(_4246_),
    .Q(\draw_game_inst.grid[54] ));
 sg13g2_dfrbp_1 _8694_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net85),
    .D(net534),
    .Q_N(_4245_),
    .Q(\draw_game_inst.grid[55] ));
 sg13g2_dfrbp_1 _8695_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net83),
    .D(net637),
    .Q_N(_4244_),
    .Q(\draw_game_inst.grid[56] ));
 sg13g2_dfrbp_1 _8696_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net81),
    .D(net645),
    .Q_N(_4243_),
    .Q(\draw_game_inst.grid[57] ));
 sg13g2_dfrbp_1 _8697_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net79),
    .D(_0241_),
    .Q_N(_4242_),
    .Q(\draw_game_inst.grid[58] ));
 sg13g2_dfrbp_1 _8698_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net77),
    .D(net540),
    .Q_N(_4241_),
    .Q(\draw_game_inst.grid[59] ));
 sg13g2_dfrbp_1 _8699_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net75),
    .D(net707),
    .Q_N(_4240_),
    .Q(\draw_game_inst.grid[60] ));
 sg13g2_dfrbp_1 _8700_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net73),
    .D(net557),
    .Q_N(_4239_),
    .Q(\draw_game_inst.grid[61] ));
 sg13g2_dfrbp_1 _8701_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net71),
    .D(_0245_),
    .Q_N(_4238_),
    .Q(\draw_game_inst.grid[62] ));
 sg13g2_dfrbp_1 _8702_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net69),
    .D(net549),
    .Q_N(_4237_),
    .Q(\draw_game_inst.grid[63] ));
 sg13g2_dfrbp_1 _8703_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net67),
    .D(_0247_),
    .Q_N(_0165_),
    .Q(show_welcome_screen));
 sg13g2_dfrbp_1 _8704_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net65),
    .D(_0248_),
    .Q_N(_4236_),
    .Q(btn_select_prev));
 sg13g2_dfrbp_1 _8705_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net64),
    .D(_0249_),
    .Q_N(_4235_),
    .Q(\draw_game_inst.new_tiles[0] ));
 sg13g2_dfrbp_1 _8706_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net63),
    .D(net474),
    .Q_N(_0070_),
    .Q(\draw_game_inst.new_tiles[1] ));
 sg13g2_dfrbp_1 _8707_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net62),
    .D(net607),
    .Q_N(_0071_),
    .Q(\draw_game_inst.new_tiles[2] ));
 sg13g2_dfrbp_1 _8708_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net61),
    .D(net612),
    .Q_N(_0072_),
    .Q(\draw_game_inst.new_tiles[3] ));
 sg13g2_dfrbp_1 _8709_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net60),
    .D(net641),
    .Q_N(_0073_),
    .Q(\draw_game_inst.new_tiles[4] ));
 sg13g2_dfrbp_1 _8710_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net59),
    .D(net793),
    .Q_N(_0074_),
    .Q(\draw_game_inst.new_tiles[5] ));
 sg13g2_dfrbp_1 _8711_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net58),
    .D(net719),
    .Q_N(_0075_),
    .Q(\draw_game_inst.new_tiles[6] ));
 sg13g2_dfrbp_1 _8712_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net57),
    .D(net500),
    .Q_N(_0076_),
    .Q(\draw_game_inst.new_tiles[7] ));
 sg13g2_dfrbp_1 _8713_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net56),
    .D(net667),
    .Q_N(_0077_),
    .Q(\draw_game_inst.new_tiles[8] ));
 sg13g2_dfrbp_1 _8714_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net55),
    .D(net643),
    .Q_N(_0078_),
    .Q(\draw_game_inst.new_tiles[9] ));
 sg13g2_dfrbp_1 _8715_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net54),
    .D(net526),
    .Q_N(_0079_),
    .Q(\draw_game_inst.new_tiles[10] ));
 sg13g2_dfrbp_1 _8716_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net53),
    .D(net576),
    .Q_N(_0080_),
    .Q(\draw_game_inst.new_tiles[11] ));
 sg13g2_dfrbp_1 _8717_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net52),
    .D(net657),
    .Q_N(_0081_),
    .Q(\draw_game_inst.new_tiles[12] ));
 sg13g2_dfrbp_1 _8718_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net51),
    .D(net572),
    .Q_N(_0082_),
    .Q(\draw_game_inst.new_tiles[13] ));
 sg13g2_dfrbp_1 _8719_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net50),
    .D(net746),
    .Q_N(_0083_),
    .Q(\draw_game_inst.new_tiles[14] ));
 sg13g2_dfrbp_1 _8720_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net49),
    .D(net651),
    .Q_N(_0084_),
    .Q(\draw_game_inst.new_tiles[15] ));
 sg13g2_dfrbp_1 _8721_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net48),
    .D(net447),
    .Q_N(_0085_),
    .Q(\new_tiles_counter[0] ));
 sg13g2_dfrbp_1 _8722_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net47),
    .D(_0266_),
    .Q_N(_0086_),
    .Q(\draw_game_inst.new_tiles_counter[0] ));
 sg13g2_dfrbp_1 _8723_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net46),
    .D(net838),
    .Q_N(_4234_),
    .Q(\draw_game_inst.new_tiles_counter[1] ));
 sg13g2_dfrbp_1 _8724_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net45),
    .D(net845),
    .Q_N(_0087_),
    .Q(\draw_game_inst.new_tiles_counter[2] ));
 sg13g2_dfrbp_1 _8725_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net44),
    .D(_0269_),
    .Q_N(_4233_),
    .Q(\new_tiles_counter[4] ));
 sg13g2_dfrbp_1 _8726_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net43),
    .D(net433),
    .Q_N(_0168_),
    .Q(retro_colors));
 sg13g2_dfrbp_1 _8727_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net41),
    .D(_0271_),
    .Q_N(_4232_),
    .Q(\btn_up_debounce.button_sync_0 ));
 sg13g2_dfrbp_1 _8728_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net40),
    .D(_0272_),
    .Q_N(_0175_),
    .Q(\btn_up_debounce.debounce_counter[0] ));
 sg13g2_dfrbp_1 _8729_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net39),
    .D(_0273_),
    .Q_N(_4231_),
    .Q(\btn_up_debounce.debounce_counter[1] ));
 sg13g2_dfrbp_1 _8730_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net38),
    .D(net503),
    .Q_N(_4230_),
    .Q(\btn_up_debounce.debounce_counter[2] ));
 sg13g2_dfrbp_1 _8731_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net37),
    .D(_0275_),
    .Q_N(_4229_),
    .Q(\btn_up_debounce.debounce_counter[3] ));
 sg13g2_dfrbp_1 _8732_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net36),
    .D(_0276_),
    .Q_N(_4228_),
    .Q(\btn_up_debounce.debounce_counter[4] ));
 sg13g2_dfrbp_1 _8733_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net35),
    .D(net713),
    .Q_N(_4227_),
    .Q(\btn_up_debounce.debounce_counter[5] ));
 sg13g2_dfrbp_1 _8734_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net34),
    .D(_0278_),
    .Q_N(_4226_),
    .Q(\btn_up_debounce.debounce_counter[6] ));
 sg13g2_dfrbp_1 _8735_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net33),
    .D(_0279_),
    .Q_N(_4225_),
    .Q(\btn_up_debounce.debounce_counter[7] ));
 sg13g2_dfrbp_1 _8736_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net32),
    .D(_0280_),
    .Q_N(_4224_),
    .Q(\btn_up_debounce.debounce_counter[8] ));
 sg13g2_dfrbp_1 _8737_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net31),
    .D(_0281_),
    .Q_N(_4223_),
    .Q(\btn_up_debounce.debounce_counter[9] ));
 sg13g2_dfrbp_1 _8738_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net30),
    .D(net595),
    .Q_N(_4222_),
    .Q(\btn_up_debounce.debounce_counter[10] ));
 sg13g2_dfrbp_1 _8739_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net29),
    .D(_0283_),
    .Q_N(_4221_),
    .Q(\btn_up_debounce.debounce_counter[11] ));
 sg13g2_dfrbp_1 _8740_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net28),
    .D(net654),
    .Q_N(_4220_),
    .Q(\btn_up_debounce.debounce_counter[12] ));
 sg13g2_dfrbp_1 _8741_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net27),
    .D(_0285_),
    .Q_N(_4219_),
    .Q(\btn_up_debounce.debounce_counter[13] ));
 sg13g2_dfrbp_1 _8742_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net26),
    .D(_0286_),
    .Q_N(_4218_),
    .Q(\btn_up_debounce.debounce_counter[14] ));
 sg13g2_dfrbp_1 _8743_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net25),
    .D(_0287_),
    .Q_N(_4217_),
    .Q(\btn_up_debounce.debounce_counter[15] ));
 sg13g2_dfrbp_1 _8744_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net415),
    .D(_0288_),
    .Q_N(_4216_),
    .Q(\btn_up_debounce.debounce_counter[16] ));
 sg13g2_dfrbp_1 _8745_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net414),
    .D(net722),
    .Q_N(_4215_),
    .Q(\btn_up_debounce.debounce_counter[17] ));
 sg13g2_dfrbp_1 _8746_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net413),
    .D(_0290_),
    .Q_N(_4214_),
    .Q(\btn_right_debounce.button_sync_1 ));
 sg13g2_dfrbp_1 _8747_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net412),
    .D(net877),
    .Q_N(_4213_),
    .Q(\btn_up_debounce.debounced ));
 sg13g2_dfrbp_1 _8748_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net410),
    .D(_0292_),
    .Q_N(_4212_),
    .Q(\btn_down_debounce.button_sync_0 ));
 sg13g2_dfrbp_1 _8749_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net409),
    .D(_0293_),
    .Q_N(_0174_),
    .Q(\btn_down_debounce.debounce_counter[0] ));
 sg13g2_dfrbp_1 _8750_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net408),
    .D(net873),
    .Q_N(_4211_),
    .Q(\btn_down_debounce.debounce_counter[1] ));
 sg13g2_dfrbp_1 _8751_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net407),
    .D(net730),
    .Q_N(_4210_),
    .Q(\btn_down_debounce.debounce_counter[2] ));
 sg13g2_dfrbp_1 _8752_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net406),
    .D(net710),
    .Q_N(_4209_),
    .Q(\btn_down_debounce.debounce_counter[3] ));
 sg13g2_dfrbp_1 _8753_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net405),
    .D(_0297_),
    .Q_N(_4208_),
    .Q(\btn_down_debounce.debounce_counter[4] ));
 sg13g2_dfrbp_1 _8754_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net404),
    .D(net702),
    .Q_N(_4207_),
    .Q(\btn_down_debounce.debounce_counter[5] ));
 sg13g2_dfrbp_1 _8755_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net403),
    .D(_0299_),
    .Q_N(_4206_),
    .Q(\btn_down_debounce.debounce_counter[6] ));
 sg13g2_dfrbp_1 _8756_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net402),
    .D(_0300_),
    .Q_N(_4205_),
    .Q(\btn_down_debounce.debounce_counter[7] ));
 sg13g2_dfrbp_1 _8757_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net401),
    .D(_0301_),
    .Q_N(_4204_),
    .Q(\btn_down_debounce.debounce_counter[8] ));
 sg13g2_dfrbp_1 _8758_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net400),
    .D(_0302_),
    .Q_N(_4203_),
    .Q(\btn_down_debounce.debounce_counter[9] ));
 sg13g2_dfrbp_1 _8759_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net399),
    .D(net603),
    .Q_N(_4202_),
    .Q(\btn_down_debounce.debounce_counter[10] ));
 sg13g2_dfrbp_1 _8760_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net398),
    .D(_0304_),
    .Q_N(_4201_),
    .Q(\btn_down_debounce.debounce_counter[11] ));
 sg13g2_dfrbp_1 _8761_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net397),
    .D(net610),
    .Q_N(_4200_),
    .Q(\btn_down_debounce.debounce_counter[12] ));
 sg13g2_dfrbp_1 _8762_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net396),
    .D(_0306_),
    .Q_N(_4199_),
    .Q(\btn_down_debounce.debounce_counter[13] ));
 sg13g2_dfrbp_1 _8763_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net395),
    .D(_0307_),
    .Q_N(_4198_),
    .Q(\btn_down_debounce.debounce_counter[14] ));
 sg13g2_dfrbp_1 _8764_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net394),
    .D(_0308_),
    .Q_N(_4197_),
    .Q(\btn_down_debounce.debounce_counter[15] ));
 sg13g2_dfrbp_1 _8765_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net393),
    .D(net585),
    .Q_N(_4196_),
    .Q(\btn_down_debounce.debounce_counter[16] ));
 sg13g2_dfrbp_1 _8766_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net392),
    .D(net494),
    .Q_N(_4195_),
    .Q(\btn_down_debounce.debounce_counter[17] ));
 sg13g2_dfrbp_1 _8767_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net391),
    .D(net770),
    .Q_N(_4194_),
    .Q(\btn_down_debounce.debounced ));
 sg13g2_dfrbp_1 _8768_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net389),
    .D(_0312_),
    .Q_N(_4193_),
    .Q(\btn_left_debounce.button_sync_0 ));
 sg13g2_dfrbp_1 _8769_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net388),
    .D(_0313_),
    .Q_N(_0173_),
    .Q(\btn_left_debounce.debounce_counter[0] ));
 sg13g2_dfrbp_1 _8770_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net387),
    .D(_0314_),
    .Q_N(_4192_),
    .Q(\btn_left_debounce.debounce_counter[1] ));
 sg13g2_dfrbp_1 _8771_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net386),
    .D(net506),
    .Q_N(_4191_),
    .Q(\btn_left_debounce.debounce_counter[2] ));
 sg13g2_dfrbp_1 _8772_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net385),
    .D(_0316_),
    .Q_N(_4190_),
    .Q(\btn_left_debounce.debounce_counter[3] ));
 sg13g2_dfrbp_1 _8773_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net384),
    .D(_0317_),
    .Q_N(_4189_),
    .Q(\btn_left_debounce.debounce_counter[4] ));
 sg13g2_dfrbp_1 _8774_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net383),
    .D(net791),
    .Q_N(_4188_),
    .Q(\btn_left_debounce.debounce_counter[5] ));
 sg13g2_dfrbp_1 _8775_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net382),
    .D(_0319_),
    .Q_N(_4187_),
    .Q(\btn_left_debounce.debounce_counter[6] ));
 sg13g2_dfrbp_1 _8776_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net381),
    .D(_0320_),
    .Q_N(_4186_),
    .Q(\btn_left_debounce.debounce_counter[7] ));
 sg13g2_dfrbp_1 _8777_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net380),
    .D(_0321_),
    .Q_N(_4185_),
    .Q(\btn_left_debounce.debounce_counter[8] ));
 sg13g2_dfrbp_1 _8778_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net379),
    .D(net847),
    .Q_N(_4184_),
    .Q(\btn_left_debounce.debounce_counter[9] ));
 sg13g2_dfrbp_1 _8779_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net378),
    .D(net512),
    .Q_N(_4183_),
    .Q(\btn_left_debounce.debounce_counter[10] ));
 sg13g2_dfrbp_1 _8780_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net377),
    .D(_0324_),
    .Q_N(_4182_),
    .Q(\btn_left_debounce.debounce_counter[11] ));
 sg13g2_dfrbp_1 _8781_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net376),
    .D(net629),
    .Q_N(_4181_),
    .Q(\btn_left_debounce.debounce_counter[12] ));
 sg13g2_dfrbp_1 _8782_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net375),
    .D(_0326_),
    .Q_N(_4180_),
    .Q(\btn_left_debounce.debounce_counter[13] ));
 sg13g2_dfrbp_1 _8783_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net310),
    .D(_0327_),
    .Q_N(_4179_),
    .Q(\btn_left_debounce.debounce_counter[14] ));
 sg13g2_dfrbp_1 _8784_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net309),
    .D(_0328_),
    .Q_N(_4178_),
    .Q(\btn_left_debounce.debounce_counter[15] ));
 sg13g2_dfrbp_1 _8785_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net308),
    .D(_0329_),
    .Q_N(_4177_),
    .Q(\btn_left_debounce.debounce_counter[16] ));
 sg13g2_dfrbp_1 _8786_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net307),
    .D(net744),
    .Q_N(_4176_),
    .Q(\btn_left_debounce.debounce_counter[17] ));
 sg13g2_dfrbp_1 _8787_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net306),
    .D(_0331_),
    .Q_N(_4175_),
    .Q(\btn_down_debounce.button_sync_1 ));
 sg13g2_dfrbp_1 _8788_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net305),
    .D(net824),
    .Q_N(_4174_),
    .Q(\btn_left_debounce.debounced ));
 sg13g2_dfrbp_1 _8789_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net303),
    .D(_0333_),
    .Q_N(_4173_),
    .Q(\btn_right_debounce.button_sync_0 ));
 sg13g2_dfrbp_1 _8790_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net302),
    .D(_0334_),
    .Q_N(_0172_),
    .Q(\btn_right_debounce.debounce_counter[0] ));
 sg13g2_dfrbp_1 _8791_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net301),
    .D(net833),
    .Q_N(_4172_),
    .Q(\btn_right_debounce.debounce_counter[1] ));
 sg13g2_dfrbp_1 _8792_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net300),
    .D(net583),
    .Q_N(_4171_),
    .Q(\btn_right_debounce.debounce_counter[2] ));
 sg13g2_dfrbp_1 _8793_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net299),
    .D(net789),
    .Q_N(_4170_),
    .Q(\btn_right_debounce.debounce_counter[3] ));
 sg13g2_dfrbp_1 _8794_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net298),
    .D(net752),
    .Q_N(_4169_),
    .Q(\btn_right_debounce.debounce_counter[4] ));
 sg13g2_dfrbp_1 _8795_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net294),
    .D(net761),
    .Q_N(_4168_),
    .Q(\btn_right_debounce.debounce_counter[5] ));
 sg13g2_dfrbp_1 _8796_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net293),
    .D(net749),
    .Q_N(_4167_),
    .Q(\btn_right_debounce.debounce_counter[6] ));
 sg13g2_dfrbp_1 _8797_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net292),
    .D(net812),
    .Q_N(_4166_),
    .Q(\btn_right_debounce.debounce_counter[7] ));
 sg13g2_dfrbp_1 _8798_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net291),
    .D(_0342_),
    .Q_N(_4165_),
    .Q(\btn_right_debounce.debounce_counter[8] ));
 sg13g2_dfrbp_1 _8799_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net290),
    .D(_0343_),
    .Q_N(_4164_),
    .Q(\btn_right_debounce.debounce_counter[9] ));
 sg13g2_dfrbp_1 _8800_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net289),
    .D(net568),
    .Q_N(_4163_),
    .Q(\btn_right_debounce.debounce_counter[10] ));
 sg13g2_dfrbp_1 _8801_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net288),
    .D(_0345_),
    .Q_N(_4162_),
    .Q(\btn_right_debounce.debounce_counter[11] ));
 sg13g2_dfrbp_1 _8802_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net287),
    .D(net672),
    .Q_N(_4161_),
    .Q(\btn_right_debounce.debounce_counter[12] ));
 sg13g2_dfrbp_1 _8803_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net286),
    .D(net777),
    .Q_N(_4160_),
    .Q(\btn_right_debounce.debounce_counter[13] ));
 sg13g2_dfrbp_1 _8804_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net285),
    .D(_0348_),
    .Q_N(_4159_),
    .Q(\btn_right_debounce.debounce_counter[14] ));
 sg13g2_dfrbp_1 _8805_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net284),
    .D(net688),
    .Q_N(_4158_),
    .Q(\btn_right_debounce.debounce_counter[15] ));
 sg13g2_dfrbp_1 _8806_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net283),
    .D(net590),
    .Q_N(_4157_),
    .Q(\btn_right_debounce.debounce_counter[16] ));
 sg13g2_dfrbp_1 _8807_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net282),
    .D(net461),
    .Q_N(_4156_),
    .Q(\btn_right_debounce.debounce_counter[17] ));
 sg13g2_dfrbp_1 _8808_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net281),
    .D(_0352_),
    .Q_N(_4155_),
    .Q(\btn_left_debounce.button_sync_1 ));
 sg13g2_dfrbp_1 _8809_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net280),
    .D(net686),
    .Q_N(_4154_),
    .Q(\btn_right_debounce.debounced ));
 sg13g2_dfrbp_1 _8810_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net205),
    .D(_0354_),
    .Q_N(_4308_),
    .Q(\game_logic_inst.prev_any_button_pressed ));
 sg13g2_dfrbp_1 _8811_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net254),
    .D(net416),
    .Q_N(_4309_),
    .Q(\gamepad_pmod.driver.pmod_clk_prev ));
 sg13g2_dfrbp_1 _8812_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net278),
    .D(net417),
    .Q_N(_4153_),
    .Q(\gamepad_pmod.driver.pmod_latch_prev ));
 sg13g2_dfrbp_1 _8813_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net277),
    .D(net487),
    .Q_N(_4152_),
    .Q(\gamepad_pmod.driver.shift_reg[0] ));
 sg13g2_dfrbp_1 _8814_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net275),
    .D(net715),
    .Q_N(_4151_),
    .Q(\gamepad_pmod.driver.shift_reg[1] ));
 sg13g2_dfrbp_1 _8815_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net273),
    .D(net786),
    .Q_N(_4150_),
    .Q(\gamepad_pmod.driver.shift_reg[2] ));
 sg13g2_dfrbp_1 _8816_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net271),
    .D(net772),
    .Q_N(_4149_),
    .Q(\gamepad_pmod.driver.shift_reg[3] ));
 sg13g2_dfrbp_1 _8817_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net269),
    .D(_0359_),
    .Q_N(_4148_),
    .Q(\gamepad_pmod.driver.shift_reg[4] ));
 sg13g2_dfrbp_1 _8818_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net267),
    .D(_0360_),
    .Q_N(_4147_),
    .Q(\gamepad_pmod.driver.shift_reg[5] ));
 sg13g2_dfrbp_1 _8819_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net264),
    .D(net663),
    .Q_N(_4146_),
    .Q(\gamepad_pmod.driver.shift_reg[6] ));
 sg13g2_dfrbp_1 _8820_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net262),
    .D(_0362_),
    .Q_N(_4145_),
    .Q(\gamepad_pmod.driver.shift_reg[7] ));
 sg13g2_dfrbp_1 _8821_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net260),
    .D(net478),
    .Q_N(_4144_),
    .Q(\gamepad_pmod.driver.shift_reg[8] ));
 sg13g2_dfrbp_1 _8822_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net258),
    .D(net774),
    .Q_N(_4143_),
    .Q(\gamepad_pmod.driver.shift_reg[9] ));
 sg13g2_dfrbp_1 _8823_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net256),
    .D(net767),
    .Q_N(_4142_),
    .Q(\gamepad_pmod.driver.shift_reg[10] ));
 sg13g2_dfrbp_1 _8824_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net253),
    .D(net626),
    .Q_N(_4141_),
    .Q(\gamepad_pmod.driver.shift_reg[11] ));
 sg13g2_dfrbp_1 _8825_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net251),
    .D(_0367_),
    .Q_N(_4140_),
    .Q(\gamepad_pmod.driver.pmod_data_sync[0] ));
 sg13g2_dfrbp_1 _8826_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net250),
    .D(_0368_),
    .Q_N(_4139_),
    .Q(\gamepad_pmod.driver.pmod_data_sync[1] ));
 sg13g2_dfrbp_1 _8827_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net249),
    .D(_0369_),
    .Q_N(_4138_),
    .Q(\gamepad_pmod.driver.pmod_clk_sync[0] ));
 sg13g2_dfrbp_1 _8828_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net248),
    .D(_0370_),
    .Q_N(_4137_),
    .Q(\gamepad_pmod.driver.pmod_clk_sync[1] ));
 sg13g2_dfrbp_1 _8829_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net247),
    .D(_0371_),
    .Q_N(_4136_),
    .Q(\game_logic_inst.lfsr_value[0] ));
 sg13g2_dfrbp_1 _8830_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net246),
    .D(_0372_),
    .Q_N(_4135_),
    .Q(\game_logic_inst.lfsr_value[1] ));
 sg13g2_dfrbp_1 _8831_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net245),
    .D(_0373_),
    .Q_N(_4134_),
    .Q(\game_logic_inst.lfsr_value[2] ));
 sg13g2_dfrbp_1 _8832_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net244),
    .D(_0374_),
    .Q_N(_4133_),
    .Q(\game_logic_inst.lfsr_value[3] ));
 sg13g2_dfrbp_1 _8833_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net243),
    .D(_0375_),
    .Q_N(_4132_),
    .Q(\game_logic_inst.lfsr_value[4] ));
 sg13g2_dfrbp_1 _8834_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net242),
    .D(_0376_),
    .Q_N(_4131_),
    .Q(\game_logic_inst.lfsr_value[5] ));
 sg13g2_dfrbp_1 _8835_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net241),
    .D(_0377_),
    .Q_N(_4130_),
    .Q(\game_logic_inst.lfsr_value[6] ));
 sg13g2_dfrbp_1 _8836_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net240),
    .D(_0378_),
    .Q_N(_4129_),
    .Q(\game_logic_inst.lfsr_value[7] ));
 sg13g2_dfrbp_1 _8837_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net239),
    .D(_0379_),
    .Q_N(_4128_),
    .Q(\game_logic_inst.lfsr_value[8] ));
 sg13g2_dfrbp_1 _8838_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net238),
    .D(_0380_),
    .Q_N(_4127_),
    .Q(\game_logic_inst.lfsr_value[9] ));
 sg13g2_dfrbp_1 _8839_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net237),
    .D(_0381_),
    .Q_N(_4126_),
    .Q(\game_logic_inst.lfsr_value[10] ));
 sg13g2_dfrbp_1 _8840_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net236),
    .D(_0382_),
    .Q_N(_4125_),
    .Q(\game_logic_inst.lfsr_value[11] ));
 sg13g2_dfrbp_1 _8841_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net235),
    .D(_0383_),
    .Q_N(_4124_),
    .Q(\game_logic_inst.lfsr_value[12] ));
 sg13g2_dfrbp_1 _8842_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net234),
    .D(_0384_),
    .Q_N(_4123_),
    .Q(\game_logic_inst.lfsr_value[13] ));
 sg13g2_dfrbp_1 _8843_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net233),
    .D(_0385_),
    .Q_N(_4122_),
    .Q(\game_logic_inst.lfsr_value[14] ));
 sg13g2_dfrbp_1 _8844_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net232),
    .D(_0386_),
    .Q_N(_4121_),
    .Q(\game_logic_inst.lfsr_value[15] ));
 sg13g2_dfrbp_1 _8845_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net231),
    .D(_0387_),
    .Q_N(_4120_),
    .Q(\lfsr_inst.lfsr[16] ));
 sg13g2_dfrbp_1 _8846_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net230),
    .D(_0388_),
    .Q_N(_4119_),
    .Q(\lfsr_inst.lfsr[17] ));
 sg13g2_dfrbp_1 _8847_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net229),
    .D(_0389_),
    .Q_N(_4118_),
    .Q(\lfsr_inst.lfsr[18] ));
 sg13g2_dfrbp_1 _8848_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net228),
    .D(_0390_),
    .Q_N(_4117_),
    .Q(\lfsr_inst.lfsr[19] ));
 sg13g2_dfrbp_1 _8849_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net227),
    .D(_0391_),
    .Q_N(_4116_),
    .Q(\lfsr_inst.lfsr[20] ));
 sg13g2_dfrbp_1 _8850_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net226),
    .D(_0392_),
    .Q_N(_4115_),
    .Q(\lfsr_inst.lfsr[21] ));
 sg13g2_dfrbp_1 _8851_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net225),
    .D(_0393_),
    .Q_N(_4114_),
    .Q(\lfsr_inst.lfsr[22] ));
 sg13g2_dfrbp_1 _8852_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net224),
    .D(_0394_),
    .Q_N(_4113_),
    .Q(\lfsr_inst.lfsr[23] ));
 sg13g2_dfrbp_1 _8853_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net223),
    .D(_0395_),
    .Q_N(_4112_),
    .Q(\lfsr_inst.lfsr[24] ));
 sg13g2_dfrbp_1 _8854_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net222),
    .D(_0396_),
    .Q_N(_4111_),
    .Q(\lfsr_inst.lfsr[25] ));
 sg13g2_dfrbp_1 _8855_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net221),
    .D(_0397_),
    .Q_N(_4110_),
    .Q(\lfsr_inst.lfsr[26] ));
 sg13g2_dfrbp_1 _8856_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net220),
    .D(_0398_),
    .Q_N(_4109_),
    .Q(\lfsr_inst.lfsr[27] ));
 sg13g2_dfrbp_1 _8857_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net219),
    .D(_0399_),
    .Q_N(_4108_),
    .Q(\lfsr_inst.lfsr[28] ));
 sg13g2_dfrbp_1 _8858_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net218),
    .D(_0400_),
    .Q_N(_4107_),
    .Q(\lfsr_inst.lfsr[29] ));
 sg13g2_dfrbp_1 _8859_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net217),
    .D(_0401_),
    .Q_N(_0167_),
    .Q(\lfsr_inst.lfsr[30] ));
 sg13g2_dfrbp_1 _8860_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net265),
    .D(_0402_),
    .Q_N(_4310_),
    .Q(\lfsr_inst.lfsr[31] ));
 sg13g2_dfrbp_1 _8861_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net216),
    .D(_0067_),
    .Q_N(_4106_),
    .Q(hsync));
 sg13g2_dfrbp_1 _8862_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net215),
    .D(_0403_),
    .Q_N(_0171_),
    .Q(\draw_game_inst.board_y[0] ));
 sg13g2_dfrbp_1 _8863_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net213),
    .D(_0404_),
    .Q_N(_0093_),
    .Q(\draw_game_inst.board_y[1] ));
 sg13g2_dfrbp_1 _8864_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net211),
    .D(_0405_),
    .Q_N(_0092_),
    .Q(\draw_game_inst.board_y[2] ));
 sg13g2_dfrbp_1 _8865_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net209),
    .D(_0406_),
    .Q_N(_0091_),
    .Q(\draw_game_inst.board_y[3] ));
 sg13g2_dfrbp_1 _8866_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net207),
    .D(_0407_),
    .Q_N(_0090_),
    .Q(\draw_game_inst.board_y[4] ));
 sg13g2_dfrbp_1 _8867_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net203),
    .D(_0408_),
    .Q_N(_4105_),
    .Q(\draw_game_inst.board_y[5] ));
 sg13g2_dfrbp_1 _8868_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net194),
    .D(_0409_),
    .Q_N(_0089_),
    .Q(\draw_game_inst.board_y[6] ));
 sg13g2_dfrbp_1 _8869_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net190),
    .D(_0410_),
    .Q_N(_0088_),
    .Q(\draw_game_inst.y[7] ));
 sg13g2_dfrbp_1 _8870_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net186),
    .D(_0411_),
    .Q_N(_4104_),
    .Q(\draw_game_inst.y[8] ));
 sg13g2_dfrbp_1 _8871_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net295),
    .D(_0412_),
    .Q_N(_4311_),
    .Q(\draw_game_inst.y[9] ));
 sg13g2_dfrbp_1 _8872_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net182),
    .D(_0068_),
    .Q_N(_4103_),
    .Q(\vga_sync_gen.vsync ));
 sg13g2_dfrbp_1 _8873_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net178),
    .D(_0413_),
    .Q_N(_4102_),
    .Q(\gamepad_pmod.driver.pmod_latch_sync[0] ));
 sg13g2_dfrbp_1 _8874_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net176),
    .D(_0414_),
    .Q_N(_4101_),
    .Q(\gamepad_pmod.driver.pmod_latch_sync[1] ));
 sg13g2_dfrbp_1 _8875_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net174),
    .D(net551),
    .Q_N(_4100_),
    .Q(\gamepad_pmod.decoder.data_reg[0] ));
 sg13g2_dfrbp_1 _8876_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net170),
    .D(net498),
    .Q_N(_4099_),
    .Q(\gamepad_pmod.decoder.data_reg[1] ));
 sg13g2_dfrbp_1 _8877_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net166),
    .D(net466),
    .Q_N(_4098_),
    .Q(\gamepad_pmod.decoder.data_reg[2] ));
 sg13g2_dfrbp_1 _8878_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net162),
    .D(net470),
    .Q_N(_4097_),
    .Q(\gamepad_pmod.decoder.data_reg[3] ));
 sg13g2_dfrbp_1 _8879_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net158),
    .D(net649),
    .Q_N(_4096_),
    .Q(\gamepad_pmod.decoder.data_reg[4] ));
 sg13g2_dfrbp_1 _8880_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net154),
    .D(_0420_),
    .Q_N(_4095_),
    .Q(\gamepad_pmod.decoder.data_reg[5] ));
 sg13g2_dfrbp_1 _8881_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net150),
    .D(net678),
    .Q_N(_4094_),
    .Q(\gamepad_pmod.decoder.data_reg[6] ));
 sg13g2_dfrbp_1 _8882_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net146),
    .D(_0422_),
    .Q_N(_4093_),
    .Q(\gamepad_pmod.decoder.data_reg[7] ));
 sg13g2_dfrbp_1 _8883_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net142),
    .D(net759),
    .Q_N(_4092_),
    .Q(\gamepad_pmod.decoder.data_reg[8] ));
 sg13g2_dfrbp_1 _8884_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net138),
    .D(net704),
    .Q_N(_4091_),
    .Q(\gamepad_pmod.decoder.data_reg[9] ));
 sg13g2_dfrbp_1 _8885_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net134),
    .D(net532),
    .Q_N(_4090_),
    .Q(\gamepad_pmod.decoder.data_reg[10] ));
 sg13g2_dfrbp_1 _8886_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net130),
    .D(net468),
    .Q_N(_4089_),
    .Q(\gamepad_pmod.decoder.data_reg[11] ));
 sg13g2_dfrbp_1 _8887_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net126),
    .D(_0427_),
    .Q_N(_0170_),
    .Q(\draw_game_inst.board_x[0] ));
 sg13g2_dfrbp_1 _8888_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net124),
    .D(net999),
    .Q_N(_4088_),
    .Q(\draw_game_inst.board_x[1] ));
 sg13g2_dfrbp_1 _8889_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net122),
    .D(net830),
    .Q_N(_4087_),
    .Q(\draw_game_inst.board_x[2] ));
 sg13g2_dfrbp_1 _8890_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net120),
    .D(_0430_),
    .Q_N(_0095_),
    .Q(\draw_game_inst.board_x[3] ));
 sg13g2_dfrbp_1 _8891_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net118),
    .D(_0431_),
    .Q_N(_0096_),
    .Q(\draw_game_inst.board_x[4] ));
 sg13g2_dfrbp_1 _8892_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net116),
    .D(_0432_),
    .Q_N(_0094_),
    .Q(\draw_game_inst.board_x[5] ));
 sg13g2_dfrbp_1 _8893_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net114),
    .D(_0433_),
    .Q_N(_4086_),
    .Q(\draw_game_inst.x[6] ));
 sg13g2_dfrbp_1 _8894_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net112),
    .D(_0434_),
    .Q_N(_4085_),
    .Q(\draw_game_inst.x[7] ));
 sg13g2_dfrbp_1 _8895_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net110),
    .D(_0435_),
    .Q_N(_4084_),
    .Q(\draw_game_inst.x[8] ));
 sg13g2_dfrbp_1 _8896_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net108),
    .D(_0436_),
    .Q_N(_4083_),
    .Q(\draw_game_inst.x[9] ));
 sg13g2_dfrbp_1 _8897_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net106),
    .D(_0437_),
    .Q_N(_4082_),
    .Q(\welcome_screen_inst.welcome_counter[0] ));
 sg13g2_dfrbp_1 _8898_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net102),
    .D(net803),
    .Q_N(_4081_),
    .Q(\welcome_screen_inst.welcome_counter[1] ));
 sg13g2_dfrbp_1 _8899_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net98),
    .D(net805),
    .Q_N(_4080_),
    .Q(\welcome_screen_inst.welcome_counter[2] ));
 sg13g2_dfrbp_1 _8900_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net94),
    .D(_0440_),
    .Q_N(_4079_),
    .Q(\welcome_screen_inst.welcome_counter[3] ));
 sg13g2_dfrbp_1 _8901_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net296),
    .D(net836),
    .Q_N(_4312_),
    .Q(\welcome_screen_inst.welcome_counter[4] ));
 sg13g2_dfrbp_1 _8902_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net297),
    .D(net635),
    .Q_N(_4313_),
    .Q(\game_logic_inst.current_direction[1] ));
 sg13g2_dfrbp_1 _8903_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net311),
    .D(net956),
    .Q_N(_4314_),
    .Q(\game_logic_inst.current_direction[2] ));
 sg13g2_dfrbp_1 _8904_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net90),
    .D(_0002_),
    .Q_N(_4078_),
    .Q(\game_logic_inst.current_direction[3] ));
 sg13g2_dfrbp_1 _8905_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net86),
    .D(net828),
    .Q_N(_4077_),
    .Q(\game_logic_inst.debug_move_reg ));
 sg13g2_dfrbp_1 _8906_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net82),
    .D(_0443_),
    .Q_N(_4076_),
    .Q(\game_logic_inst.valid_move ));
 sg13g2_dfrbp_1 _8907_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net78),
    .D(_0444_),
    .Q_N(_0097_),
    .Q(\game_logic_inst.calculate_move ));
 sg13g2_dfrbp_1 _8908_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net74),
    .D(_0445_),
    .Q_N(_0169_),
    .Q(\game_logic_inst.lfsr_shift[0] ));
 sg13g2_dfrbp_1 _8909_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net72),
    .D(_0446_),
    .Q_N(_4075_),
    .Q(\game_logic_inst.lfsr_shift[1] ));
 sg13g2_dfrbp_1 _8910_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net70),
    .D(_0447_),
    .Q_N(_0166_),
    .Q(\game_logic_inst.game_started ));
 sg13g2_dfrbp_1 _8911_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net68),
    .D(net797),
    .Q_N(_4074_),
    .Q(\game_logic_inst.add_new_tiles[0] ));
 sg13g2_dfrbp_1 _8912_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net42),
    .D(net442),
    .Q_N(_4073_),
    .Q(\game_logic_inst.add_new_tiles[1] ));
 sg13g2_dfrbp_1 _8913_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net390),
    .D(_0450_),
    .Q_N(_4072_),
    .Q(\game_logic_inst.added_tile_index[0] ));
 sg13g2_dfrbp_1 _8914_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net304),
    .D(_0451_),
    .Q_N(_4071_),
    .Q(\game_logic_inst.added_tile_index[1] ));
 sg13g2_dfrbp_1 _8915_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net279),
    .D(_0452_),
    .Q_N(_4070_),
    .Q(\game_logic_inst.added_tile_index[2] ));
 sg13g2_dfrbp_1 _8916_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net276),
    .D(_0453_),
    .Q_N(_4069_),
    .Q(\game_logic_inst.added_tile_index[3] ));
 sg13g2_dfrbp_1 _8917_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net312),
    .D(_0454_),
    .Q_N(_4315_),
    .Q(\debug_controller_inst.data_out_en ));
 sg13g2_dfrbp_1 _8918_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net313),
    .D(net960),
    .Q_N(_0099_),
    .Q(\debug_controller_inst.grid_in[0] ));
 sg13g2_dfrbp_1 _8919_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net314),
    .D(net938),
    .Q_N(_0100_),
    .Q(\debug_controller_inst.grid_in[1] ));
 sg13g2_dfrbp_1 _8920_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net315),
    .D(net929),
    .Q_N(_0101_),
    .Q(\debug_controller_inst.grid_in[2] ));
 sg13g2_dfrbp_1 _8921_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net316),
    .D(net906),
    .Q_N(_0102_),
    .Q(\debug_controller_inst.grid_in[3] ));
 sg13g2_dfrbp_1 _8922_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net317),
    .D(_0047_),
    .Q_N(_0103_),
    .Q(\debug_controller_inst.grid_in[4] ));
 sg13g2_dfrbp_1 _8923_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net318),
    .D(_0058_),
    .Q_N(_0105_),
    .Q(\debug_controller_inst.grid_in[5] ));
 sg13g2_dfrbp_1 _8924_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net319),
    .D(_0063_),
    .Q_N(_0107_),
    .Q(\debug_controller_inst.grid_in[6] ));
 sg13g2_dfrbp_1 _8925_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net320),
    .D(_0064_),
    .Q_N(_0109_),
    .Q(\debug_controller_inst.grid_in[7] ));
 sg13g2_dfrbp_1 _8926_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net321),
    .D(net904),
    .Q_N(_0111_),
    .Q(\debug_controller_inst.grid_in[8] ));
 sg13g2_dfrbp_1 _8927_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net322),
    .D(net921),
    .Q_N(_0113_),
    .Q(\debug_controller_inst.grid_in[9] ));
 sg13g2_dfrbp_1 _8928_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net323),
    .D(net969),
    .Q_N(_0115_),
    .Q(\debug_controller_inst.grid_in[10] ));
 sg13g2_dfrbp_1 _8929_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net324),
    .D(net944),
    .Q_N(_0117_),
    .Q(\debug_controller_inst.grid_in[11] ));
 sg13g2_dfrbp_1 _8930_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net325),
    .D(_0006_),
    .Q_N(_0119_),
    .Q(\debug_controller_inst.grid_in[12] ));
 sg13g2_dfrbp_1 _8931_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net326),
    .D(_0007_),
    .Q_N(_0121_),
    .Q(\debug_controller_inst.grid_in[13] ));
 sg13g2_dfrbp_1 _8932_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net327),
    .D(_0008_),
    .Q_N(_0123_),
    .Q(\debug_controller_inst.grid_in[14] ));
 sg13g2_dfrbp_1 _8933_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net328),
    .D(_0009_),
    .Q_N(_0125_),
    .Q(\debug_controller_inst.grid_in[15] ));
 sg13g2_dfrbp_1 _8934_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net329),
    .D(_0010_),
    .Q_N(_0104_),
    .Q(\debug_controller_inst.grid_in[16] ));
 sg13g2_dfrbp_1 _8935_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net330),
    .D(_0011_),
    .Q_N(_0106_),
    .Q(\debug_controller_inst.grid_in[17] ));
 sg13g2_dfrbp_1 _8936_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net331),
    .D(_0012_),
    .Q_N(_0108_),
    .Q(\debug_controller_inst.grid_in[18] ));
 sg13g2_dfrbp_1 _8937_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net332),
    .D(_0013_),
    .Q_N(_0110_),
    .Q(\debug_controller_inst.grid_in[19] ));
 sg13g2_dfrbp_1 _8938_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net333),
    .D(_0015_),
    .Q_N(_0127_),
    .Q(\debug_controller_inst.grid_in[20] ));
 sg13g2_dfrbp_1 _8939_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net334),
    .D(_0016_),
    .Q_N(_0128_),
    .Q(\debug_controller_inst.grid_in[21] ));
 sg13g2_dfrbp_1 _8940_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net335),
    .D(_0017_),
    .Q_N(_0129_),
    .Q(\debug_controller_inst.grid_in[22] ));
 sg13g2_dfrbp_1 _8941_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net336),
    .D(net913),
    .Q_N(_0130_),
    .Q(\debug_controller_inst.grid_in[23] ));
 sg13g2_dfrbp_1 _8942_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net337),
    .D(net964),
    .Q_N(_0131_),
    .Q(\debug_controller_inst.grid_in[24] ));
 sg13g2_dfrbp_1 _8943_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net338),
    .D(net932),
    .Q_N(_0133_),
    .Q(\debug_controller_inst.grid_in[25] ));
 sg13g2_dfrbp_1 _8944_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net339),
    .D(net979),
    .Q_N(_0135_),
    .Q(\debug_controller_inst.grid_in[26] ));
 sg13g2_dfrbp_1 _8945_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net340),
    .D(net987),
    .Q_N(_0137_),
    .Q(\debug_controller_inst.grid_in[27] ));
 sg13g2_dfrbp_1 _8946_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net341),
    .D(_0023_),
    .Q_N(_0139_),
    .Q(\debug_controller_inst.grid_in[28] ));
 sg13g2_dfrbp_1 _8947_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net342),
    .D(_0024_),
    .Q_N(_0141_),
    .Q(\debug_controller_inst.grid_in[29] ));
 sg13g2_dfrbp_1 _8948_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net343),
    .D(_0026_),
    .Q_N(_0143_),
    .Q(\debug_controller_inst.grid_in[30] ));
 sg13g2_dfrbp_1 _8949_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net344),
    .D(_0027_),
    .Q_N(_0145_),
    .Q(\debug_controller_inst.grid_in[31] ));
 sg13g2_dfrbp_1 _8950_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net345),
    .D(net990),
    .Q_N(_0112_),
    .Q(\debug_controller_inst.grid_in[32] ));
 sg13g2_dfrbp_1 _8951_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net346),
    .D(_0029_),
    .Q_N(_0114_),
    .Q(\debug_controller_inst.grid_in[33] ));
 sg13g2_dfrbp_1 _8952_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net347),
    .D(_0030_),
    .Q_N(_0116_),
    .Q(\debug_controller_inst.grid_in[34] ));
 sg13g2_dfrbp_1 _8953_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net348),
    .D(net1022),
    .Q_N(_0118_),
    .Q(\debug_controller_inst.grid_in[35] ));
 sg13g2_dfrbp_1 _8954_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net349),
    .D(_0032_),
    .Q_N(_0132_),
    .Q(\debug_controller_inst.grid_in[36] ));
 sg13g2_dfrbp_1 _8955_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net350),
    .D(_0033_),
    .Q_N(_0134_),
    .Q(\debug_controller_inst.grid_in[37] ));
 sg13g2_dfrbp_1 _8956_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net351),
    .D(_0034_),
    .Q_N(_0136_),
    .Q(\debug_controller_inst.grid_in[38] ));
 sg13g2_dfrbp_1 _8957_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net352),
    .D(net1030),
    .Q_N(_0138_),
    .Q(\debug_controller_inst.grid_in[39] ));
 sg13g2_dfrbp_1 _8958_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net353),
    .D(_0037_),
    .Q_N(_0147_),
    .Q(\debug_controller_inst.grid_in[40] ));
 sg13g2_dfrbp_1 _8959_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net354),
    .D(net934),
    .Q_N(_0148_),
    .Q(\debug_controller_inst.grid_in[41] ));
 sg13g2_dfrbp_1 _8960_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net355),
    .D(net918),
    .Q_N(_0149_),
    .Q(\debug_controller_inst.grid_in[42] ));
 sg13g2_dfrbp_1 _8961_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net356),
    .D(net923),
    .Q_N(_0150_),
    .Q(\debug_controller_inst.grid_in[43] ));
 sg13g2_dfrbp_1 _8962_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net357),
    .D(net992),
    .Q_N(_0151_),
    .Q(\debug_controller_inst.grid_in[44] ));
 sg13g2_dfrbp_1 _8963_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net358),
    .D(net941),
    .Q_N(_0153_),
    .Q(\debug_controller_inst.grid_in[45] ));
 sg13g2_dfrbp_1 _8964_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net359),
    .D(net984),
    .Q_N(_0155_),
    .Q(\debug_controller_inst.grid_in[46] ));
 sg13g2_dfrbp_1 _8965_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net360),
    .D(_0044_),
    .Q_N(_0157_),
    .Q(\debug_controller_inst.grid_in[47] ));
 sg13g2_dfrbp_1 _8966_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net361),
    .D(_0045_),
    .Q_N(_0120_),
    .Q(\debug_controller_inst.grid_in[48] ));
 sg13g2_dfrbp_1 _8967_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net362),
    .D(_0046_),
    .Q_N(_0122_),
    .Q(\debug_controller_inst.grid_in[49] ));
 sg13g2_dfrbp_1 _8968_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net363),
    .D(_0048_),
    .Q_N(_0124_),
    .Q(\debug_controller_inst.grid_in[50] ));
 sg13g2_dfrbp_1 _8969_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net364),
    .D(_0049_),
    .Q_N(_0126_),
    .Q(\debug_controller_inst.grid_in[51] ));
 sg13g2_dfrbp_1 _8970_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net365),
    .D(_0050_),
    .Q_N(_0140_),
    .Q(\debug_controller_inst.grid_in[52] ));
 sg13g2_dfrbp_1 _8971_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net366),
    .D(net899),
    .Q_N(_0142_),
    .Q(\debug_controller_inst.grid_in[53] ));
 sg13g2_dfrbp_1 _8972_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net367),
    .D(net972),
    .Q_N(_0144_),
    .Q(\debug_controller_inst.grid_in[54] ));
 sg13g2_dfrbp_1 _8973_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net368),
    .D(_0053_),
    .Q_N(_0146_),
    .Q(\debug_controller_inst.grid_in[55] ));
 sg13g2_dfrbp_1 _8974_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net369),
    .D(_0054_),
    .Q_N(_0152_),
    .Q(\debug_controller_inst.grid_in[56] ));
 sg13g2_dfrbp_1 _8975_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net370),
    .D(_0055_),
    .Q_N(_0154_),
    .Q(\debug_controller_inst.grid_in[57] ));
 sg13g2_dfrbp_1 _8976_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net371),
    .D(net910),
    .Q_N(_0156_),
    .Q(\debug_controller_inst.grid_in[58] ));
 sg13g2_dfrbp_1 _8977_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net372),
    .D(net976),
    .Q_N(_0158_),
    .Q(\debug_controller_inst.grid_in[59] ));
 sg13g2_dfrbp_1 _8978_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net373),
    .D(_0059_),
    .Q_N(_0159_),
    .Q(\debug_controller_inst.grid_in[60] ));
 sg13g2_dfrbp_1 _8979_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net374),
    .D(_0060_),
    .Q_N(_0160_),
    .Q(\debug_controller_inst.grid_in[61] ));
 sg13g2_dfrbp_1 _8980_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net257),
    .D(_0061_),
    .Q_N(_0161_),
    .Q(\debug_controller_inst.grid_in[62] ));
 sg13g2_dfrbp_1 _8981_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net274),
    .D(_0062_),
    .Q_N(_0162_),
    .Q(\debug_controller_inst.grid_in[63] ));
 sg13g2_dfrbp_1 _8982_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net272),
    .D(net888),
    .Q_N(_0069_),
    .Q(\game_logic_inst.should_transpose ));
 sg13g2_dfrbp_1 _8983_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net268),
    .D(_0456_),
    .Q_N(_0098_),
    .Q(\game_logic_inst.current_row_index[0] ));
 sg13g2_dfrbp_1 _8984_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net263),
    .D(net916),
    .Q_N(_4068_),
    .Q(\game_logic_inst.current_row_index[1] ));
 sg13g2_dfrbp_1 _8985_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net259),
    .D(_0458_),
    .Q_N(_4067_),
    .Q(uio_out[4]));
 sg13g2_dfrbp_1 _8986_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net255),
    .D(_0459_),
    .Q_N(_4066_),
    .Q(uio_out[5]));
 sg13g2_dfrbp_1 _8987_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net214),
    .D(_0460_),
    .Q_N(_4065_),
    .Q(uio_out[6]));
 sg13g2_dfrbp_1 _8988_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net210),
    .D(_0461_),
    .Q_N(_4064_),
    .Q(uio_out[7]));
 sg13g2_dfrbp_1 _8989_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net206),
    .D(_0462_),
    .Q_N(_4063_),
    .Q(debug_btn_up));
 sg13g2_dfrbp_1 _8990_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net202),
    .D(_0463_),
    .Q_N(_4062_),
    .Q(debug_btn_down));
 sg13g2_dfrbp_1 _8991_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net192),
    .D(_0464_),
    .Q_N(_4061_),
    .Q(debug_btn_left));
 sg13g2_dfrbp_1 _8992_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net188),
    .D(_0465_),
    .Q_N(_4060_),
    .Q(debug_btn_right));
 sg13g2_dfrbp_1 _8993_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net184),
    .D(_0466_),
    .Q_N(_4059_),
    .Q(\debug_controller_inst.grid_out_valid ));
 sg13g2_dfrbp_1 _8994_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net180),
    .D(_0467_),
    .Q_N(_4058_),
    .Q(\debug_controller_inst.grid_out_data[0] ));
 sg13g2_dfrbp_1 _8995_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net168),
    .D(_0468_),
    .Q_N(_4057_),
    .Q(\debug_controller_inst.grid_out_data[1] ));
 sg13g2_dfrbp_1 _8996_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net160),
    .D(_0469_),
    .Q_N(_4056_),
    .Q(\debug_controller_inst.grid_out_data[2] ));
 sg13g2_dfrbp_1 _8997_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net152),
    .D(_0470_),
    .Q_N(_4055_),
    .Q(\debug_controller_inst.grid_out_data[3] ));
 sg13g2_dfrbp_1 _8998_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net144),
    .D(_0471_),
    .Q_N(_4054_),
    .Q(\debug_controller_inst.grid_out_addr[0] ));
 sg13g2_dfrbp_1 _8999_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net136),
    .D(_0472_),
    .Q_N(_4053_),
    .Q(\debug_controller_inst.grid_out_addr[1] ));
 sg13g2_dfrbp_1 _9000_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net128),
    .D(net952),
    .Q_N(_4052_),
    .Q(\debug_controller_inst.grid_out_addr[2] ));
 sg13g2_dfrbp_1 _9001_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net100),
    .D(_0474_),
    .Q_N(_4051_),
    .Q(\debug_controller_inst.grid_out_addr[3] ));
 sg13g2_dfrbp_1 _9002_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net92),
    .D(_0475_),
    .Q_N(_4050_),
    .Q(\btn_up_debounce.button_sync_1 ));
 sg13g2_dfrbp_1 _9003_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net88),
    .D(net439),
    .Q_N(_0163_),
    .Q(\debug_controller_inst.grid_addr[0] ));
 sg13g2_dfrbp_1 _9004_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net80),
    .D(_0477_),
    .Q_N(_4049_),
    .Q(\debug_controller_inst.grid_addr[1] ));
 sg13g2_dfrbp_1 _9005_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net66),
    .D(_0478_),
    .Q_N(_0164_),
    .Q(\debug_controller_inst.grid_addr[2] ));
 sg13g2_dfrbp_1 _9006_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net270),
    .D(_0479_),
    .Q_N(_4048_),
    .Q(\debug_controller_inst.grid_addr[3] ));
 sg13g2_dfrbp_1 _9007_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net261),
    .D(net852),
    .Q_N(_4047_),
    .Q(\welcome_screen_grid[52] ));
 sg13g2_dfrbp_1 _9008_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net252),
    .D(net820),
    .Q_N(_4046_),
    .Q(\welcome_screen_grid[56] ));
 sg13g2_dfrbp_1 _9009_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net208),
    .D(net859),
    .Q_N(_4045_),
    .Q(\welcome_screen_grid[60] ));
 sg13g2_dfrbp_1 _9010_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net164),
    .D(net724),
    .Q_N(_4044_),
    .Q(\welcome_screen_grid[44] ));
 sg13g2_dfrbp_1 _9011_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net148),
    .D(net717),
    .Q_N(_4043_),
    .Q(\welcome_screen_grid[40] ));
 sg13g2_dfrbp_1 _9012_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net132),
    .D(net696),
    .Q_N(_4042_),
    .Q(\welcome_screen_grid[11] ));
 sg13g2_dfrbp_1 _9013_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net96),
    .D(net665),
    .Q_N(_4041_),
    .Q(\welcome_screen_grid[32] ));
 sg13g2_dfrbp_1 _9014_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net76),
    .D(net756),
    .Q_N(_4040_),
    .Q(\welcome_screen_grid[0] ));
 sg13g2_dfrbp_1 _9015_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net266),
    .D(net842),
    .Q_N(_4039_),
    .Q(\welcome_screen_grid[20] ));
 sg13g2_dfrbp_1 _9016_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net212),
    .D(net795),
    .Q_N(_4038_),
    .Q(\welcome_screen_grid[36] ));
 sg13g2_dfrbp_1 _9017_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net156),
    .D(net861),
    .Q_N(_4037_),
    .Q(\welcome_screen_grid[16] ));
 sg13g2_dfrbp_1 _9018_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net104),
    .D(net885),
    .Q_N(_4036_),
    .Q(\welcome_screen_grid[48] ));
 sg13g2_dfrbp_1 _9019_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net411),
    .D(net857),
    .Q_N(_4035_),
    .Q(\welcome_screen_grid[28] ));
 sg13g2_dfrbp_1 _9020_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net172),
    .D(net880),
    .Q_N(_4034_),
    .Q(\welcome_screen_grid[24] ));
 sg13g2_dfrbp_1 _9021_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net84),
    .D(net814),
    .Q_N(_4033_),
    .Q(\welcome_screen_grid[12] ));
 sg13g2_dfrbp_1 _9022_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net140),
    .D(net779),
    .Q_N(_4032_),
    .Q(\welcome_screen_grid[4] ));
 sg13g2_tiehi _8742__26 (.L_HI(net26));
 sg13g2_tiehi _8741__27 (.L_HI(net27));
 sg13g2_tiehi _8740__28 (.L_HI(net28));
 sg13g2_tiehi _8739__29 (.L_HI(net29));
 sg13g2_tiehi _8738__30 (.L_HI(net30));
 sg13g2_tiehi _8737__31 (.L_HI(net31));
 sg13g2_tiehi _8736__32 (.L_HI(net32));
 sg13g2_tiehi _8735__33 (.L_HI(net33));
 sg13g2_tiehi _8734__34 (.L_HI(net34));
 sg13g2_tiehi _8733__35 (.L_HI(net35));
 sg13g2_tiehi _8732__36 (.L_HI(net36));
 sg13g2_tiehi _8731__37 (.L_HI(net37));
 sg13g2_tiehi _8730__38 (.L_HI(net38));
 sg13g2_tiehi _8729__39 (.L_HI(net39));
 sg13g2_tiehi _8728__40 (.L_HI(net40));
 sg13g2_tiehi _8727__41 (.L_HI(net41));
 sg13g2_tiehi _8912__42 (.L_HI(net42));
 sg13g2_tiehi _8726__43 (.L_HI(net43));
 sg13g2_tiehi _8725__44 (.L_HI(net44));
 sg13g2_tiehi _8724__45 (.L_HI(net45));
 sg13g2_tiehi _8723__46 (.L_HI(net46));
 sg13g2_tiehi _8722__47 (.L_HI(net47));
 sg13g2_tiehi _8721__48 (.L_HI(net48));
 sg13g2_tiehi _8720__49 (.L_HI(net49));
 sg13g2_tiehi _8719__50 (.L_HI(net50));
 sg13g2_tiehi _8718__51 (.L_HI(net51));
 sg13g2_tiehi _8717__52 (.L_HI(net52));
 sg13g2_tiehi _8716__53 (.L_HI(net53));
 sg13g2_tiehi _8715__54 (.L_HI(net54));
 sg13g2_tiehi _8714__55 (.L_HI(net55));
 sg13g2_tiehi _8713__56 (.L_HI(net56));
 sg13g2_tiehi _8712__57 (.L_HI(net57));
 sg13g2_tiehi _8711__58 (.L_HI(net58));
 sg13g2_tiehi _8710__59 (.L_HI(net59));
 sg13g2_tiehi _8709__60 (.L_HI(net60));
 sg13g2_tiehi _8708__61 (.L_HI(net61));
 sg13g2_tiehi _8707__62 (.L_HI(net62));
 sg13g2_tiehi _8706__63 (.L_HI(net63));
 sg13g2_tiehi _8705__64 (.L_HI(net64));
 sg13g2_tiehi _8704__65 (.L_HI(net65));
 sg13g2_tiehi _9005__66 (.L_HI(net66));
 sg13g2_tiehi _8703__67 (.L_HI(net67));
 sg13g2_tiehi _8911__68 (.L_HI(net68));
 sg13g2_tiehi _8702__69 (.L_HI(net69));
 sg13g2_tiehi _8910__70 (.L_HI(net70));
 sg13g2_tiehi _8701__71 (.L_HI(net71));
 sg13g2_tiehi _8909__72 (.L_HI(net72));
 sg13g2_tiehi _8700__73 (.L_HI(net73));
 sg13g2_tiehi _8908__74 (.L_HI(net74));
 sg13g2_tiehi _8699__75 (.L_HI(net75));
 sg13g2_tiehi _9014__76 (.L_HI(net76));
 sg13g2_tiehi _8698__77 (.L_HI(net77));
 sg13g2_tiehi _8907__78 (.L_HI(net78));
 sg13g2_tiehi _8697__79 (.L_HI(net79));
 sg13g2_tiehi _9004__80 (.L_HI(net80));
 sg13g2_tiehi _8696__81 (.L_HI(net81));
 sg13g2_tiehi _8906__82 (.L_HI(net82));
 sg13g2_tiehi _8695__83 (.L_HI(net83));
 sg13g2_tiehi _9021__84 (.L_HI(net84));
 sg13g2_tiehi _8694__85 (.L_HI(net85));
 sg13g2_tiehi _8905__86 (.L_HI(net86));
 sg13g2_tiehi _8693__87 (.L_HI(net87));
 sg13g2_tiehi _9003__88 (.L_HI(net88));
 sg13g2_tiehi _8692__89 (.L_HI(net89));
 sg13g2_tiehi _8904__90 (.L_HI(net90));
 sg13g2_tiehi _8691__91 (.L_HI(net91));
 sg13g2_tiehi _9002__92 (.L_HI(net92));
 sg13g2_tiehi _8690__93 (.L_HI(net93));
 sg13g2_tiehi _8900__94 (.L_HI(net94));
 sg13g2_tiehi _8689__95 (.L_HI(net95));
 sg13g2_tiehi _9013__96 (.L_HI(net96));
 sg13g2_tiehi _8688__97 (.L_HI(net97));
 sg13g2_tiehi _8899__98 (.L_HI(net98));
 sg13g2_tiehi _8687__99 (.L_HI(net99));
 sg13g2_tiehi _9001__100 (.L_HI(net100));
 sg13g2_tiehi _8686__101 (.L_HI(net101));
 sg13g2_tiehi _8898__102 (.L_HI(net102));
 sg13g2_tiehi _8685__103 (.L_HI(net103));
 sg13g2_tiehi _9018__104 (.L_HI(net104));
 sg13g2_tiehi _8684__105 (.L_HI(net105));
 sg13g2_tiehi _8897__106 (.L_HI(net106));
 sg13g2_tiehi _8683__107 (.L_HI(net107));
 sg13g2_tiehi _8896__108 (.L_HI(net108));
 sg13g2_tiehi _8682__109 (.L_HI(net109));
 sg13g2_tiehi _8895__110 (.L_HI(net110));
 sg13g2_tiehi _8681__111 (.L_HI(net111));
 sg13g2_tiehi _8894__112 (.L_HI(net112));
 sg13g2_tiehi _8680__113 (.L_HI(net113));
 sg13g2_tiehi _8893__114 (.L_HI(net114));
 sg13g2_tiehi _8679__115 (.L_HI(net115));
 sg13g2_tiehi _8892__116 (.L_HI(net116));
 sg13g2_tiehi _8678__117 (.L_HI(net117));
 sg13g2_tiehi _8891__118 (.L_HI(net118));
 sg13g2_tiehi _8677__119 (.L_HI(net119));
 sg13g2_tiehi _8890__120 (.L_HI(net120));
 sg13g2_tiehi _8676__121 (.L_HI(net121));
 sg13g2_tiehi _8889__122 (.L_HI(net122));
 sg13g2_tiehi _8675__123 (.L_HI(net123));
 sg13g2_tiehi _8888__124 (.L_HI(net124));
 sg13g2_tiehi _8674__125 (.L_HI(net125));
 sg13g2_tiehi _8887__126 (.L_HI(net126));
 sg13g2_tiehi _8673__127 (.L_HI(net127));
 sg13g2_tiehi _9000__128 (.L_HI(net128));
 sg13g2_tiehi _8672__129 (.L_HI(net129));
 sg13g2_tiehi _8886__130 (.L_HI(net130));
 sg13g2_tiehi _8671__131 (.L_HI(net131));
 sg13g2_tiehi _9012__132 (.L_HI(net132));
 sg13g2_tiehi _8670__133 (.L_HI(net133));
 sg13g2_tiehi _8885__134 (.L_HI(net134));
 sg13g2_tiehi _8669__135 (.L_HI(net135));
 sg13g2_tiehi _8999__136 (.L_HI(net136));
 sg13g2_tiehi _8668__137 (.L_HI(net137));
 sg13g2_tiehi _8884__138 (.L_HI(net138));
 sg13g2_tiehi _8667__139 (.L_HI(net139));
 sg13g2_tiehi _9022__140 (.L_HI(net140));
 sg13g2_tiehi _8666__141 (.L_HI(net141));
 sg13g2_tiehi _8883__142 (.L_HI(net142));
 sg13g2_tiehi _8665__143 (.L_HI(net143));
 sg13g2_tiehi _8998__144 (.L_HI(net144));
 sg13g2_tiehi _8664__145 (.L_HI(net145));
 sg13g2_tiehi _8882__146 (.L_HI(net146));
 sg13g2_tiehi _8663__147 (.L_HI(net147));
 sg13g2_tiehi _9011__148 (.L_HI(net148));
 sg13g2_tiehi _8662__149 (.L_HI(net149));
 sg13g2_tiehi _8881__150 (.L_HI(net150));
 sg13g2_tiehi _8661__151 (.L_HI(net151));
 sg13g2_tiehi _8997__152 (.L_HI(net152));
 sg13g2_tiehi _8660__153 (.L_HI(net153));
 sg13g2_tiehi _8880__154 (.L_HI(net154));
 sg13g2_tiehi _8659__155 (.L_HI(net155));
 sg13g2_tiehi _9017__156 (.L_HI(net156));
 sg13g2_tiehi _8658__157 (.L_HI(net157));
 sg13g2_tiehi _8879__158 (.L_HI(net158));
 sg13g2_tiehi _8657__159 (.L_HI(net159));
 sg13g2_tiehi _8996__160 (.L_HI(net160));
 sg13g2_tiehi _8656__161 (.L_HI(net161));
 sg13g2_tiehi _8878__162 (.L_HI(net162));
 sg13g2_tiehi _8655__163 (.L_HI(net163));
 sg13g2_tiehi _9010__164 (.L_HI(net164));
 sg13g2_tiehi _8654__165 (.L_HI(net165));
 sg13g2_tiehi _8877__166 (.L_HI(net166));
 sg13g2_tiehi _8653__167 (.L_HI(net167));
 sg13g2_tiehi _8995__168 (.L_HI(net168));
 sg13g2_tiehi _8652__169 (.L_HI(net169));
 sg13g2_tiehi _8876__170 (.L_HI(net170));
 sg13g2_tiehi _8651__171 (.L_HI(net171));
 sg13g2_tiehi _9020__172 (.L_HI(net172));
 sg13g2_tiehi _8650__173 (.L_HI(net173));
 sg13g2_tiehi _8875__174 (.L_HI(net174));
 sg13g2_tiehi _8649__175 (.L_HI(net175));
 sg13g2_tiehi _8874__176 (.L_HI(net176));
 sg13g2_tiehi _8648__177 (.L_HI(net177));
 sg13g2_tiehi _8873__178 (.L_HI(net178));
 sg13g2_tiehi _8647__179 (.L_HI(net179));
 sg13g2_tiehi _8994__180 (.L_HI(net180));
 sg13g2_tiehi _8646__181 (.L_HI(net181));
 sg13g2_tiehi _8872__182 (.L_HI(net182));
 sg13g2_tiehi _8645__183 (.L_HI(net183));
 sg13g2_tiehi _8993__184 (.L_HI(net184));
 sg13g2_tiehi _8644__185 (.L_HI(net185));
 sg13g2_tiehi _8870__186 (.L_HI(net186));
 sg13g2_tiehi _8643__187 (.L_HI(net187));
 sg13g2_tiehi _8992__188 (.L_HI(net188));
 sg13g2_tiehi _8642__189 (.L_HI(net189));
 sg13g2_tiehi _8869__190 (.L_HI(net190));
 sg13g2_tiehi _8641__191 (.L_HI(net191));
 sg13g2_tiehi _8991__192 (.L_HI(net192));
 sg13g2_tiehi _8640__193 (.L_HI(net193));
 sg13g2_tiehi _8868__194 (.L_HI(net194));
 sg13g2_tiehi _8639__195 (.L_HI(net195));
 sg13g2_tiehi _8638__196 (.L_HI(net196));
 sg13g2_tiehi _8637__197 (.L_HI(net197));
 sg13g2_tiehi _8636__198 (.L_HI(net198));
 sg13g2_tiehi _8635__199 (.L_HI(net199));
 sg13g2_tiehi _8634__200 (.L_HI(net200));
 sg13g2_tiehi _8633__201 (.L_HI(net201));
 sg13g2_tiehi _8990__202 (.L_HI(net202));
 sg13g2_tiehi _8867__203 (.L_HI(net203));
 sg13g2_tiehi _8632__204 (.L_HI(net204));
 sg13g2_tiehi _8810__205 (.L_HI(net205));
 sg13g2_tiehi _8989__206 (.L_HI(net206));
 sg13g2_tiehi _8866__207 (.L_HI(net207));
 sg13g2_tiehi _9009__208 (.L_HI(net208));
 sg13g2_tiehi _8865__209 (.L_HI(net209));
 sg13g2_tiehi _8988__210 (.L_HI(net210));
 sg13g2_tiehi _8864__211 (.L_HI(net211));
 sg13g2_tiehi _9016__212 (.L_HI(net212));
 sg13g2_tiehi _8863__213 (.L_HI(net213));
 sg13g2_tiehi _8987__214 (.L_HI(net214));
 sg13g2_tiehi _8862__215 (.L_HI(net215));
 sg13g2_tiehi _8861__216 (.L_HI(net216));
 sg13g2_tiehi _8859__217 (.L_HI(net217));
 sg13g2_tiehi _8858__218 (.L_HI(net218));
 sg13g2_tiehi _8857__219 (.L_HI(net219));
 sg13g2_tiehi _8856__220 (.L_HI(net220));
 sg13g2_tiehi _8855__221 (.L_HI(net221));
 sg13g2_tiehi _8854__222 (.L_HI(net222));
 sg13g2_tiehi _8853__223 (.L_HI(net223));
 sg13g2_tiehi _8852__224 (.L_HI(net224));
 sg13g2_tiehi _8851__225 (.L_HI(net225));
 sg13g2_tiehi _8850__226 (.L_HI(net226));
 sg13g2_tiehi _8849__227 (.L_HI(net227));
 sg13g2_tiehi _8848__228 (.L_HI(net228));
 sg13g2_tiehi _8847__229 (.L_HI(net229));
 sg13g2_tiehi _8846__230 (.L_HI(net230));
 sg13g2_tiehi _8845__231 (.L_HI(net231));
 sg13g2_tiehi _8844__232 (.L_HI(net232));
 sg13g2_tiehi _8843__233 (.L_HI(net233));
 sg13g2_tiehi _8842__234 (.L_HI(net234));
 sg13g2_tiehi _8841__235 (.L_HI(net235));
 sg13g2_tiehi _8840__236 (.L_HI(net236));
 sg13g2_tiehi _8839__237 (.L_HI(net237));
 sg13g2_tiehi _8838__238 (.L_HI(net238));
 sg13g2_tiehi _8837__239 (.L_HI(net239));
 sg13g2_tiehi _8836__240 (.L_HI(net240));
 sg13g2_tiehi _8835__241 (.L_HI(net241));
 sg13g2_tiehi _8834__242 (.L_HI(net242));
 sg13g2_tiehi _8833__243 (.L_HI(net243));
 sg13g2_tiehi _8832__244 (.L_HI(net244));
 sg13g2_tiehi _8831__245 (.L_HI(net245));
 sg13g2_tiehi _8830__246 (.L_HI(net246));
 sg13g2_tiehi _8829__247 (.L_HI(net247));
 sg13g2_tiehi _8828__248 (.L_HI(net248));
 sg13g2_tiehi _8827__249 (.L_HI(net249));
 sg13g2_tiehi _8826__250 (.L_HI(net250));
 sg13g2_tiehi _8825__251 (.L_HI(net251));
 sg13g2_tiehi _9008__252 (.L_HI(net252));
 sg13g2_tiehi _8824__253 (.L_HI(net253));
 sg13g2_tiehi _8811__254 (.L_HI(net254));
 sg13g2_tiehi _8986__255 (.L_HI(net255));
 sg13g2_tiehi _8823__256 (.L_HI(net256));
 sg13g2_tiehi _8980__257 (.L_HI(net257));
 sg13g2_tiehi _8822__258 (.L_HI(net258));
 sg13g2_tiehi _8985__259 (.L_HI(net259));
 sg13g2_tiehi _8821__260 (.L_HI(net260));
 sg13g2_tiehi _9007__261 (.L_HI(net261));
 sg13g2_tiehi _8820__262 (.L_HI(net262));
 sg13g2_tiehi _8984__263 (.L_HI(net263));
 sg13g2_tiehi _8819__264 (.L_HI(net264));
 sg13g2_tiehi _8860__265 (.L_HI(net265));
 sg13g2_tiehi _9015__266 (.L_HI(net266));
 sg13g2_tiehi _8818__267 (.L_HI(net267));
 sg13g2_tiehi _8983__268 (.L_HI(net268));
 sg13g2_tiehi _8817__269 (.L_HI(net269));
 sg13g2_tiehi _9006__270 (.L_HI(net270));
 sg13g2_tiehi _8816__271 (.L_HI(net271));
 sg13g2_tiehi _8982__272 (.L_HI(net272));
 sg13g2_tiehi _8815__273 (.L_HI(net273));
 sg13g2_tiehi _8981__274 (.L_HI(net274));
 sg13g2_tiehi _8814__275 (.L_HI(net275));
 sg13g2_tiehi _8916__276 (.L_HI(net276));
 sg13g2_tiehi _8813__277 (.L_HI(net277));
 sg13g2_tiehi _8812__278 (.L_HI(net278));
 sg13g2_tiehi _8915__279 (.L_HI(net279));
 sg13g2_tiehi _8809__280 (.L_HI(net280));
 sg13g2_tiehi _8808__281 (.L_HI(net281));
 sg13g2_tiehi _8807__282 (.L_HI(net282));
 sg13g2_tiehi _8806__283 (.L_HI(net283));
 sg13g2_tiehi _8805__284 (.L_HI(net284));
 sg13g2_tiehi _8804__285 (.L_HI(net285));
 sg13g2_tiehi _8803__286 (.L_HI(net286));
 sg13g2_tiehi _8802__287 (.L_HI(net287));
 sg13g2_tiehi _8801__288 (.L_HI(net288));
 sg13g2_tiehi _8800__289 (.L_HI(net289));
 sg13g2_tiehi _8799__290 (.L_HI(net290));
 sg13g2_tiehi _8798__291 (.L_HI(net291));
 sg13g2_tiehi _8797__292 (.L_HI(net292));
 sg13g2_tiehi _8796__293 (.L_HI(net293));
 sg13g2_tiehi _8795__294 (.L_HI(net294));
 sg13g2_tiehi _8871__295 (.L_HI(net295));
 sg13g2_tiehi _8901__296 (.L_HI(net296));
 sg13g2_tiehi _8902__297 (.L_HI(net297));
 sg13g2_tiehi _8794__298 (.L_HI(net298));
 sg13g2_tiehi _8793__299 (.L_HI(net299));
 sg13g2_tiehi _8792__300 (.L_HI(net300));
 sg13g2_tiehi _8791__301 (.L_HI(net301));
 sg13g2_tiehi _8790__302 (.L_HI(net302));
 sg13g2_tiehi _8789__303 (.L_HI(net303));
 sg13g2_tiehi _8914__304 (.L_HI(net304));
 sg13g2_tiehi _8788__305 (.L_HI(net305));
 sg13g2_tiehi _8787__306 (.L_HI(net306));
 sg13g2_tiehi _8786__307 (.L_HI(net307));
 sg13g2_tiehi _8785__308 (.L_HI(net308));
 sg13g2_tiehi _8784__309 (.L_HI(net309));
 sg13g2_tiehi _8783__310 (.L_HI(net310));
 sg13g2_tiehi _8903__311 (.L_HI(net311));
 sg13g2_tiehi _8917__312 (.L_HI(net312));
 sg13g2_tiehi _8918__313 (.L_HI(net313));
 sg13g2_tiehi _8919__314 (.L_HI(net314));
 sg13g2_tiehi _8920__315 (.L_HI(net315));
 sg13g2_tiehi _8921__316 (.L_HI(net316));
 sg13g2_tiehi _8922__317 (.L_HI(net317));
 sg13g2_tiehi _8923__318 (.L_HI(net318));
 sg13g2_tiehi _8924__319 (.L_HI(net319));
 sg13g2_tiehi _8925__320 (.L_HI(net320));
 sg13g2_tiehi _8926__321 (.L_HI(net321));
 sg13g2_tiehi _8927__322 (.L_HI(net322));
 sg13g2_tiehi _8928__323 (.L_HI(net323));
 sg13g2_tiehi _8929__324 (.L_HI(net324));
 sg13g2_tiehi _8930__325 (.L_HI(net325));
 sg13g2_tiehi _8931__326 (.L_HI(net326));
 sg13g2_tiehi _8932__327 (.L_HI(net327));
 sg13g2_tiehi _8933__328 (.L_HI(net328));
 sg13g2_tiehi _8934__329 (.L_HI(net329));
 sg13g2_tiehi _8935__330 (.L_HI(net330));
 sg13g2_tiehi _8936__331 (.L_HI(net331));
 sg13g2_tiehi _8937__332 (.L_HI(net332));
 sg13g2_tiehi _8938__333 (.L_HI(net333));
 sg13g2_tiehi _8939__334 (.L_HI(net334));
 sg13g2_tiehi _8940__335 (.L_HI(net335));
 sg13g2_tiehi _8941__336 (.L_HI(net336));
 sg13g2_tiehi _8942__337 (.L_HI(net337));
 sg13g2_tiehi _8943__338 (.L_HI(net338));
 sg13g2_tiehi _8944__339 (.L_HI(net339));
 sg13g2_tiehi _8945__340 (.L_HI(net340));
 sg13g2_tiehi _8946__341 (.L_HI(net341));
 sg13g2_tiehi _8947__342 (.L_HI(net342));
 sg13g2_tiehi _8948__343 (.L_HI(net343));
 sg13g2_tiehi _8949__344 (.L_HI(net344));
 sg13g2_tiehi _8950__345 (.L_HI(net345));
 sg13g2_tiehi _8951__346 (.L_HI(net346));
 sg13g2_tiehi _8952__347 (.L_HI(net347));
 sg13g2_tiehi _8953__348 (.L_HI(net348));
 sg13g2_tiehi _8954__349 (.L_HI(net349));
 sg13g2_tiehi _8955__350 (.L_HI(net350));
 sg13g2_tiehi _8956__351 (.L_HI(net351));
 sg13g2_tiehi _8957__352 (.L_HI(net352));
 sg13g2_tiehi _8958__353 (.L_HI(net353));
 sg13g2_tiehi _8959__354 (.L_HI(net354));
 sg13g2_tiehi _8960__355 (.L_HI(net355));
 sg13g2_tiehi _8961__356 (.L_HI(net356));
 sg13g2_tiehi _8962__357 (.L_HI(net357));
 sg13g2_tiehi _8963__358 (.L_HI(net358));
 sg13g2_tiehi _8964__359 (.L_HI(net359));
 sg13g2_tiehi _8965__360 (.L_HI(net360));
 sg13g2_tiehi _8966__361 (.L_HI(net361));
 sg13g2_tiehi _8967__362 (.L_HI(net362));
 sg13g2_tiehi _8968__363 (.L_HI(net363));
 sg13g2_tiehi _8969__364 (.L_HI(net364));
 sg13g2_tiehi _8970__365 (.L_HI(net365));
 sg13g2_tiehi _8971__366 (.L_HI(net366));
 sg13g2_tiehi _8972__367 (.L_HI(net367));
 sg13g2_tiehi _8973__368 (.L_HI(net368));
 sg13g2_tiehi _8974__369 (.L_HI(net369));
 sg13g2_tiehi _8975__370 (.L_HI(net370));
 sg13g2_tiehi _8976__371 (.L_HI(net371));
 sg13g2_tiehi _8977__372 (.L_HI(net372));
 sg13g2_tiehi _8978__373 (.L_HI(net373));
 sg13g2_tiehi _8979__374 (.L_HI(net374));
 sg13g2_tiehi _8782__375 (.L_HI(net375));
 sg13g2_tiehi _8781__376 (.L_HI(net376));
 sg13g2_tiehi _8780__377 (.L_HI(net377));
 sg13g2_tiehi _8779__378 (.L_HI(net378));
 sg13g2_tiehi _8778__379 (.L_HI(net379));
 sg13g2_tiehi _8777__380 (.L_HI(net380));
 sg13g2_tiehi _8776__381 (.L_HI(net381));
 sg13g2_tiehi _8775__382 (.L_HI(net382));
 sg13g2_tiehi _8774__383 (.L_HI(net383));
 sg13g2_tiehi _8773__384 (.L_HI(net384));
 sg13g2_tiehi _8772__385 (.L_HI(net385));
 sg13g2_tiehi _8771__386 (.L_HI(net386));
 sg13g2_tiehi _8770__387 (.L_HI(net387));
 sg13g2_tiehi _8769__388 (.L_HI(net388));
 sg13g2_tiehi _8768__389 (.L_HI(net389));
 sg13g2_tiehi _8913__390 (.L_HI(net390));
 sg13g2_tiehi _8767__391 (.L_HI(net391));
 sg13g2_tiehi _8766__392 (.L_HI(net392));
 sg13g2_tiehi _8765__393 (.L_HI(net393));
 sg13g2_tiehi _8764__394 (.L_HI(net394));
 sg13g2_tiehi _8763__395 (.L_HI(net395));
 sg13g2_tiehi _8762__396 (.L_HI(net396));
 sg13g2_tiehi _8761__397 (.L_HI(net397));
 sg13g2_tiehi _8760__398 (.L_HI(net398));
 sg13g2_tiehi _8759__399 (.L_HI(net399));
 sg13g2_tiehi _8758__400 (.L_HI(net400));
 sg13g2_tiehi _8757__401 (.L_HI(net401));
 sg13g2_tiehi _8756__402 (.L_HI(net402));
 sg13g2_tiehi _8755__403 (.L_HI(net403));
 sg13g2_tiehi _8754__404 (.L_HI(net404));
 sg13g2_tiehi _8753__405 (.L_HI(net405));
 sg13g2_tiehi _8752__406 (.L_HI(net406));
 sg13g2_tiehi _8751__407 (.L_HI(net407));
 sg13g2_tiehi _8750__408 (.L_HI(net408));
 sg13g2_tiehi _8749__409 (.L_HI(net409));
 sg13g2_tiehi _8748__410 (.L_HI(net410));
 sg13g2_tiehi _9019__411 (.L_HI(net411));
 sg13g2_tiehi _8747__412 (.L_HI(net412));
 sg13g2_tiehi _8746__413 (.L_HI(net413));
 sg13g2_tiehi _8745__414 (.L_HI(net414));
 sg13g2_tiehi _8744__415 (.L_HI(net415));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_2048_vga_game_18 (.L_LO(net18));
 sg13g2_tielo tt_um_2048_vga_game_19 (.L_LO(net19));
 sg13g2_tielo tt_um_2048_vga_game_20 (.L_LO(net20));
 sg13g2_tielo tt_um_2048_vga_game_21 (.L_LO(net21));
 sg13g2_tielo tt_um_2048_vga_game_22 (.L_LO(net22));
 sg13g2_tielo tt_um_2048_vga_game_23 (.L_LO(net23));
 sg13g2_tielo tt_um_2048_vga_game_24 (.L_LO(net24));
 sg13g2_tiehi _8743__25 (.L_HI(net25));
 sg13g2_buf_1 _9422_ (.A(\debug_controller_inst.data_out_en ),
    .X(uio_oe[4]));
 sg13g2_buf_1 _9423_ (.A(\debug_controller_inst.data_out_en ),
    .X(uio_oe[5]));
 sg13g2_buf_1 _9424_ (.A(\debug_controller_inst.data_out_en ),
    .X(uio_oe[6]));
 sg13g2_buf_1 _9425_ (.A(\debug_controller_inst.data_out_en ),
    .X(uio_oe[7]));
 sg13g2_buf_1 _9426_ (.A(\vga_sync_gen.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _9427_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_4 fanout1725 (.X(net1725),
    .A(_1286_));
 sg13g2_buf_4 fanout1726 (.X(net1726),
    .A(_1282_));
 sg13g2_buf_1 fanout1727 (.A(_1282_),
    .X(net1727));
 sg13g2_buf_4 fanout1728 (.X(net1728),
    .A(_0867_));
 sg13g2_buf_4 fanout1729 (.X(net1729),
    .A(_1790_));
 sg13g2_buf_4 fanout1730 (.X(net1730),
    .A(_1602_));
 sg13g2_buf_2 fanout1731 (.A(net1732),
    .X(net1731));
 sg13g2_buf_4 fanout1732 (.X(net1732),
    .A(_1466_));
 sg13g2_buf_4 fanout1733 (.X(net1733),
    .A(net1736));
 sg13g2_buf_4 fanout1734 (.X(net1734),
    .A(net1736));
 sg13g2_buf_1 fanout1735 (.A(net1736),
    .X(net1735));
 sg13g2_buf_4 fanout1736 (.X(net1736),
    .A(_0775_));
 sg13g2_buf_2 fanout1737 (.A(net1738),
    .X(net1737));
 sg13g2_buf_4 fanout1738 (.X(net1738),
    .A(net1741));
 sg13g2_buf_4 fanout1739 (.X(net1739),
    .A(net1741));
 sg13g2_buf_2 fanout1740 (.A(net1741),
    .X(net1740));
 sg13g2_buf_2 fanout1741 (.A(_0774_),
    .X(net1741));
 sg13g2_buf_4 fanout1742 (.X(net1742),
    .A(_1822_));
 sg13g2_buf_2 fanout1743 (.A(_1479_),
    .X(net1743));
 sg13g2_buf_2 fanout1744 (.A(net1745),
    .X(net1744));
 sg13g2_buf_2 fanout1745 (.A(net1746),
    .X(net1745));
 sg13g2_buf_2 fanout1746 (.A(net1749),
    .X(net1746));
 sg13g2_buf_4 fanout1747 (.X(net1747),
    .A(net1748));
 sg13g2_buf_4 fanout1748 (.X(net1748),
    .A(net1749));
 sg13g2_buf_2 fanout1749 (.A(_0870_),
    .X(net1749));
 sg13g2_buf_2 fanout1750 (.A(net1751),
    .X(net1750));
 sg13g2_buf_2 fanout1751 (.A(net1753),
    .X(net1751));
 sg13g2_buf_2 fanout1752 (.A(net1753),
    .X(net1752));
 sg13g2_buf_2 fanout1753 (.A(net1757),
    .X(net1753));
 sg13g2_buf_2 fanout1754 (.A(net1757),
    .X(net1754));
 sg13g2_buf_2 fanout1755 (.A(net1757),
    .X(net1755));
 sg13g2_buf_2 fanout1756 (.A(net1757),
    .X(net1756));
 sg13g2_buf_2 fanout1757 (.A(_0865_),
    .X(net1757));
 sg13g2_buf_2 fanout1758 (.A(net1761),
    .X(net1758));
 sg13g2_buf_2 fanout1759 (.A(net1760),
    .X(net1759));
 sg13g2_buf_2 fanout1760 (.A(net1761),
    .X(net1760));
 sg13g2_buf_2 fanout1761 (.A(_0706_),
    .X(net1761));
 sg13g2_buf_2 fanout1762 (.A(_0705_),
    .X(net1762));
 sg13g2_buf_2 fanout1763 (.A(_0705_),
    .X(net1763));
 sg13g2_buf_2 fanout1764 (.A(_0600_),
    .X(net1764));
 sg13g2_buf_2 fanout1765 (.A(_3595_),
    .X(net1765));
 sg13g2_buf_2 fanout1766 (.A(_3595_),
    .X(net1766));
 sg13g2_buf_2 fanout1767 (.A(net1769),
    .X(net1767));
 sg13g2_buf_2 fanout1768 (.A(net1769),
    .X(net1768));
 sg13g2_buf_1 fanout1769 (.A(_3554_),
    .X(net1769));
 sg13g2_buf_2 fanout1770 (.A(_3512_),
    .X(net1770));
 sg13g2_buf_2 fanout1771 (.A(_3512_),
    .X(net1771));
 sg13g2_buf_2 fanout1772 (.A(net1774),
    .X(net1772));
 sg13g2_buf_2 fanout1773 (.A(net1774),
    .X(net1773));
 sg13g2_buf_1 fanout1774 (.A(_3469_),
    .X(net1774));
 sg13g2_buf_4 fanout1775 (.X(net1775),
    .A(_0521_));
 sg13g2_buf_4 fanout1776 (.X(net1776),
    .A(_0520_));
 sg13g2_buf_1 fanout1777 (.A(_0520_),
    .X(net1777));
 sg13g2_buf_2 fanout1778 (.A(net1779),
    .X(net1778));
 sg13g2_buf_2 fanout1779 (.A(_3711_),
    .X(net1779));
 sg13g2_buf_2 fanout1780 (.A(net1781),
    .X(net1780));
 sg13g2_buf_1 fanout1781 (.A(net1782),
    .X(net1781));
 sg13g2_buf_1 fanout1782 (.A(_3711_),
    .X(net1782));
 sg13g2_buf_2 fanout1783 (.A(_0626_),
    .X(net1783));
 sg13g2_buf_4 fanout1784 (.X(net1784),
    .A(_3634_));
 sg13g2_buf_2 fanout1785 (.A(_3399_),
    .X(net1785));
 sg13g2_buf_2 fanout1786 (.A(_3399_),
    .X(net1786));
 sg13g2_buf_4 fanout1787 (.X(net1787),
    .A(_1900_));
 sg13g2_buf_4 fanout1788 (.X(net1788),
    .A(_1858_));
 sg13g2_buf_4 fanout1789 (.X(net1789),
    .A(_1702_));
 sg13g2_buf_4 fanout1790 (.X(net1790),
    .A(_1625_));
 sg13g2_buf_2 fanout1791 (.A(_0591_),
    .X(net1791));
 sg13g2_buf_4 fanout1792 (.X(net1792),
    .A(net1793));
 sg13g2_buf_4 fanout1793 (.X(net1793),
    .A(_3263_));
 sg13g2_buf_4 fanout1794 (.X(net1794),
    .A(_2024_));
 sg13g2_buf_2 fanout1795 (.A(_2001_),
    .X(net1795));
 sg13g2_buf_4 fanout1796 (.X(net1796),
    .A(_1750_));
 sg13g2_buf_4 fanout1797 (.X(net1797),
    .A(_1739_));
 sg13g2_buf_4 fanout1798 (.X(net1798),
    .A(_1642_));
 sg13g2_buf_4 fanout1799 (.X(net1799),
    .A(net1800));
 sg13g2_buf_4 fanout1800 (.X(net1800),
    .A(_1614_));
 sg13g2_buf_4 fanout1801 (.X(net1801),
    .A(_1553_));
 sg13g2_buf_4 fanout1802 (.X(net1802),
    .A(net1803));
 sg13g2_buf_2 fanout1803 (.A(_1539_),
    .X(net1803));
 sg13g2_buf_4 fanout1804 (.X(net1804),
    .A(_1511_));
 sg13g2_buf_2 fanout1805 (.A(_1511_),
    .X(net1805));
 sg13g2_buf_4 fanout1806 (.X(net1806),
    .A(_1510_));
 sg13g2_buf_4 fanout1807 (.X(net1807),
    .A(net1809));
 sg13g2_buf_1 fanout1808 (.A(net1809),
    .X(net1808));
 sg13g2_buf_4 fanout1809 (.X(net1809),
    .A(_1493_));
 sg13g2_buf_4 fanout1810 (.X(net1810),
    .A(net1812));
 sg13g2_buf_2 fanout1811 (.A(net1812),
    .X(net1811));
 sg13g2_buf_4 fanout1812 (.X(net1812),
    .A(_1492_));
 sg13g2_buf_4 fanout1813 (.X(net1813),
    .A(_1482_));
 sg13g2_buf_2 fanout1814 (.A(_1482_),
    .X(net1814));
 sg13g2_buf_2 fanout1815 (.A(net1816),
    .X(net1815));
 sg13g2_buf_2 fanout1816 (.A(_3872_),
    .X(net1816));
 sg13g2_buf_4 fanout1817 (.X(net1817),
    .A(_3779_));
 sg13g2_buf_4 fanout1818 (.X(net1818),
    .A(_3663_));
 sg13g2_buf_2 fanout1819 (.A(_3663_),
    .X(net1819));
 sg13g2_buf_4 fanout1820 (.X(net1820),
    .A(_3628_));
 sg13g2_buf_1 fanout1821 (.A(_3628_),
    .X(net1821));
 sg13g2_buf_2 fanout1822 (.A(net1823),
    .X(net1822));
 sg13g2_buf_2 fanout1823 (.A(_3262_),
    .X(net1823));
 sg13g2_buf_4 fanout1824 (.X(net1824),
    .A(net1828));
 sg13g2_buf_2 fanout1825 (.A(net1828),
    .X(net1825));
 sg13g2_buf_4 fanout1826 (.X(net1826),
    .A(net1827));
 sg13g2_buf_4 fanout1827 (.X(net1827),
    .A(net1828));
 sg13g2_buf_2 fanout1828 (.A(net1832),
    .X(net1828));
 sg13g2_buf_4 fanout1829 (.X(net1829),
    .A(net1831));
 sg13g2_buf_4 fanout1830 (.X(net1830),
    .A(net1831));
 sg13g2_buf_2 fanout1831 (.A(net1832),
    .X(net1831));
 sg13g2_buf_2 fanout1832 (.A(_3258_),
    .X(net1832));
 sg13g2_buf_4 fanout1833 (.X(net1833),
    .A(_1823_));
 sg13g2_buf_4 fanout1834 (.X(net1834),
    .A(net1836));
 sg13g2_buf_2 fanout1835 (.A(net1836),
    .X(net1835));
 sg13g2_buf_4 fanout1836 (.X(net1836),
    .A(_1814_));
 sg13g2_buf_4 fanout1837 (.X(net1837),
    .A(_1770_));
 sg13g2_buf_2 fanout1838 (.A(_1770_),
    .X(net1838));
 sg13g2_buf_4 fanout1839 (.X(net1839),
    .A(net1840));
 sg13g2_buf_4 fanout1840 (.X(net1840),
    .A(_1757_));
 sg13g2_buf_4 fanout1841 (.X(net1841),
    .A(_1749_));
 sg13g2_buf_4 fanout1842 (.X(net1842),
    .A(_1738_));
 sg13g2_buf_2 fanout1843 (.A(_1738_),
    .X(net1843));
 sg13g2_buf_4 fanout1844 (.X(net1844),
    .A(_1641_));
 sg13g2_buf_4 fanout1845 (.X(net1845),
    .A(net1846));
 sg13g2_buf_4 fanout1846 (.X(net1846),
    .A(_1640_));
 sg13g2_buf_4 fanout1847 (.X(net1847),
    .A(net1849));
 sg13g2_buf_2 fanout1848 (.A(net1849),
    .X(net1848));
 sg13g2_buf_4 fanout1849 (.X(net1849),
    .A(_1636_));
 sg13g2_buf_4 fanout1850 (.X(net1850),
    .A(_1616_));
 sg13g2_buf_8 fanout1851 (.A(_1608_),
    .X(net1851));
 sg13g2_buf_4 fanout1852 (.X(net1852),
    .A(_1608_));
 sg13g2_buf_2 fanout1853 (.A(net1854),
    .X(net1853));
 sg13g2_buf_4 fanout1854 (.X(net1854),
    .A(net1855));
 sg13g2_buf_4 fanout1855 (.X(net1855),
    .A(_1608_));
 sg13g2_buf_4 fanout1856 (.X(net1856),
    .A(net1857));
 sg13g2_buf_4 fanout1857 (.X(net1857),
    .A(_1591_));
 sg13g2_buf_4 fanout1858 (.X(net1858),
    .A(net1860));
 sg13g2_buf_4 fanout1859 (.X(net1859),
    .A(net1860));
 sg13g2_buf_8 fanout1860 (.A(_1590_),
    .X(net1860));
 sg13g2_buf_4 fanout1861 (.X(net1861),
    .A(net1862));
 sg13g2_buf_2 fanout1862 (.A(net1863),
    .X(net1862));
 sg13g2_buf_4 fanout1863 (.X(net1863),
    .A(_1552_));
 sg13g2_buf_4 fanout1864 (.X(net1864),
    .A(_1552_));
 sg13g2_buf_4 fanout1865 (.X(net1865),
    .A(net1866));
 sg13g2_buf_8 fanout1866 (.A(_1551_),
    .X(net1866));
 sg13g2_buf_4 fanout1867 (.X(net1867),
    .A(_1549_));
 sg13g2_buf_4 fanout1868 (.X(net1868),
    .A(_1534_));
 sg13g2_buf_4 fanout1869 (.X(net1869),
    .A(net1870));
 sg13g2_buf_4 fanout1870 (.X(net1870),
    .A(_1532_));
 sg13g2_buf_4 fanout1871 (.X(net1871),
    .A(net1873));
 sg13g2_buf_4 fanout1872 (.X(net1872),
    .A(net1873));
 sg13g2_buf_4 fanout1873 (.X(net1873),
    .A(_1531_));
 sg13g2_buf_4 fanout1874 (.X(net1874),
    .A(_1508_));
 sg13g2_buf_4 fanout1875 (.X(net1875),
    .A(_1508_));
 sg13g2_buf_4 fanout1876 (.X(net1876),
    .A(_1494_));
 sg13g2_buf_4 fanout1877 (.X(net1877),
    .A(_1490_));
 sg13g2_buf_4 fanout1878 (.X(net1878),
    .A(net1879));
 sg13g2_buf_8 fanout1879 (.A(_1489_),
    .X(net1879));
 sg13g2_buf_4 fanout1880 (.X(net1880),
    .A(_1488_));
 sg13g2_buf_2 fanout1881 (.A(_1488_),
    .X(net1881));
 sg13g2_buf_4 fanout1882 (.X(net1882),
    .A(_1487_));
 sg13g2_buf_4 fanout1883 (.X(net1883),
    .A(_1487_));
 sg13g2_buf_4 fanout1884 (.X(net1884),
    .A(_1485_));
 sg13g2_buf_4 fanout1885 (.X(net1885),
    .A(net1886));
 sg13g2_buf_4 fanout1886 (.X(net1886),
    .A(_1484_));
 sg13g2_buf_4 fanout1887 (.X(net1887),
    .A(_1483_));
 sg13g2_buf_4 fanout1888 (.X(net1888),
    .A(net1891));
 sg13g2_buf_4 fanout1889 (.X(net1889),
    .A(net1891));
 sg13g2_buf_2 fanout1890 (.A(net1891),
    .X(net1890));
 sg13g2_buf_4 fanout1891 (.X(net1891),
    .A(_1411_));
 sg13g2_buf_4 fanout1892 (.X(net1892),
    .A(_1400_));
 sg13g2_buf_4 fanout1893 (.X(net1893),
    .A(net1894));
 sg13g2_buf_4 fanout1894 (.X(net1894),
    .A(net1897));
 sg13g2_buf_4 fanout1895 (.X(net1895),
    .A(net1897));
 sg13g2_buf_2 fanout1896 (.A(net1897),
    .X(net1896));
 sg13g2_buf_2 fanout1897 (.A(_1396_),
    .X(net1897));
 sg13g2_buf_4 fanout1898 (.X(net1898),
    .A(net1899));
 sg13g2_buf_4 fanout1899 (.X(net1899),
    .A(_1395_));
 sg13g2_buf_4 fanout1900 (.X(net1900),
    .A(_1395_));
 sg13g2_buf_4 fanout1901 (.X(net1901),
    .A(_1395_));
 sg13g2_buf_4 fanout1902 (.X(net1902),
    .A(_1392_));
 sg13g2_buf_2 fanout1903 (.A(net1904),
    .X(net1903));
 sg13g2_buf_4 fanout1904 (.X(net1904),
    .A(_1392_));
 sg13g2_buf_4 fanout1905 (.X(net1905),
    .A(net1906));
 sg13g2_buf_4 fanout1906 (.X(net1906),
    .A(_1392_));
 sg13g2_buf_4 fanout1907 (.X(net1907),
    .A(_1391_));
 sg13g2_buf_4 fanout1908 (.X(net1908),
    .A(_1391_));
 sg13g2_buf_4 fanout1909 (.X(net1909),
    .A(net1911));
 sg13g2_buf_4 fanout1910 (.X(net1910),
    .A(net1911));
 sg13g2_buf_4 fanout1911 (.X(net1911),
    .A(_1391_));
 sg13g2_buf_4 fanout1912 (.X(net1912),
    .A(_1390_));
 sg13g2_buf_4 fanout1913 (.X(net1913),
    .A(_1390_));
 sg13g2_buf_2 fanout1914 (.A(net1915),
    .X(net1914));
 sg13g2_buf_4 fanout1915 (.X(net1915),
    .A(_1019_));
 sg13g2_buf_2 fanout1916 (.A(_0869_),
    .X(net1916));
 sg13g2_buf_4 fanout1917 (.X(net1917),
    .A(_0869_));
 sg13g2_buf_4 fanout1918 (.X(net1918),
    .A(_0638_));
 sg13g2_buf_2 fanout1919 (.A(_0546_),
    .X(net1919));
 sg13g2_buf_2 fanout1920 (.A(net1921),
    .X(net1920));
 sg13g2_buf_2 fanout1921 (.A(_3662_),
    .X(net1921));
 sg13g2_buf_2 fanout1922 (.A(_3627_),
    .X(net1922));
 sg13g2_buf_1 fanout1923 (.A(_3627_),
    .X(net1923));
 sg13g2_buf_4 fanout1924 (.X(net1924),
    .A(net1925));
 sg13g2_buf_2 fanout1925 (.A(net1926),
    .X(net1925));
 sg13g2_buf_2 fanout1926 (.A(_3255_),
    .X(net1926));
 sg13g2_buf_4 fanout1927 (.X(net1927),
    .A(net1928));
 sg13g2_buf_8 fanout1928 (.A(_1669_),
    .X(net1928));
 sg13g2_buf_4 fanout1929 (.X(net1929),
    .A(net1931));
 sg13g2_buf_4 fanout1930 (.X(net1930),
    .A(net1931));
 sg13g2_buf_2 fanout1931 (.A(_1617_),
    .X(net1931));
 sg13g2_buf_4 fanout1932 (.X(net1932),
    .A(net1933));
 sg13g2_buf_4 fanout1933 (.X(net1933),
    .A(_1609_));
 sg13g2_buf_4 fanout1934 (.X(net1934),
    .A(net1937));
 sg13g2_buf_4 fanout1935 (.X(net1935),
    .A(net1937));
 sg13g2_buf_1 fanout1936 (.A(net1937),
    .X(net1936));
 sg13g2_buf_2 fanout1937 (.A(_1609_),
    .X(net1937));
 sg13g2_buf_4 fanout1938 (.X(net1938),
    .A(net1941));
 sg13g2_buf_2 fanout1939 (.A(net1941),
    .X(net1939));
 sg13g2_buf_4 fanout1940 (.X(net1940),
    .A(net1941));
 sg13g2_buf_2 fanout1941 (.A(_1589_),
    .X(net1941));
 sg13g2_buf_4 fanout1942 (.X(net1942),
    .A(net1944));
 sg13g2_buf_2 fanout1943 (.A(net1944),
    .X(net1943));
 sg13g2_buf_4 fanout1944 (.X(net1944),
    .A(_1588_));
 sg13g2_buf_4 fanout1945 (.X(net1945),
    .A(_1573_));
 sg13g2_buf_2 fanout1946 (.A(_1573_),
    .X(net1946));
 sg13g2_buf_4 fanout1947 (.X(net1947),
    .A(_1569_));
 sg13g2_buf_4 fanout1948 (.X(net1948),
    .A(net1949));
 sg13g2_buf_4 fanout1949 (.X(net1949),
    .A(_1568_));
 sg13g2_buf_4 fanout1950 (.X(net1950),
    .A(_1535_));
 sg13g2_buf_4 fanout1951 (.X(net1951),
    .A(_1535_));
 sg13g2_buf_4 fanout1952 (.X(net1952),
    .A(net1953));
 sg13g2_buf_4 fanout1953 (.X(net1953),
    .A(net1954));
 sg13g2_buf_4 fanout1954 (.X(net1954),
    .A(_1529_));
 sg13g2_buf_4 fanout1955 (.X(net1955),
    .A(net1957));
 sg13g2_buf_1 fanout1956 (.A(net1957),
    .X(net1956));
 sg13g2_buf_4 fanout1957 (.X(net1957),
    .A(_1520_));
 sg13g2_buf_8 fanout1958 (.A(_1507_),
    .X(net1958));
 sg13g2_buf_4 fanout1959 (.X(net1959),
    .A(net1961));
 sg13g2_buf_4 fanout1960 (.X(net1960),
    .A(net1961));
 sg13g2_buf_4 fanout1961 (.X(net1961),
    .A(_1505_));
 sg13g2_buf_2 fanout1962 (.A(net1963),
    .X(net1962));
 sg13g2_buf_4 fanout1963 (.X(net1963),
    .A(net1964));
 sg13g2_buf_8 fanout1964 (.A(_1505_),
    .X(net1964));
 sg13g2_buf_8 fanout1965 (.A(net1970),
    .X(net1965));
 sg13g2_buf_2 fanout1966 (.A(net1970),
    .X(net1966));
 sg13g2_buf_4 fanout1967 (.X(net1967),
    .A(net1970));
 sg13g2_buf_2 fanout1968 (.A(net1969),
    .X(net1968));
 sg13g2_buf_4 fanout1969 (.X(net1969),
    .A(net1970));
 sg13g2_buf_2 fanout1970 (.A(_1504_),
    .X(net1970));
 sg13g2_buf_4 fanout1971 (.X(net1971),
    .A(_1498_));
 sg13g2_buf_1 fanout1972 (.A(_1498_),
    .X(net1972));
 sg13g2_buf_4 fanout1973 (.X(net1973),
    .A(_1497_));
 sg13g2_buf_4 fanout1974 (.X(net1974),
    .A(_1495_));
 sg13g2_buf_2 fanout1975 (.A(_1495_),
    .X(net1975));
 sg13g2_buf_4 fanout1976 (.X(net1976),
    .A(_1486_));
 sg13g2_buf_2 fanout1977 (.A(_1486_),
    .X(net1977));
 sg13g2_buf_4 fanout1978 (.X(net1978),
    .A(_1426_));
 sg13g2_buf_2 fanout1979 (.A(net1980),
    .X(net1979));
 sg13g2_buf_4 fanout1980 (.X(net1980),
    .A(_1419_));
 sg13g2_buf_4 fanout1981 (.X(net1981),
    .A(net1982));
 sg13g2_buf_2 fanout1982 (.A(net1984),
    .X(net1982));
 sg13g2_buf_4 fanout1983 (.X(net1983),
    .A(net1984));
 sg13g2_buf_4 fanout1984 (.X(net1984),
    .A(_1413_));
 sg13g2_buf_4 fanout1985 (.X(net1985),
    .A(net1986));
 sg13g2_buf_2 fanout1986 (.A(net1990),
    .X(net1986));
 sg13g2_buf_4 fanout1987 (.X(net1987),
    .A(net1990));
 sg13g2_buf_4 fanout1988 (.X(net1988),
    .A(net1990));
 sg13g2_buf_2 fanout1989 (.A(net1990),
    .X(net1989));
 sg13g2_buf_2 fanout1990 (.A(_1412_),
    .X(net1990));
 sg13g2_buf_4 fanout1991 (.X(net1991),
    .A(net1995));
 sg13g2_buf_2 fanout1992 (.A(net1995),
    .X(net1992));
 sg13g2_buf_4 fanout1993 (.X(net1993),
    .A(net1994));
 sg13g2_buf_4 fanout1994 (.X(net1994),
    .A(net1995));
 sg13g2_buf_4 fanout1995 (.X(net1995),
    .A(_1410_));
 sg13g2_buf_4 fanout1996 (.X(net1996),
    .A(_1399_));
 sg13g2_buf_2 fanout1997 (.A(net1998),
    .X(net1997));
 sg13g2_buf_4 fanout1998 (.X(net1998),
    .A(net1999));
 sg13g2_buf_2 fanout1999 (.A(_0543_),
    .X(net1999));
 sg13g2_buf_2 fanout2000 (.A(net2001),
    .X(net2000));
 sg13g2_buf_2 fanout2001 (.A(_0542_),
    .X(net2001));
 sg13g2_buf_2 fanout2002 (.A(net2004),
    .X(net2002));
 sg13g2_buf_1 fanout2003 (.A(net2004),
    .X(net2003));
 sg13g2_buf_4 fanout2004 (.X(net2004),
    .A(_0541_));
 sg13g2_buf_4 fanout2005 (.X(net2005),
    .A(_0540_));
 sg13g2_buf_4 fanout2006 (.X(net2006),
    .A(net2008));
 sg13g2_buf_2 fanout2007 (.A(net2008),
    .X(net2007));
 sg13g2_buf_2 fanout2008 (.A(_0539_),
    .X(net2008));
 sg13g2_buf_4 fanout2009 (.X(net2009),
    .A(net2010));
 sg13g2_buf_2 fanout2010 (.A(net2011),
    .X(net2010));
 sg13g2_buf_4 fanout2011 (.X(net2011),
    .A(_0538_));
 sg13g2_buf_2 fanout2012 (.A(net2013),
    .X(net2012));
 sg13g2_buf_2 fanout2013 (.A(net2014),
    .X(net2013));
 sg13g2_buf_2 fanout2014 (.A(net2015),
    .X(net2014));
 sg13g2_buf_2 fanout2015 (.A(_0537_),
    .X(net2015));
 sg13g2_buf_2 fanout2016 (.A(net2017),
    .X(net2016));
 sg13g2_buf_2 fanout2017 (.A(net2019),
    .X(net2017));
 sg13g2_buf_2 fanout2018 (.A(net2019),
    .X(net2018));
 sg13g2_buf_2 fanout2019 (.A(_0536_),
    .X(net2019));
 sg13g2_buf_4 fanout2020 (.X(net2020),
    .A(_0535_));
 sg13g2_buf_4 fanout2021 (.X(net2021),
    .A(net2022));
 sg13g2_buf_2 fanout2022 (.A(net2023),
    .X(net2022));
 sg13g2_buf_8 fanout2023 (.A(_4002_),
    .X(net2023));
 sg13g2_buf_4 fanout2024 (.X(net2024),
    .A(net2026));
 sg13g2_buf_1 fanout2025 (.A(net2026),
    .X(net2025));
 sg13g2_buf_4 fanout2026 (.X(net2026),
    .A(_4001_));
 sg13g2_buf_4 fanout2027 (.X(net2027),
    .A(net2028));
 sg13g2_buf_4 fanout2028 (.X(net2028),
    .A(_3999_));
 sg13g2_buf_4 fanout2029 (.X(net2029),
    .A(net2031));
 sg13g2_buf_2 fanout2030 (.A(net2031),
    .X(net2030));
 sg13g2_buf_4 fanout2031 (.X(net2031),
    .A(net2032));
 sg13g2_buf_4 fanout2032 (.X(net2032),
    .A(_3998_));
 sg13g2_buf_4 fanout2033 (.X(net2033),
    .A(net2034));
 sg13g2_buf_4 fanout2034 (.X(net2034),
    .A(net2037));
 sg13g2_buf_4 fanout2035 (.X(net2035),
    .A(net2037));
 sg13g2_buf_4 fanout2036 (.X(net2036),
    .A(net2037));
 sg13g2_buf_4 fanout2037 (.X(net2037),
    .A(_3998_));
 sg13g2_buf_4 fanout2038 (.X(net2038),
    .A(net2041));
 sg13g2_buf_4 fanout2039 (.X(net2039),
    .A(net2041));
 sg13g2_buf_1 fanout2040 (.A(net2041),
    .X(net2040));
 sg13g2_buf_4 fanout2041 (.X(net2041),
    .A(_3997_));
 sg13g2_buf_4 fanout2042 (.X(net2042),
    .A(net2044));
 sg13g2_buf_4 fanout2043 (.X(net2043),
    .A(_3997_));
 sg13g2_buf_2 fanout2044 (.A(_3997_),
    .X(net2044));
 sg13g2_buf_4 fanout2045 (.X(net2045),
    .A(net2047));
 sg13g2_buf_2 fanout2046 (.A(net2047),
    .X(net2046));
 sg13g2_buf_4 fanout2047 (.X(net2047),
    .A(_3996_));
 sg13g2_buf_4 fanout2048 (.X(net2048),
    .A(net2050));
 sg13g2_buf_4 fanout2049 (.X(net2049),
    .A(net2050));
 sg13g2_buf_4 fanout2050 (.X(net2050),
    .A(_3996_));
 sg13g2_buf_4 fanout2051 (.X(net2051),
    .A(_3994_));
 sg13g2_buf_2 fanout2052 (.A(_3994_),
    .X(net2052));
 sg13g2_buf_2 fanout2053 (.A(net2054),
    .X(net2053));
 sg13g2_buf_4 fanout2054 (.X(net2054),
    .A(net2060));
 sg13g2_buf_2 fanout2055 (.A(net2056),
    .X(net2055));
 sg13g2_buf_2 fanout2056 (.A(net2060),
    .X(net2056));
 sg13g2_buf_2 fanout2057 (.A(net2059),
    .X(net2057));
 sg13g2_buf_2 fanout2058 (.A(net2059),
    .X(net2058));
 sg13g2_buf_2 fanout2059 (.A(net2060),
    .X(net2059));
 sg13g2_buf_2 fanout2060 (.A(_3977_),
    .X(net2060));
 sg13g2_buf_2 fanout2061 (.A(net2064),
    .X(net2061));
 sg13g2_buf_2 fanout2062 (.A(net2064),
    .X(net2062));
 sg13g2_buf_1 fanout2063 (.A(net2064),
    .X(net2063));
 sg13g2_buf_1 fanout2064 (.A(_3960_),
    .X(net2064));
 sg13g2_buf_2 fanout2065 (.A(net2068),
    .X(net2065));
 sg13g2_buf_2 fanout2066 (.A(net2068),
    .X(net2066));
 sg13g2_buf_2 fanout2067 (.A(net2068),
    .X(net2067));
 sg13g2_buf_2 fanout2068 (.A(_3960_),
    .X(net2068));
 sg13g2_buf_4 fanout2069 (.X(net2069),
    .A(_3932_));
 sg13g2_buf_4 fanout2070 (.X(net2070),
    .A(_3931_));
 sg13g2_buf_2 fanout2071 (.A(net2073),
    .X(net2071));
 sg13g2_buf_1 fanout2072 (.A(net2073),
    .X(net2072));
 sg13g2_buf_2 fanout2073 (.A(net2074),
    .X(net2073));
 sg13g2_buf_2 fanout2074 (.A(net951),
    .X(net2074));
 sg13g2_buf_2 fanout2075 (.A(net2076),
    .X(net2075));
 sg13g2_buf_2 fanout2076 (.A(net2077),
    .X(net2076));
 sg13g2_buf_2 fanout2077 (.A(net1031),
    .X(net2077));
 sg13g2_buf_2 fanout2078 (.A(net2080),
    .X(net2078));
 sg13g2_buf_1 fanout2079 (.A(net2080),
    .X(net2079));
 sg13g2_buf_2 fanout2080 (.A(net2081),
    .X(net2080));
 sg13g2_buf_4 fanout2081 (.X(net2081),
    .A(net2083));
 sg13g2_buf_4 fanout2082 (.X(net2082),
    .A(net2083));
 sg13g2_buf_4 fanout2083 (.X(net2083),
    .A(net982));
 sg13g2_buf_4 fanout2084 (.X(net2084),
    .A(\debug_controller_inst.grid_out_addr[2] ));
 sg13g2_buf_2 fanout2085 (.A(\debug_controller_inst.grid_out_addr[2] ),
    .X(net2085));
 sg13g2_buf_4 fanout2086 (.X(net2086),
    .A(net2087));
 sg13g2_buf_4 fanout2087 (.X(net2087),
    .A(net1032));
 sg13g2_buf_4 fanout2088 (.X(net2088),
    .A(net2089));
 sg13g2_buf_4 fanout2089 (.X(net2089),
    .A(net983));
 sg13g2_buf_4 fanout2090 (.X(net2090),
    .A(net2091));
 sg13g2_buf_4 fanout2091 (.X(net2091),
    .A(net940));
 sg13g2_buf_4 fanout2092 (.X(net2092),
    .A(net2093));
 sg13g2_buf_4 fanout2093 (.X(net2093),
    .A(net991));
 sg13g2_buf_4 fanout2094 (.X(net2094),
    .A(\game_logic_inst.current_row_index[1] ));
 sg13g2_buf_4 fanout2095 (.X(net2095),
    .A(net2096));
 sg13g2_buf_4 fanout2096 (.X(net2096),
    .A(\game_logic_inst.current_row_index[1] ));
 sg13g2_buf_8 fanout2097 (.A(\game_logic_inst.current_row_index[0] ),
    .X(net2097));
 sg13g2_buf_8 fanout2098 (.A(net2099),
    .X(net2098));
 sg13g2_buf_4 fanout2099 (.X(net2099),
    .A(\game_logic_inst.current_row_index[0] ));
 sg13g2_buf_2 fanout2100 (.A(\game_logic_inst.added_tile_index[3] ),
    .X(net2100));
 sg13g2_buf_2 fanout2101 (.A(net2102),
    .X(net2101));
 sg13g2_buf_2 fanout2102 (.A(\game_logic_inst.added_tile_index[2] ),
    .X(net2102));
 sg13g2_buf_4 fanout2103 (.X(net2103),
    .A(net915));
 sg13g2_buf_2 fanout2104 (.A(net2110),
    .X(net2104));
 sg13g2_buf_2 fanout2105 (.A(net2106),
    .X(net2105));
 sg13g2_buf_4 fanout2106 (.X(net2106),
    .A(net2110));
 sg13g2_buf_2 fanout2107 (.A(net2108),
    .X(net2107));
 sg13g2_buf_2 fanout2108 (.A(net2110),
    .X(net2108));
 sg13g2_buf_1 fanout2109 (.A(net2110),
    .X(net2109));
 sg13g2_buf_2 fanout2110 (.A(\game_logic_inst.game_started ),
    .X(net2110));
 sg13g2_buf_2 fanout2111 (.A(net2112),
    .X(net2111));
 sg13g2_buf_2 fanout2112 (.A(net2113),
    .X(net2112));
 sg13g2_buf_2 fanout2113 (.A(\game_logic_inst.game_started ),
    .X(net2113));
 sg13g2_buf_2 fanout2114 (.A(net2117),
    .X(net2114));
 sg13g2_buf_2 fanout2115 (.A(net2116),
    .X(net2115));
 sg13g2_buf_2 fanout2116 (.A(net2117),
    .X(net2116));
 sg13g2_buf_2 fanout2117 (.A(\game_logic_inst.game_started ),
    .X(net2117));
 sg13g2_buf_2 fanout2118 (.A(net2119),
    .X(net2118));
 sg13g2_buf_2 fanout2119 (.A(net2120),
    .X(net2119));
 sg13g2_buf_2 fanout2120 (.A(net2121),
    .X(net2120));
 sg13g2_buf_4 fanout2121 (.X(net2121),
    .A(\game_logic_inst.calculate_move ));
 sg13g2_buf_2 fanout2122 (.A(net1007),
    .X(net2122));
 sg13g2_buf_4 fanout2123 (.X(net2123),
    .A(net2125));
 sg13g2_buf_4 fanout2124 (.X(net2124),
    .A(\draw_game_inst.x[7] ));
 sg13g2_buf_2 fanout2125 (.A(\draw_game_inst.x[7] ),
    .X(net2125));
 sg13g2_buf_8 fanout2126 (.A(net2127),
    .X(net2126));
 sg13g2_buf_4 fanout2127 (.X(net2127),
    .A(\draw_game_inst.x[6] ));
 sg13g2_buf_4 fanout2128 (.X(net2128),
    .A(net1015));
 sg13g2_buf_4 fanout2129 (.X(net2129),
    .A(net1015));
 sg13g2_buf_2 fanout2130 (.A(net2131),
    .X(net2130));
 sg13g2_buf_2 fanout2131 (.A(net2133),
    .X(net2131));
 sg13g2_buf_4 fanout2132 (.X(net2132),
    .A(net2133));
 sg13g2_buf_2 fanout2133 (.A(_0094_),
    .X(net2133));
 sg13g2_buf_4 fanout2134 (.X(net2134),
    .A(net2135));
 sg13g2_buf_4 fanout2135 (.X(net2135),
    .A(net2139));
 sg13g2_buf_4 fanout2136 (.X(net2136),
    .A(net2137));
 sg13g2_buf_4 fanout2137 (.X(net2137),
    .A(net2138));
 sg13g2_buf_4 fanout2138 (.X(net2138),
    .A(net2139));
 sg13g2_buf_2 fanout2139 (.A(\draw_game_inst.board_x[5] ),
    .X(net2139));
 sg13g2_buf_4 fanout2140 (.X(net2140),
    .A(net2141));
 sg13g2_buf_4 fanout2141 (.X(net2141),
    .A(net2142));
 sg13g2_buf_4 fanout2142 (.X(net2142),
    .A(net2143));
 sg13g2_buf_4 fanout2143 (.X(net2143),
    .A(\draw_game_inst.board_x[4] ));
 sg13g2_buf_4 fanout2144 (.X(net2144),
    .A(\draw_game_inst.board_x[4] ));
 sg13g2_buf_4 fanout2145 (.X(net2145),
    .A(_0095_));
 sg13g2_buf_4 fanout2146 (.X(net2146),
    .A(_0095_));
 sg13g2_buf_4 fanout2147 (.X(net2147),
    .A(net2148));
 sg13g2_buf_2 fanout2148 (.A(net2151),
    .X(net2148));
 sg13g2_buf_4 fanout2149 (.X(net2149),
    .A(net2150));
 sg13g2_buf_2 fanout2150 (.A(net2151),
    .X(net2150));
 sg13g2_buf_4 fanout2151 (.X(net2151),
    .A(\draw_game_inst.board_x[3] ));
 sg13g2_buf_2 fanout2152 (.A(net2153),
    .X(net2152));
 sg13g2_buf_4 fanout2153 (.X(net2153),
    .A(\draw_game_inst.y[7] ));
 sg13g2_buf_4 fanout2154 (.X(net2154),
    .A(\draw_game_inst.board_y[6] ));
 sg13g2_buf_2 fanout2155 (.A(net2157),
    .X(net2155));
 sg13g2_buf_2 fanout2156 (.A(net2157),
    .X(net2156));
 sg13g2_buf_4 fanout2157 (.X(net2157),
    .A(\draw_game_inst.board_y[5] ));
 sg13g2_buf_4 fanout2158 (.X(net2158),
    .A(net2159));
 sg13g2_buf_4 fanout2159 (.X(net2159),
    .A(\draw_game_inst.board_y[5] ));
 sg13g2_buf_4 fanout2160 (.X(net2160),
    .A(net2161));
 sg13g2_buf_4 fanout2161 (.X(net2161),
    .A(_0090_));
 sg13g2_buf_4 fanout2162 (.X(net2162),
    .A(net2165));
 sg13g2_buf_2 fanout2163 (.A(net2164),
    .X(net2163));
 sg13g2_buf_4 fanout2164 (.X(net2164),
    .A(net2165));
 sg13g2_buf_2 fanout2165 (.A(\draw_game_inst.board_y[4] ),
    .X(net2165));
 sg13g2_buf_4 fanout2166 (.X(net2166),
    .A(net2167));
 sg13g2_buf_4 fanout2167 (.X(net2167),
    .A(net2182));
 sg13g2_buf_2 fanout2168 (.A(net2169),
    .X(net2168));
 sg13g2_buf_1 fanout2169 (.A(net2170),
    .X(net2169));
 sg13g2_buf_2 fanout2170 (.A(net2182),
    .X(net2170));
 sg13g2_buf_2 fanout2171 (.A(net2173),
    .X(net2171));
 sg13g2_buf_2 fanout2172 (.A(net2173),
    .X(net2172));
 sg13g2_buf_2 fanout2173 (.A(net2182),
    .X(net2173));
 sg13g2_buf_2 fanout2174 (.A(net2178),
    .X(net2174));
 sg13g2_buf_2 fanout2175 (.A(net2177),
    .X(net2175));
 sg13g2_buf_2 fanout2176 (.A(net2177),
    .X(net2176));
 sg13g2_buf_2 fanout2177 (.A(net2178),
    .X(net2177));
 sg13g2_buf_2 fanout2178 (.A(net2182),
    .X(net2178));
 sg13g2_buf_2 fanout2179 (.A(net2180),
    .X(net2179));
 sg13g2_buf_4 fanout2180 (.X(net2180),
    .A(net2181));
 sg13g2_buf_4 fanout2181 (.X(net2181),
    .A(net2182));
 sg13g2_buf_4 fanout2182 (.X(net2182),
    .A(\draw_game_inst.board_y[3] ));
 sg13g2_buf_4 fanout2183 (.X(net2183),
    .A(net2185));
 sg13g2_buf_4 fanout2184 (.X(net2184),
    .A(net2185));
 sg13g2_buf_4 fanout2185 (.X(net2185),
    .A(_0092_));
 sg13g2_buf_2 fanout2186 (.A(net2187),
    .X(net2186));
 sg13g2_buf_4 fanout2187 (.X(net2187),
    .A(net2190));
 sg13g2_buf_4 fanout2188 (.X(net2188),
    .A(net2189));
 sg13g2_buf_4 fanout2189 (.X(net2189),
    .A(net2190));
 sg13g2_buf_2 fanout2190 (.A(net1025),
    .X(net2190));
 sg13g2_buf_4 fanout2191 (.X(net2191),
    .A(net2194));
 sg13g2_buf_2 fanout2192 (.A(net2194),
    .X(net2192));
 sg13g2_buf_4 fanout2193 (.X(net2193),
    .A(net2194));
 sg13g2_buf_4 fanout2194 (.X(net2194),
    .A(\draw_game_inst.board_y[2] ));
 sg13g2_buf_2 fanout2195 (.A(net2197),
    .X(net2195));
 sg13g2_buf_2 fanout2196 (.A(net2197),
    .X(net2196));
 sg13g2_buf_4 fanout2197 (.X(net2197),
    .A(\draw_game_inst.board_y[2] ));
 sg13g2_buf_2 fanout2198 (.A(_0093_),
    .X(net2198));
 sg13g2_buf_2 fanout2199 (.A(net2200),
    .X(net2199));
 sg13g2_buf_2 fanout2200 (.A(net2202),
    .X(net2200));
 sg13g2_buf_4 fanout2201 (.X(net2201),
    .A(net2202));
 sg13g2_buf_2 fanout2202 (.A(net2224),
    .X(net2202));
 sg13g2_buf_2 fanout2203 (.A(net2206),
    .X(net2203));
 sg13g2_buf_2 fanout2204 (.A(net2205),
    .X(net2204));
 sg13g2_buf_2 fanout2205 (.A(net2206),
    .X(net2205));
 sg13g2_buf_2 fanout2206 (.A(net2224),
    .X(net2206));
 sg13g2_buf_2 fanout2207 (.A(net2209),
    .X(net2207));
 sg13g2_buf_2 fanout2208 (.A(net2209),
    .X(net2208));
 sg13g2_buf_2 fanout2209 (.A(net2224),
    .X(net2209));
 sg13g2_buf_2 fanout2210 (.A(net2211),
    .X(net2210));
 sg13g2_buf_4 fanout2211 (.X(net2211),
    .A(net2223));
 sg13g2_buf_2 fanout2212 (.A(net2213),
    .X(net2212));
 sg13g2_buf_2 fanout2213 (.A(net2223),
    .X(net2213));
 sg13g2_buf_2 fanout2214 (.A(net2217),
    .X(net2214));
 sg13g2_buf_2 fanout2215 (.A(net2217),
    .X(net2215));
 sg13g2_buf_4 fanout2216 (.X(net2216),
    .A(net2217));
 sg13g2_buf_2 fanout2217 (.A(net2222),
    .X(net2217));
 sg13g2_buf_4 fanout2218 (.X(net2218),
    .A(net2222));
 sg13g2_buf_4 fanout2219 (.X(net2219),
    .A(net2222));
 sg13g2_buf_4 fanout2220 (.X(net2220),
    .A(net2221));
 sg13g2_buf_4 fanout2221 (.X(net2221),
    .A(net2222));
 sg13g2_buf_2 fanout2222 (.A(net2223),
    .X(net2222));
 sg13g2_buf_2 fanout2223 (.A(net2224),
    .X(net2223));
 sg13g2_buf_4 fanout2224 (.X(net2224),
    .A(\draw_game_inst.board_y[1] ));
 sg13g2_buf_4 fanout2225 (.X(net2225),
    .A(net962));
 sg13g2_buf_4 fanout2226 (.X(net2226),
    .A(_0171_));
 sg13g2_buf_2 fanout2227 (.A(net2228),
    .X(net2227));
 sg13g2_buf_2 fanout2228 (.A(net2229),
    .X(net2228));
 sg13g2_buf_2 fanout2229 (.A(net2237),
    .X(net2229));
 sg13g2_buf_2 fanout2230 (.A(net2233),
    .X(net2230));
 sg13g2_buf_2 fanout2231 (.A(net2232),
    .X(net2231));
 sg13g2_buf_2 fanout2232 (.A(net2233),
    .X(net2232));
 sg13g2_buf_1 fanout2233 (.A(net2237),
    .X(net2233));
 sg13g2_buf_2 fanout2234 (.A(net2235),
    .X(net2234));
 sg13g2_buf_2 fanout2235 (.A(net2237),
    .X(net2235));
 sg13g2_buf_4 fanout2236 (.X(net2236),
    .A(net2237));
 sg13g2_buf_4 fanout2237 (.X(net2237),
    .A(\draw_game_inst.board_y[0] ));
 sg13g2_buf_4 fanout2238 (.X(net2238),
    .A(net2240));
 sg13g2_buf_4 fanout2239 (.X(net2239),
    .A(net2240));
 sg13g2_buf_4 fanout2240 (.X(net2240),
    .A(\draw_game_inst.board_y[0] ));
 sg13g2_buf_2 fanout2241 (.A(net2249),
    .X(net2241));
 sg13g2_buf_1 fanout2242 (.A(net2249),
    .X(net2242));
 sg13g2_buf_2 fanout2243 (.A(net2249),
    .X(net2243));
 sg13g2_buf_4 fanout2244 (.X(net2244),
    .A(net2249));
 sg13g2_buf_2 fanout2245 (.A(net2249),
    .X(net2245));
 sg13g2_buf_4 fanout2246 (.X(net2246),
    .A(net2247));
 sg13g2_buf_2 fanout2247 (.A(net2248),
    .X(net2247));
 sg13g2_buf_4 fanout2248 (.X(net2248),
    .A(net2249));
 sg13g2_buf_4 fanout2249 (.X(net2249),
    .A(\draw_game_inst.board_y[0] ));
 sg13g2_buf_2 fanout2250 (.A(_0167_),
    .X(net2250));
 sg13g2_buf_2 fanout2251 (.A(_0167_),
    .X(net2251));
 sg13g2_buf_2 fanout2252 (.A(net1010),
    .X(net2252));
 sg13g2_buf_2 fanout2253 (.A(net1009),
    .X(net2253));
 sg13g2_buf_4 fanout2254 (.X(net2254),
    .A(net2256));
 sg13g2_buf_4 fanout2255 (.X(net2255),
    .A(net2256));
 sg13g2_buf_2 fanout2256 (.A(show_welcome_screen),
    .X(net2256));
 sg13g2_buf_4 fanout2257 (.X(net2257),
    .A(net2258));
 sg13g2_buf_4 fanout2258 (.X(net2258),
    .A(net2259));
 sg13g2_buf_4 fanout2259 (.X(net2259),
    .A(_3978_));
 sg13g2_buf_4 fanout2260 (.X(net2260),
    .A(net2263));
 sg13g2_buf_2 fanout2261 (.A(net2263),
    .X(net2261));
 sg13g2_buf_2 fanout2262 (.A(net2263),
    .X(net2262));
 sg13g2_buf_2 fanout2263 (.A(_3978_),
    .X(net2263));
 sg13g2_buf_2 fanout2264 (.A(net2266),
    .X(net2264));
 sg13g2_buf_1 fanout2265 (.A(net2266),
    .X(net2265));
 sg13g2_buf_1 fanout2266 (.A(net2269),
    .X(net2266));
 sg13g2_buf_2 fanout2267 (.A(net2268),
    .X(net2267));
 sg13g2_buf_2 fanout2268 (.A(net2269),
    .X(net2268));
 sg13g2_buf_2 fanout2269 (.A(net2279),
    .X(net2269));
 sg13g2_buf_2 fanout2270 (.A(net2274),
    .X(net2270));
 sg13g2_buf_1 fanout2271 (.A(net2274),
    .X(net2271));
 sg13g2_buf_2 fanout2272 (.A(net2273),
    .X(net2272));
 sg13g2_buf_2 fanout2273 (.A(net2274),
    .X(net2273));
 sg13g2_buf_2 fanout2274 (.A(net2279),
    .X(net2274));
 sg13g2_buf_4 fanout2275 (.X(net2275),
    .A(net2279));
 sg13g2_buf_2 fanout2276 (.A(net2279),
    .X(net2276));
 sg13g2_buf_4 fanout2277 (.X(net2277),
    .A(net2278));
 sg13g2_buf_4 fanout2278 (.X(net2278),
    .A(net2279));
 sg13g2_buf_4 fanout2279 (.X(net2279),
    .A(rst_n));
 sg13g2_buf_2 fanout2280 (.A(net2284),
    .X(net2280));
 sg13g2_buf_2 fanout2281 (.A(net2284),
    .X(net2281));
 sg13g2_buf_2 fanout2282 (.A(net2284),
    .X(net2282));
 sg13g2_buf_2 fanout2283 (.A(net2284),
    .X(net2283));
 sg13g2_buf_1 fanout2284 (.A(net2285),
    .X(net2284));
 sg13g2_buf_2 fanout2285 (.A(net2292),
    .X(net2285));
 sg13g2_buf_4 fanout2286 (.X(net2286),
    .A(net2292));
 sg13g2_buf_2 fanout2287 (.A(net2292),
    .X(net2287));
 sg13g2_buf_4 fanout2288 (.X(net2288),
    .A(net2291));
 sg13g2_buf_4 fanout2289 (.X(net2289),
    .A(net2291));
 sg13g2_buf_4 fanout2290 (.X(net2290),
    .A(net2291));
 sg13g2_buf_4 fanout2291 (.X(net2291),
    .A(net2292));
 sg13g2_buf_2 fanout2292 (.A(rst_n),
    .X(net2292));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_4 input5 (.X(net5),
    .A(ui_in[4]));
 sg13g2_buf_4 input6 (.X(net6),
    .A(ui_in[5]));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_2 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[3]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[4]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[5]),
    .X(net14));
 sg13g2_buf_2 input15 (.A(uio_in[6]),
    .X(net15));
 sg13g2_buf_1 input16 (.A(uio_in[7]),
    .X(net16));
 sg13g2_tielo tt_um_2048_vga_game_17 (.L_LO(net17));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_leaf_49_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_2 clkbuf_leaf_50_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_2 clkbuf_leaf_51_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_2 clkbuf_leaf_52_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_2 clkbuf_leaf_53_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_2 clkbuf_leaf_54_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_2 clkbuf_leaf_55_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_2 clkbuf_leaf_56_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_2 clkbuf_leaf_57_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_2 clkbuf_leaf_58_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_2 clkbuf_leaf_59_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_2 clkbuf_leaf_60_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_4_2_0_clk));
 sg13g2_buf_1 clkload2 (.A(clknet_4_3_0_clk));
 sg13g2_buf_1 clkload3 (.A(clknet_4_4_0_clk));
 sg13g2_buf_1 clkload4 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_7_0_clk));
 sg13g2_buf_1 clkload6 (.A(clknet_4_8_0_clk));
 sg13g2_buf_1 clkload7 (.A(clknet_4_10_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_11_0_clk));
 sg13g2_buf_1 clkload9 (.A(clknet_4_12_0_clk));
 sg13g2_buf_1 clkload10 (.A(clknet_4_13_0_clk));
 sg13g2_buf_1 clkload11 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_4_15_0_clk));
 sg13g2_inv_4 clkload13 (.A(clknet_leaf_60_clk));
 sg13g2_inv_4 clkload14 (.A(clknet_leaf_3_clk));
 sg13g2_inv_1 clkload15 (.A(clknet_leaf_12_clk));
 sg13g2_inv_4 clkload16 (.A(clknet_leaf_15_clk));
 sg13g2_inv_1 clkload17 (.A(clknet_leaf_57_clk));
 sg13g2_inv_1 clkload18 (.A(clknet_leaf_0_clk));
 sg13g2_inv_4 clkload19 (.A(clknet_leaf_1_clk));
 sg13g2_inv_2 clkload20 (.A(clknet_leaf_16_clk));
 sg13g2_inv_1 clkload21 (.A(clknet_leaf_26_clk));
 sg13g2_inv_2 clkload22 (.A(clknet_leaf_24_clk));
 sg13g2_inv_2 clkload23 (.A(clknet_leaf_28_clk));
 sg13g2_inv_1 clkload24 (.A(clknet_leaf_33_clk));
 sg13g2_inv_2 clkload25 (.A(clknet_leaf_52_clk));
 sg13g2_inv_4 clkload26 (.A(clknet_leaf_53_clk));
 sg13g2_inv_4 clkload27 (.A(clknet_leaf_6_clk));
 sg13g2_inv_4 clkload28 (.A(clknet_leaf_7_clk));
 sg13g2_inv_2 clkload29 (.A(clknet_leaf_49_clk));
 sg13g2_inv_2 clkload30 (.A(clknet_leaf_30_clk));
 sg13g2_inv_1 clkload31 (.A(clknet_leaf_48_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\gamepad_pmod.driver.pmod_clk_sync[1] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold2 (.A(\gamepad_pmod.driver.pmod_latch_sync[1] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0170_),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0175_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0173_),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold6 (.A(\gamepad_pmod.driver.pmod_clk_sync[0] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0174_),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0172_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0169_),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold10 (.A(\lfsr_inst.lfsr[26] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold11 (.A(\lfsr_inst.lfsr[20] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold12 (.A(\lfsr_inst.lfsr[22] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold13 (.A(\lfsr_inst.lfsr[16] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold14 (.A(\lfsr_inst.lfsr[19] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold15 (.A(\lfsr_inst.lfsr[25] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold16 (.A(\lfsr_inst.lfsr[23] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0168_),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0270_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold19 (.A(\gamepad_pmod.driver.pmod_latch_sync[0] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold20 (.A(\lfsr_inst.lfsr[18] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold21 (.A(\lfsr_inst.lfsr[27] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold22 (.A(\game_logic_inst.lfsr_value[10] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0163_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0476_),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0097_),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold26 (.A(_3773_),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0449_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold28 (.A(\lfsr_inst.lfsr[24] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold29 (.A(\game_logic_inst.lfsr_value[2] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold30 (.A(\lfsr_inst.lfsr[17] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0085_),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0265_),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold33 (.A(\game_logic_inst.lfsr_value[4] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold34 (.A(\debug_controller_inst.grid_in[15] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0198_),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold36 (.A(\draw_game_inst.new_tiles[0] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold37 (.A(_3394_),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold38 (.A(\game_logic_inst.lfsr_value[3] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold39 (.A(\game_logic_inst.lfsr_value[8] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold40 (.A(\game_logic_inst.lfsr_value[6] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold41 (.A(\game_logic_inst.lfsr_value[9] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold42 (.A(\game_logic_inst.lfsr_value[14] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold43 (.A(\game_logic_inst.lfsr_value[7] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold44 (.A(\lfsr_inst.lfsr[21] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold45 (.A(\btn_right_debounce.debounce_counter[17] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0351_),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold47 (.A(\game_logic_inst.lfsr_value[12] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold48 (.A(\draw_game_inst.grid[45] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0228_),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold50 (.A(\gamepad_pmod.decoder.data_reg[2] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0417_),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold52 (.A(\gamepad_pmod.decoder.data_reg[11] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0426_),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold54 (.A(\gamepad_pmod.decoder.data_reg[3] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0418_),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold56 (.A(\draw_game_inst.grid[62] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold57 (.A(_3384_),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold58 (.A(\draw_game_inst.new_tiles[1] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0250_),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold60 (.A(\game_logic_inst.lfsr_value[5] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold61 (.A(\game_logic_inst.lfsr_value[11] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold62 (.A(\gamepad_pmod.driver.shift_reg[7] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0363_),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold64 (.A(\game_logic_inst.lfsr_value[15] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold65 (.A(\draw_game_inst.grid[34] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold66 (.A(_3328_),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold67 (.A(\draw_game_inst.grid[2] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold68 (.A(_3264_),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold69 (.A(\draw_game_inst.grid[35] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0218_),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold71 (.A(\gamepad_pmod.driver.pmod_data_sync[1] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0355_),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold73 (.A(\draw_game_inst.grid[46] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold74 (.A(_3352_),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold75 (.A(\draw_game_inst.grid[33] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0216_),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold77 (.A(\btn_down_debounce.debounce_counter[17] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold78 (.A(_3542_),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0310_),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold80 (.A(\draw_game_inst.grid[6] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold81 (.A(_3272_),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold82 (.A(\gamepad_pmod.decoder.data_reg[1] ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0416_),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold84 (.A(\draw_game_inst.new_tiles[7] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0256_),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold86 (.A(\btn_up_debounce.debounce_counter[2] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold87 (.A(_3472_),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0274_),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold89 (.A(\btn_left_debounce.debounce_counter[2] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold90 (.A(_3557_),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0315_),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold92 (.A(\draw_game_inst.grid[10] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold93 (.A(_3280_),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold94 (.A(\btn_down_debounce.button_sync_0 ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold95 (.A(\btn_left_debounce.debounce_counter[10] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold96 (.A(_3571_),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0323_),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold98 (.A(\draw_game_inst.grid[1] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0184_),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold100 (.A(\draw_game_inst.grid[41] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0224_),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold102 (.A(\draw_game_inst.grid[54] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold103 (.A(_3368_),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold104 (.A(\draw_game_inst.grid[37] ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0220_),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold106 (.A(\draw_game_inst.grid[0] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0183_),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold108 (.A(\draw_game_inst.grid[39] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0222_),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold110 (.A(\draw_game_inst.new_tiles[10] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0259_),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold112 (.A(\draw_game_inst.grid[42] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold113 (.A(_3344_),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold114 (.A(\draw_game_inst.grid[47] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0230_),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold116 (.A(\gamepad_pmod.decoder.data_reg[10] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0425_),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold118 (.A(\draw_game_inst.grid[55] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0238_),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold120 (.A(\draw_game_inst.grid[38] ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold121 (.A(_3336_),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold122 (.A(\draw_game_inst.grid[43] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0226_),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold124 (.A(\draw_game_inst.grid[59] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0242_),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold126 (.A(\draw_game_inst.grid[32] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0215_),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold128 (.A(\draw_game_inst.grid[14] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold129 (.A(_3288_),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold130 (.A(\draw_game_inst.grid[52] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0235_),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold132 (.A(\game_logic_inst.lfsr_value[13] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold133 (.A(\draw_game_inst.grid[63] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0246_),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold135 (.A(\gamepad_pmod.decoder.data_reg[0] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0415_),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold137 (.A(\draw_game_inst.grid[16] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0199_),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold139 (.A(\draw_game_inst.grid[18] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold140 (.A(_3296_),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold141 (.A(\draw_game_inst.grid[61] ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0244_),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold143 (.A(\draw_game_inst.grid[53] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0236_),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold145 (.A(\draw_game_inst.grid[12] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0195_),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold147 (.A(\draw_game_inst.grid[36] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0219_),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold149 (.A(\draw_game_inst.grid[21] ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0204_),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold151 (.A(\btn_right_debounce.debounce_counter[10] ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold152 (.A(_3613_),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0344_),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold154 (.A(\draw_game_inst.grid[50] ),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold155 (.A(_3360_),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold156 (.A(\draw_game_inst.new_tiles[13] ),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0262_),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold158 (.A(\draw_game_inst.grid[51] ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0234_),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0080_),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0260_),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold162 (.A(\draw_game_inst.grid[13] ),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0196_),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold164 (.A(\draw_game_inst.grid[58] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold165 (.A(_3376_),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold166 (.A(\btn_right_debounce.debounce_counter[2] ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold167 (.A(_3599_),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0336_),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold169 (.A(\btn_down_debounce.debounce_counter[16] ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0309_),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold171 (.A(\draw_game_inst.grid[9] ),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0192_),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold173 (.A(\btn_right_debounce.debounce_counter[16] ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold174 (.A(_3623_),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0350_),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold176 (.A(\draw_game_inst.grid[25] ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0208_),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold178 (.A(\btn_up_debounce.debounce_counter[10] ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold179 (.A(_3486_),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0282_),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold181 (.A(\vga_sync_gen.vsync ),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold182 (.A(\draw_game_inst.grid[3] ),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0186_),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold184 (.A(\draw_game_inst.grid[28] ),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0211_),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold186 (.A(\btn_down_debounce.debounce_counter[10] ),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold187 (.A(_3530_),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0303_),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold189 (.A(\draw_game_inst.grid[19] ),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0202_),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold191 (.A(\draw_game_inst.new_tiles[2] ),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0251_),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold193 (.A(\btn_down_debounce.debounce_counter[12] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold194 (.A(_3533_),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0305_),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold196 (.A(\draw_game_inst.new_tiles[3] ),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0252_),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold198 (.A(\draw_game_inst.grid[31] ),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0214_),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold200 (.A(\draw_game_inst.grid[20] ),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0203_),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold202 (.A(\draw_game_inst.grid[29] ),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0212_),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold204 (.A(\draw_game_inst.grid[44] ),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0227_),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold206 (.A(\draw_game_inst.grid[24] ),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0207_),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold208 (.A(\draw_game_inst.grid[22] ),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold209 (.A(_3304_),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold210 (.A(\gamepad_pmod.driver.shift_reg[11] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0366_),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold212 (.A(\btn_left_debounce.debounce_counter[12] ),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold213 (.A(_3574_),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0325_),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold215 (.A(\draw_game_inst.grid[26] ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold216 (.A(_3312_),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold217 (.A(\draw_game_inst.grid[8] ),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0191_),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold219 (.A(\game_logic_inst.current_direction[1] ),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0000_),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold221 (.A(\draw_game_inst.grid[56] ),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0239_),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold223 (.A(\draw_game_inst.grid[27] ),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0210_),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold225 (.A(_0073_),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold226 (.A(_0253_),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold227 (.A(\draw_game_inst.new_tiles[9] ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold228 (.A(_0258_),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold229 (.A(\draw_game_inst.grid[57] ),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0240_),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold231 (.A(\draw_game_inst.grid[23] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold232 (.A(_0206_),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold233 (.A(\gamepad_pmod.decoder.data_reg[4] ),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold234 (.A(_0419_),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold235 (.A(_0084_),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0264_),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold237 (.A(\btn_up_debounce.debounce_counter[12] ),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold238 (.A(_3489_),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold239 (.A(_0284_),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0081_),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold241 (.A(_3432_),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0261_),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold243 (.A(\draw_game_inst.grid[30] ),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold244 (.A(_3320_),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold245 (.A(\draw_game_inst.grid[17] ),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold246 (.A(_0200_),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold247 (.A(\gamepad_pmod.driver.shift_reg[5] ),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold248 (.A(_0361_),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold249 (.A(\welcome_screen_grid[32] ),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold250 (.A(_0486_),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0077_),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold252 (.A(_0257_),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold253 (.A(\draw_game_inst.grid[40] ),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold254 (.A(_0223_),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold255 (.A(\btn_right_debounce.debounce_counter[12] ),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold256 (.A(_3616_),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold257 (.A(_0346_),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold258 (.A(_0098_),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold259 (.A(_3786_),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold260 (.A(\draw_game_inst.grid[11] ),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold261 (.A(_0194_),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold262 (.A(\gamepad_pmod.decoder.data_reg[6] ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold263 (.A(_0421_),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold264 (.A(\draw_game_inst.grid[49] ),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold265 (.A(_0232_),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold266 (.A(\draw_game_inst.grid[4] ),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold267 (.A(_0187_),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold268 (.A(\gamepad_pmod.decoder.data_reg[5] ),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold269 (.A(\game_logic_inst.lfsr_value[0] ),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold270 (.A(\btn_right_debounce.debounced ),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold271 (.A(_0353_),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold272 (.A(\btn_right_debounce.debounce_counter[15] ),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold273 (.A(_0349_),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold274 (.A(\new_tiles_counter[4] ),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold275 (.A(_3458_),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold276 (.A(\draw_game_inst.grid[7] ),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold277 (.A(_0190_),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold278 (.A(\draw_game_inst.grid[48] ),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold279 (.A(_0231_),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold280 (.A(\welcome_screen_grid[11] ),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold281 (.A(_0485_),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold282 (.A(\draw_game_inst.grid[5] ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold283 (.A(_0188_),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold284 (.A(\btn_down_debounce.debounce_counter[4] ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold285 (.A(_3520_),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold286 (.A(\btn_down_debounce.debounce_counter[5] ),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold287 (.A(_0298_),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold288 (.A(\gamepad_pmod.decoder.data_reg[9] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold289 (.A(_0424_),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold290 (.A(\gamepad_pmod.decoder.data_reg[7] ),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold291 (.A(\draw_game_inst.grid[60] ),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold292 (.A(_0243_),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold293 (.A(\btn_down_debounce.debounce_counter[3] ),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold294 (.A(_3518_),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold295 (.A(_0296_),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold296 (.A(\btn_up_debounce.debounce_counter[5] ),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold297 (.A(_3478_),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold298 (.A(_0277_),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold299 (.A(\gamepad_pmod.driver.shift_reg[0] ),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold300 (.A(_0356_),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold301 (.A(\welcome_screen_grid[40] ),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold302 (.A(_0484_),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold303 (.A(\draw_game_inst.new_tiles[6] ),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold304 (.A(_0255_),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold305 (.A(\btn_up_debounce.debounce_counter[17] ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold306 (.A(_3499_),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold307 (.A(_0289_),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold308 (.A(\welcome_screen_grid[44] ),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold309 (.A(_0483_),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold310 (.A(\btn_up_debounce.debounce_counter[7] ),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold311 (.A(_3481_),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold312 (.A(\gamepad_pmod.driver.shift_reg[4] ),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold313 (.A(\btn_down_debounce.debounce_counter[2] ),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold314 (.A(_3516_),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold315 (.A(_0295_),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold316 (.A(\btn_up_debounce.debounce_counter[6] ),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold317 (.A(\btn_down_debounce.debounce_counter[13] ),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold318 (.A(_3535_),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold319 (.A(\btn_up_debounce.debounce_counter[15] ),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold320 (.A(_3495_),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold321 (.A(\btn_up_debounce.debounce_counter[4] ),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold322 (.A(_3476_),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold323 (.A(\btn_down_debounce.debounce_counter[8] ),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold324 (.A(_3527_),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold325 (.A(\btn_left_debounce.debounce_counter[3] ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold326 (.A(_3559_),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold327 (.A(\btn_left_debounce.debounce_counter[17] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold328 (.A(_3584_),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold329 (.A(_0330_),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold330 (.A(\draw_game_inst.new_tiles[14] ),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold331 (.A(_0263_),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold332 (.A(\btn_right_debounce.debounce_counter[6] ),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold333 (.A(_3606_),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold334 (.A(_0340_),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold335 (.A(\btn_right_debounce.debounce_counter[4] ),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold336 (.A(_3603_),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold337 (.A(_0338_),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold338 (.A(\draw_game_inst.board_y[6] ),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold339 (.A(\btn_left_debounce.debounce_counter[4] ),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold340 (.A(\welcome_screen_grid[0] ),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold341 (.A(_0487_),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold342 (.A(\game_logic_inst.lfsr_value[1] ),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold343 (.A(\gamepad_pmod.decoder.data_reg[8] ),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold344 (.A(_0423_),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold345 (.A(\btn_right_debounce.debounce_counter[5] ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold346 (.A(_0339_),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold347 (.A(\btn_left_debounce.debounce_counter[6] ),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold348 (.A(_3564_),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold349 (.A(\btn_left_debounce.debounce_counter[13] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold350 (.A(_3576_),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold351 (.A(\gamepad_pmod.driver.shift_reg[10] ),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold352 (.A(_0365_),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold353 (.A(\gamepad_pmod.driver.shift_reg[6] ),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold354 (.A(\btn_down_debounce.button_sync_1 ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold355 (.A(_0311_),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold356 (.A(\gamepad_pmod.driver.shift_reg[3] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold357 (.A(_0358_),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold358 (.A(\gamepad_pmod.driver.shift_reg[9] ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold359 (.A(_0364_),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold360 (.A(\btn_right_debounce.debounce_counter[13] ),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold361 (.A(_3618_),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold362 (.A(_0347_),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold363 (.A(\welcome_screen_grid[4] ),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold364 (.A(_0495_),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold365 (.A(\btn_left_debounce.debounce_counter[7] ),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold366 (.A(\btn_up_debounce.debounce_counter[3] ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold367 (.A(_3474_),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold368 (.A(\gamepad_pmod.driver.pmod_clk_prev ),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold369 (.A(\btn_left_debounce.debounce_counter[14] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold370 (.A(\gamepad_pmod.driver.shift_reg[2] ),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold371 (.A(_0357_),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold372 (.A(\btn_right_debounce.debounce_counter[3] ),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold373 (.A(_3601_),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold374 (.A(_0337_),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold375 (.A(\btn_left_debounce.debounce_counter[5] ),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold376 (.A(_0318_),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold377 (.A(\draw_game_inst.new_tiles[5] ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold378 (.A(_0254_),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold379 (.A(\welcome_screen_grid[36] ),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold380 (.A(_0489_),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold381 (.A(\game_logic_inst.add_new_tiles[0] ),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold382 (.A(_0448_),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold383 (.A(\draw_game_inst.new_tiles_counter[0] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold384 (.A(_3449_),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold385 (.A(\btn_up_debounce.debounce_counter[14] ),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold386 (.A(_3493_),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold387 (.A(\welcome_screen_inst.welcome_counter[1] ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold388 (.A(_0438_),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold389 (.A(\welcome_screen_inst.welcome_counter[2] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold390 (.A(_0439_),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold391 (.A(\btn_up_debounce.debounce_counter[8] ),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold392 (.A(\btn_down_debounce.debounce_counter[6] ),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold393 (.A(\btn_right_debounce.debounce_counter[8] ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold394 (.A(_3610_),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold395 (.A(\btn_left_debounce.debounce_counter[15] ),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold396 (.A(\btn_right_debounce.debounce_counter[7] ),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold397 (.A(_0341_),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold398 (.A(\welcome_screen_grid[12] ),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold399 (.A(_0494_),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold400 (.A(\btn_up_debounce.debounce_counter[13] ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold401 (.A(_3491_),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold402 (.A(\btn_up_debounce.debounce_counter[16] ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold403 (.A(\btn_left_debounce.debounce_counter[16] ),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold404 (.A(\welcome_screen_grid[56] ),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold405 (.A(_0481_),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold406 (.A(\btn_left_debounce.debounce_counter[8] ),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold407 (.A(\btn_down_debounce.debounce_counter[7] ),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold408 (.A(\btn_left_debounce.debounced ),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold409 (.A(_0332_),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold410 (.A(\btn_up_debounce.debounce_counter[0] ),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold411 (.A(_3470_),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold412 (.A(\game_logic_inst.debug_move_reg ),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold413 (.A(_0442_),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold414 (.A(\draw_game_inst.board_x[2] ),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold415 (.A(_0429_),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold416 (.A(\btn_right_debounce.debounce_counter[0] ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold417 (.A(_3597_),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold418 (.A(_0335_),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold419 (.A(\welcome_screen_inst.welcome_counter[4] ),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold420 (.A(_3715_),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold421 (.A(_0441_),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold422 (.A(\draw_game_inst.new_tiles_counter[1] ),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold423 (.A(_0267_),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold424 (.A(\btn_left_debounce.debounce_counter[11] ),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold425 (.A(_3573_),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold426 (.A(\welcome_screen_grid[20] ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold427 (.A(_0488_),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold428 (.A(_0087_),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold429 (.A(_3457_),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold430 (.A(_0268_),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold431 (.A(\btn_left_debounce.debounce_counter[9] ),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold432 (.A(_0322_),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold433 (.A(_0089_),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold434 (.A(\btn_right_debounce.debounce_counter[11] ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold435 (.A(_3615_),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold436 (.A(\welcome_screen_grid[52] ),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold437 (.A(_0480_),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold438 (.A(\btn_up_debounce.debounce_counter[9] ),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold439 (.A(\btn_down_debounce.debounce_counter[11] ),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold440 (.A(_3532_),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold441 (.A(\welcome_screen_grid[28] ),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold442 (.A(_0492_),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold443 (.A(\welcome_screen_grid[60] ),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold444 (.A(_0482_),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold445 (.A(\welcome_screen_grid[16] ),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold446 (.A(_0490_),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold447 (.A(\btn_left_debounce.debounce_counter[1] ),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold448 (.A(_3555_),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold449 (.A(uio_out[5]),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold450 (.A(uio_out[6]),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold451 (.A(\btn_up_debounce.debounce_counter[11] ),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold452 (.A(\btn_down_debounce.debounce_counter[14] ),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold453 (.A(\btn_down_debounce.debounce_counter[9] ),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold454 (.A(_0124_),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold455 (.A(_1304_),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold456 (.A(\btn_down_debounce.debounce_counter[1] ),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold457 (.A(_3503_),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold458 (.A(_0294_),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold459 (.A(\btn_down_debounce.debounce_counter[15] ),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold460 (.A(\btn_right_debounce.debounce_counter[9] ),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold461 (.A(\btn_up_debounce.debounced ),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold462 (.A(_0291_),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold463 (.A(_0122_),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold464 (.A(\welcome_screen_grid[24] ),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold465 (.A(_0493_),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold466 (.A(_0120_),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold467 (.A(_1293_),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold468 (.A(\draw_game_inst.y[8] ),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold469 (.A(\welcome_screen_grid[48] ),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold470 (.A(_0491_),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold471 (.A(\lfsr_inst.lfsr[30] ),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold472 (.A(\game_logic_inst.should_transpose ),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold473 (.A(_0455_),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold474 (.A(\btn_right_debounce.debounce_counter[14] ),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold475 (.A(\btn_up_debounce.button_sync_0 ),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold476 (.A(_0125_),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold477 (.A(_1305_),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold478 (.A(_1309_),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold479 (.A(uio_out[4]),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold480 (.A(\debug_controller_inst.grid_out_addr[3] ),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold481 (.A(\draw_game_inst.y[9] ),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold482 (.A(uio_out[7]),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold483 (.A(_0142_),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold484 (.A(_0051_),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold485 (.A(_0107_),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold486 (.A(_0915_),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold487 (.A(_0111_),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold488 (.A(_0948_),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold489 (.A(_0065_),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold490 (.A(_0102_),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold491 (.A(_0036_),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold492 (.A(_0105_),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold493 (.A(_0899_),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold494 (.A(_0156_),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold495 (.A(_0056_),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold496 (.A(_0130_),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold497 (.A(_1088_),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold498 (.A(_0018_),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold499 (.A(_0104_),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold500 (.A(_0166_),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold501 (.A(_0457_),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold502 (.A(_0149_),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold503 (.A(_0039_),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold504 (.A(_0113_),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold505 (.A(_0958_),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold506 (.A(_0066_),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold507 (.A(_0150_),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold508 (.A(_0040_),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold509 (.A(_0109_),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold510 (.A(_0162_),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold511 (.A(_1389_),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold512 (.A(\lfsr_inst.lfsr[31] ),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold513 (.A(_0101_),
    .X(net928));
 sg13g2_dlygate4sd3_1 hold514 (.A(_0025_),
    .X(net929));
 sg13g2_dlygate4sd3_1 hold515 (.A(_0133_),
    .X(net930));
 sg13g2_dlygate4sd3_1 hold516 (.A(_1108_),
    .X(net931));
 sg13g2_dlygate4sd3_1 hold517 (.A(_0020_),
    .X(net932));
 sg13g2_dlygate4sd3_1 hold518 (.A(_0148_),
    .X(net933));
 sg13g2_dlygate4sd3_1 hold519 (.A(_0038_),
    .X(net934));
 sg13g2_dlygate4sd3_1 hold520 (.A(_0103_),
    .X(net935));
 sg13g2_dlygate4sd3_1 hold521 (.A(_0100_),
    .X(net936));
 sg13g2_dlygate4sd3_1 hold522 (.A(_0791_),
    .X(net937));
 sg13g2_dlygate4sd3_1 hold523 (.A(_0014_),
    .X(net938));
 sg13g2_dlygate4sd3_1 hold524 (.A(_0139_),
    .X(net939));
 sg13g2_dlygate4sd3_1 hold525 (.A(\debug_controller_inst.grid_out_data[1] ),
    .X(net940));
 sg13g2_dlygate4sd3_1 hold526 (.A(_0042_),
    .X(net941));
 sg13g2_dlygate4sd3_1 hold527 (.A(_0117_),
    .X(net942));
 sg13g2_dlygate4sd3_1 hold528 (.A(_0976_),
    .X(net943));
 sg13g2_dlygate4sd3_1 hold529 (.A(_0005_),
    .X(net944));
 sg13g2_dlygate4sd3_1 hold530 (.A(\draw_game_inst.x[9] ),
    .X(net945));
 sg13g2_dlygate4sd3_1 hold531 (.A(_0146_),
    .X(net946));
 sg13g2_dlygate4sd3_1 hold532 (.A(_1331_),
    .X(net947));
 sg13g2_dlygate4sd3_1 hold533 (.A(_0129_),
    .X(net948));
 sg13g2_dlygate4sd3_1 hold534 (.A(_0143_),
    .X(net949));
 sg13g2_dlygate4sd3_1 hold535 (.A(_1153_),
    .X(net950));
 sg13g2_dlygate4sd3_1 hold536 (.A(\debug_controller_inst.grid_addr[2] ),
    .X(net951));
 sg13g2_dlygate4sd3_1 hold537 (.A(_0473_),
    .X(net952));
 sg13g2_dlygate4sd3_1 hold538 (.A(_0145_),
    .X(net953));
 sg13g2_dlygate4sd3_1 hold539 (.A(_1161_),
    .X(net954));
 sg13g2_dlygate4sd3_1 hold540 (.A(\game_logic_inst.current_direction[2] ),
    .X(net955));
 sg13g2_dlygate4sd3_1 hold541 (.A(_0001_),
    .X(net956));
 sg13g2_dlygate4sd3_1 hold542 (.A(_0127_),
    .X(net957));
 sg13g2_dlygate4sd3_1 hold543 (.A(_0161_),
    .X(net958));
 sg13g2_dlygate4sd3_1 hold544 (.A(_0099_),
    .X(net959));
 sg13g2_dlygate4sd3_1 hold545 (.A(_0003_),
    .X(net960));
 sg13g2_dlygate4sd3_1 hold546 (.A(_0160_),
    .X(net961));
 sg13g2_dlygate4sd3_1 hold547 (.A(_0171_),
    .X(net962));
 sg13g2_dlygate4sd3_1 hold548 (.A(_0131_),
    .X(net963));
 sg13g2_dlygate4sd3_1 hold549 (.A(_0019_),
    .X(net964));
 sg13g2_dlygate4sd3_1 hold550 (.A(_0147_),
    .X(net965));
 sg13g2_dlygate4sd3_1 hold551 (.A(_0128_),
    .X(net966));
 sg13g2_dlygate4sd3_1 hold552 (.A(_0115_),
    .X(net967));
 sg13g2_dlygate4sd3_1 hold553 (.A(_0967_),
    .X(net968));
 sg13g2_dlygate4sd3_1 hold554 (.A(_0004_),
    .X(net969));
 sg13g2_dlygate4sd3_1 hold555 (.A(_0144_),
    .X(net970));
 sg13g2_dlygate4sd3_1 hold556 (.A(_1326_),
    .X(net971));
 sg13g2_dlygate4sd3_1 hold557 (.A(_0052_),
    .X(net972));
 sg13g2_dlygate4sd3_1 hold558 (.A(_0141_),
    .X(net973));
 sg13g2_dlygate4sd3_1 hold559 (.A(_0158_),
    .X(net974));
 sg13g2_dlygate4sd3_1 hold560 (.A(_1356_),
    .X(net975));
 sg13g2_dlygate4sd3_1 hold561 (.A(_0057_),
    .X(net976));
 sg13g2_dlygate4sd3_1 hold562 (.A(_0135_),
    .X(net977));
 sg13g2_dlygate4sd3_1 hold563 (.A(_1116_),
    .X(net978));
 sg13g2_dlygate4sd3_1 hold564 (.A(_0021_),
    .X(net979));
 sg13g2_dlygate4sd3_1 hold565 (.A(_0140_),
    .X(net980));
 sg13g2_dlygate4sd3_1 hold566 (.A(_0106_),
    .X(net981));
 sg13g2_dlygate4sd3_1 hold567 (.A(\debug_controller_inst.grid_addr[0] ),
    .X(net982));
 sg13g2_dlygate4sd3_1 hold568 (.A(\debug_controller_inst.grid_out_data[2] ),
    .X(net983));
 sg13g2_dlygate4sd3_1 hold569 (.A(_0043_),
    .X(net984));
 sg13g2_dlygate4sd3_1 hold570 (.A(_0137_),
    .X(net985));
 sg13g2_dlygate4sd3_1 hold571 (.A(_1124_),
    .X(net986));
 sg13g2_dlygate4sd3_1 hold572 (.A(_0022_),
    .X(net987));
 sg13g2_dlygate4sd3_1 hold573 (.A(\gamepad_pmod.driver.pmod_data_sync[0] ),
    .X(net988));
 sg13g2_dlygate4sd3_1 hold574 (.A(_0112_),
    .X(net989));
 sg13g2_dlygate4sd3_1 hold575 (.A(_0028_),
    .X(net990));
 sg13g2_dlygate4sd3_1 hold576 (.A(\debug_controller_inst.grid_out_data[0] ),
    .X(net991));
 sg13g2_dlygate4sd3_1 hold577 (.A(_0041_),
    .X(net992));
 sg13g2_dlygate4sd3_1 hold578 (.A(\game_logic_inst.lfsr_shift[1] ),
    .X(net993));
 sg13g2_dlygate4sd3_1 hold579 (.A(_3756_),
    .X(net994));
 sg13g2_dlygate4sd3_1 hold580 (.A(\draw_game_inst.board_x[1] ),
    .X(net995));
 sg13g2_dlygate4sd3_1 hold581 (.A(_3215_),
    .X(net996));
 sg13g2_dlygate4sd3_1 hold582 (.A(_0110_),
    .X(net997));
 sg13g2_dlygate4sd3_1 hold583 (.A(\draw_game_inst.board_x[0] ),
    .X(net998));
 sg13g2_dlygate4sd3_1 hold584 (.A(_0428_),
    .X(net999));
 sg13g2_dlygate4sd3_1 hold585 (.A(_0108_),
    .X(net1000));
 sg13g2_dlygate4sd3_1 hold586 (.A(_0132_),
    .X(net1001));
 sg13g2_dlygate4sd3_1 hold587 (.A(_0165_),
    .X(net1002));
 sg13g2_dlygate4sd3_1 hold588 (.A(_0513_),
    .X(net1003));
 sg13g2_dlygate4sd3_1 hold589 (.A(_0527_),
    .X(net1004));
 sg13g2_dlygate4sd3_1 hold590 (.A(\welcome_screen_inst.welcome_counter[3] ),
    .X(net1005));
 sg13g2_dlygate4sd3_1 hold591 (.A(_3712_),
    .X(net1006));
 sg13g2_dlygate4sd3_1 hold592 (.A(\draw_game_inst.x[8] ),
    .X(net1007));
 sg13g2_dlygate4sd3_1 hold593 (.A(_0154_),
    .X(net1008));
 sg13g2_dlygate4sd3_1 hold594 (.A(\lfsr_inst.lfsr[28] ),
    .X(net1009));
 sg13g2_dlygate4sd3_1 hold595 (.A(\lfsr_inst.lfsr[29] ),
    .X(net1010));
 sg13g2_dlygate4sd3_1 hold596 (.A(_0164_),
    .X(net1011));
 sg13g2_dlygate4sd3_1 hold597 (.A(_3900_),
    .X(net1012));
 sg13g2_dlygate4sd3_1 hold598 (.A(\btn_left_debounce.button_sync_0 ),
    .X(net1013));
 sg13g2_dlygate4sd3_1 hold599 (.A(\welcome_screen_inst.welcome_counter[0] ),
    .X(net1014));
 sg13g2_dlygate4sd3_1 hold600 (.A(\draw_game_inst.x[6] ),
    .X(net1015));
 sg13g2_dlygate4sd3_1 hold601 (.A(_0152_),
    .X(net1016));
 sg13g2_dlygate4sd3_1 hold602 (.A(_0116_),
    .X(net1017));
 sg13g2_dlygate4sd3_1 hold603 (.A(_1185_),
    .X(net1018));
 sg13g2_dlygate4sd3_1 hold604 (.A(_0136_),
    .X(net1019));
 sg13g2_dlygate4sd3_1 hold605 (.A(_0118_),
    .X(net1020));
 sg13g2_dlygate4sd3_1 hold606 (.A(_1191_),
    .X(net1021));
 sg13g2_dlygate4sd3_1 hold607 (.A(_0031_),
    .X(net1022));
 sg13g2_dlygate4sd3_1 hold608 (.A(_0114_),
    .X(net1023));
 sg13g2_dlygate4sd3_1 hold609 (.A(_1179_),
    .X(net1024));
 sg13g2_dlygate4sd3_1 hold610 (.A(\draw_game_inst.board_y[2] ),
    .X(net1025));
 sg13g2_dlygate4sd3_1 hold611 (.A(\btn_right_debounce.button_sync_0 ),
    .X(net1026));
 sg13g2_dlygate4sd3_1 hold612 (.A(_0123_),
    .X(net1027));
 sg13g2_dlygate4sd3_1 hold613 (.A(_0119_),
    .X(net1028));
 sg13g2_dlygate4sd3_1 hold614 (.A(_0138_),
    .X(net1029));
 sg13g2_dlygate4sd3_1 hold615 (.A(_0035_),
    .X(net1030));
 sg13g2_dlygate4sd3_1 hold616 (.A(\debug_controller_inst.grid_addr[1] ),
    .X(net1031));
 sg13g2_dlygate4sd3_1 hold617 (.A(\debug_controller_inst.grid_out_data[3] ),
    .X(net1032));
 sg13g2_dlygate4sd3_1 hold618 (.A(_0134_),
    .X(net1033));
 sg13g2_dlygate4sd3_1 hold619 (.A(\gamepad_pmod.decoder.data_reg[6] ),
    .X(net1034));
 sg13g2_dlygate4sd3_1 hold620 (.A(_0121_),
    .X(net1035));
 sg13g2_dlygate4sd3_1 hold621 (.A(_0157_),
    .X(net1036));
 sg13g2_dlygate4sd3_1 hold622 (.A(\draw_game_inst.new_tiles_counter[2] ),
    .X(net1037));
 sg13g2_dlygate4sd3_1 hold623 (.A(_0179_),
    .X(net1038));
 sg13g2_dlygate4sd3_1 hold624 (.A(_0159_),
    .X(net1039));
 sg13g2_dlygate4sd3_1 hold625 (.A(\draw_game_inst.x[9] ),
    .X(net1040));
 sg13g2_dlygate4sd3_1 hold626 (.A(\game_logic_inst.valid_move ),
    .X(net1041));
 sg13g2_dlygate4sd3_1 hold627 (.A(\draw_game_inst.y[9] ),
    .X(net1042));
 sg13g2_dlygate4sd3_1 hold628 (.A(_3249_),
    .X(net1043));
 sg13g2_dlygate4sd3_1 hold629 (.A(_0086_),
    .X(net1044));
 sg13g2_dlygate4sd3_1 hold630 (.A(_0121_),
    .X(net1045));
 sg13g2_dlygate4sd3_1 hold631 (.A(_0140_),
    .X(net1046));
 sg13g2_dlygate4sd3_1 hold632 (.A(_0110_),
    .X(net1047));
 sg13g2_dlygate4sd3_1 hold633 (.A(_0110_),
    .X(net1048));
 sg13g2_antennanp ANTENNA_1 (.A(\btn_left_debounce.button_sync_0 ));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_fill_1 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_fill_1 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_fill_1 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_fill_1 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_fill_1 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_8 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_707 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_8 FILLER_5_728 ();
 sg13g2_decap_8 FILLER_5_735 ();
 sg13g2_decap_8 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_8 FILLER_5_756 ();
 sg13g2_decap_8 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_8 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_8 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_854 ();
 sg13g2_fill_1 FILLER_5_861 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_518 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_8 FILLER_6_539 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_8 FILLER_6_553 ();
 sg13g2_decap_8 FILLER_6_560 ();
 sg13g2_decap_8 FILLER_6_567 ();
 sg13g2_decap_8 FILLER_6_574 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_decap_8 FILLER_6_595 ();
 sg13g2_decap_8 FILLER_6_602 ();
 sg13g2_decap_8 FILLER_6_609 ();
 sg13g2_decap_8 FILLER_6_616 ();
 sg13g2_decap_8 FILLER_6_623 ();
 sg13g2_decap_8 FILLER_6_630 ();
 sg13g2_decap_8 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_651 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_decap_8 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_679 ();
 sg13g2_decap_8 FILLER_6_686 ();
 sg13g2_decap_8 FILLER_6_693 ();
 sg13g2_decap_8 FILLER_6_700 ();
 sg13g2_decap_8 FILLER_6_707 ();
 sg13g2_decap_8 FILLER_6_714 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_decap_8 FILLER_6_742 ();
 sg13g2_decap_8 FILLER_6_749 ();
 sg13g2_decap_8 FILLER_6_756 ();
 sg13g2_decap_8 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_777 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_833 ();
 sg13g2_decap_8 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_6_847 ();
 sg13g2_decap_8 FILLER_6_854 ();
 sg13g2_fill_1 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_fill_1 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_8 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_546 ();
 sg13g2_decap_8 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_560 ();
 sg13g2_decap_8 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_decap_8 FILLER_8_581 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_decap_8 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_623 ();
 sg13g2_decap_8 FILLER_8_630 ();
 sg13g2_decap_8 FILLER_8_637 ();
 sg13g2_decap_8 FILLER_8_644 ();
 sg13g2_decap_8 FILLER_8_651 ();
 sg13g2_decap_8 FILLER_8_658 ();
 sg13g2_decap_8 FILLER_8_665 ();
 sg13g2_decap_8 FILLER_8_672 ();
 sg13g2_decap_8 FILLER_8_679 ();
 sg13g2_decap_8 FILLER_8_686 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_8 FILLER_8_700 ();
 sg13g2_decap_8 FILLER_8_707 ();
 sg13g2_decap_8 FILLER_8_714 ();
 sg13g2_decap_8 FILLER_8_721 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_decap_8 FILLER_8_735 ();
 sg13g2_decap_8 FILLER_8_742 ();
 sg13g2_decap_8 FILLER_8_749 ();
 sg13g2_decap_8 FILLER_8_756 ();
 sg13g2_decap_8 FILLER_8_763 ();
 sg13g2_decap_8 FILLER_8_770 ();
 sg13g2_decap_8 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_784 ();
 sg13g2_decap_8 FILLER_8_791 ();
 sg13g2_decap_8 FILLER_8_798 ();
 sg13g2_decap_8 FILLER_8_805 ();
 sg13g2_decap_8 FILLER_8_812 ();
 sg13g2_decap_8 FILLER_8_819 ();
 sg13g2_decap_8 FILLER_8_826 ();
 sg13g2_decap_8 FILLER_8_833 ();
 sg13g2_decap_8 FILLER_8_840 ();
 sg13g2_decap_8 FILLER_8_847 ();
 sg13g2_decap_8 FILLER_8_854 ();
 sg13g2_fill_1 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_4 FILLER_9_140 ();
 sg13g2_fill_2 FILLER_9_144 ();
 sg13g2_decap_8 FILLER_9_150 ();
 sg13g2_fill_2 FILLER_9_157 ();
 sg13g2_decap_8 FILLER_9_164 ();
 sg13g2_decap_8 FILLER_9_171 ();
 sg13g2_decap_8 FILLER_9_178 ();
 sg13g2_decap_8 FILLER_9_185 ();
 sg13g2_decap_8 FILLER_9_192 ();
 sg13g2_decap_8 FILLER_9_199 ();
 sg13g2_decap_8 FILLER_9_206 ();
 sg13g2_decap_8 FILLER_9_213 ();
 sg13g2_decap_8 FILLER_9_220 ();
 sg13g2_decap_8 FILLER_9_227 ();
 sg13g2_decap_8 FILLER_9_234 ();
 sg13g2_decap_8 FILLER_9_241 ();
 sg13g2_decap_8 FILLER_9_248 ();
 sg13g2_decap_8 FILLER_9_255 ();
 sg13g2_decap_8 FILLER_9_262 ();
 sg13g2_decap_8 FILLER_9_269 ();
 sg13g2_decap_8 FILLER_9_276 ();
 sg13g2_decap_8 FILLER_9_283 ();
 sg13g2_decap_8 FILLER_9_290 ();
 sg13g2_decap_8 FILLER_9_297 ();
 sg13g2_decap_8 FILLER_9_304 ();
 sg13g2_decap_8 FILLER_9_311 ();
 sg13g2_decap_8 FILLER_9_318 ();
 sg13g2_decap_8 FILLER_9_325 ();
 sg13g2_decap_8 FILLER_9_332 ();
 sg13g2_decap_8 FILLER_9_339 ();
 sg13g2_decap_8 FILLER_9_346 ();
 sg13g2_decap_4 FILLER_9_353 ();
 sg13g2_fill_2 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_375 ();
 sg13g2_decap_8 FILLER_9_382 ();
 sg13g2_decap_8 FILLER_9_389 ();
 sg13g2_decap_8 FILLER_9_396 ();
 sg13g2_decap_8 FILLER_9_403 ();
 sg13g2_decap_8 FILLER_9_410 ();
 sg13g2_decap_8 FILLER_9_417 ();
 sg13g2_decap_8 FILLER_9_424 ();
 sg13g2_decap_8 FILLER_9_431 ();
 sg13g2_decap_8 FILLER_9_438 ();
 sg13g2_decap_8 FILLER_9_445 ();
 sg13g2_decap_8 FILLER_9_452 ();
 sg13g2_decap_8 FILLER_9_459 ();
 sg13g2_decap_8 FILLER_9_466 ();
 sg13g2_decap_8 FILLER_9_473 ();
 sg13g2_decap_8 FILLER_9_480 ();
 sg13g2_decap_8 FILLER_9_487 ();
 sg13g2_decap_8 FILLER_9_494 ();
 sg13g2_decap_8 FILLER_9_501 ();
 sg13g2_decap_8 FILLER_9_508 ();
 sg13g2_decap_8 FILLER_9_515 ();
 sg13g2_decap_8 FILLER_9_522 ();
 sg13g2_fill_2 FILLER_9_529 ();
 sg13g2_fill_1 FILLER_9_531 ();
 sg13g2_decap_8 FILLER_9_542 ();
 sg13g2_decap_8 FILLER_9_549 ();
 sg13g2_decap_8 FILLER_9_556 ();
 sg13g2_decap_8 FILLER_9_563 ();
 sg13g2_decap_8 FILLER_9_570 ();
 sg13g2_decap_8 FILLER_9_577 ();
 sg13g2_decap_8 FILLER_9_584 ();
 sg13g2_decap_8 FILLER_9_591 ();
 sg13g2_decap_8 FILLER_9_598 ();
 sg13g2_decap_8 FILLER_9_605 ();
 sg13g2_decap_8 FILLER_9_612 ();
 sg13g2_decap_8 FILLER_9_619 ();
 sg13g2_decap_8 FILLER_9_626 ();
 sg13g2_decap_8 FILLER_9_633 ();
 sg13g2_decap_8 FILLER_9_640 ();
 sg13g2_decap_8 FILLER_9_647 ();
 sg13g2_decap_8 FILLER_9_654 ();
 sg13g2_decap_8 FILLER_9_661 ();
 sg13g2_decap_8 FILLER_9_668 ();
 sg13g2_decap_8 FILLER_9_675 ();
 sg13g2_decap_8 FILLER_9_682 ();
 sg13g2_decap_8 FILLER_9_689 ();
 sg13g2_decap_8 FILLER_9_696 ();
 sg13g2_decap_8 FILLER_9_703 ();
 sg13g2_decap_8 FILLER_9_710 ();
 sg13g2_decap_8 FILLER_9_717 ();
 sg13g2_decap_8 FILLER_9_724 ();
 sg13g2_decap_8 FILLER_9_731 ();
 sg13g2_decap_8 FILLER_9_738 ();
 sg13g2_decap_8 FILLER_9_745 ();
 sg13g2_decap_8 FILLER_9_752 ();
 sg13g2_decap_8 FILLER_9_759 ();
 sg13g2_decap_8 FILLER_9_766 ();
 sg13g2_decap_8 FILLER_9_773 ();
 sg13g2_decap_8 FILLER_9_780 ();
 sg13g2_decap_8 FILLER_9_787 ();
 sg13g2_decap_8 FILLER_9_794 ();
 sg13g2_decap_8 FILLER_9_801 ();
 sg13g2_decap_8 FILLER_9_808 ();
 sg13g2_decap_8 FILLER_9_815 ();
 sg13g2_decap_8 FILLER_9_822 ();
 sg13g2_decap_8 FILLER_9_829 ();
 sg13g2_decap_8 FILLER_9_836 ();
 sg13g2_decap_8 FILLER_9_843 ();
 sg13g2_decap_8 FILLER_9_850 ();
 sg13g2_decap_4 FILLER_9_857 ();
 sg13g2_fill_1 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_fill_2 FILLER_10_98 ();
 sg13g2_fill_1 FILLER_10_100 ();
 sg13g2_fill_2 FILLER_10_115 ();
 sg13g2_decap_8 FILLER_10_121 ();
 sg13g2_fill_2 FILLER_10_128 ();
 sg13g2_fill_1 FILLER_10_130 ();
 sg13g2_fill_2 FILLER_10_145 ();
 sg13g2_fill_1 FILLER_10_152 ();
 sg13g2_fill_2 FILLER_10_158 ();
 sg13g2_fill_1 FILLER_10_160 ();
 sg13g2_fill_1 FILLER_10_174 ();
 sg13g2_decap_8 FILLER_10_179 ();
 sg13g2_decap_8 FILLER_10_186 ();
 sg13g2_decap_8 FILLER_10_193 ();
 sg13g2_decap_8 FILLER_10_200 ();
 sg13g2_decap_8 FILLER_10_207 ();
 sg13g2_decap_8 FILLER_10_214 ();
 sg13g2_decap_8 FILLER_10_221 ();
 sg13g2_decap_8 FILLER_10_228 ();
 sg13g2_decap_8 FILLER_10_235 ();
 sg13g2_decap_8 FILLER_10_242 ();
 sg13g2_decap_8 FILLER_10_249 ();
 sg13g2_decap_8 FILLER_10_256 ();
 sg13g2_decap_8 FILLER_10_263 ();
 sg13g2_decap_8 FILLER_10_270 ();
 sg13g2_decap_8 FILLER_10_277 ();
 sg13g2_decap_8 FILLER_10_284 ();
 sg13g2_decap_8 FILLER_10_291 ();
 sg13g2_decap_8 FILLER_10_298 ();
 sg13g2_decap_8 FILLER_10_305 ();
 sg13g2_decap_8 FILLER_10_312 ();
 sg13g2_decap_8 FILLER_10_319 ();
 sg13g2_decap_8 FILLER_10_326 ();
 sg13g2_decap_8 FILLER_10_333 ();
 sg13g2_decap_8 FILLER_10_340 ();
 sg13g2_fill_2 FILLER_10_347 ();
 sg13g2_fill_1 FILLER_10_349 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_434 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_decap_4 FILLER_10_448 ();
 sg13g2_decap_4 FILLER_10_456 ();
 sg13g2_fill_2 FILLER_10_465 ();
 sg13g2_fill_1 FILLER_10_467 ();
 sg13g2_fill_2 FILLER_10_473 ();
 sg13g2_decap_8 FILLER_10_493 ();
 sg13g2_decap_8 FILLER_10_500 ();
 sg13g2_fill_1 FILLER_10_507 ();
 sg13g2_fill_1 FILLER_10_512 ();
 sg13g2_fill_2 FILLER_10_541 ();
 sg13g2_fill_1 FILLER_10_543 ();
 sg13g2_decap_8 FILLER_10_557 ();
 sg13g2_decap_8 FILLER_10_564 ();
 sg13g2_decap_8 FILLER_10_571 ();
 sg13g2_decap_8 FILLER_10_578 ();
 sg13g2_decap_8 FILLER_10_585 ();
 sg13g2_decap_8 FILLER_10_592 ();
 sg13g2_decap_8 FILLER_10_599 ();
 sg13g2_decap_8 FILLER_10_606 ();
 sg13g2_decap_8 FILLER_10_613 ();
 sg13g2_decap_8 FILLER_10_620 ();
 sg13g2_decap_8 FILLER_10_627 ();
 sg13g2_decap_8 FILLER_10_634 ();
 sg13g2_decap_8 FILLER_10_641 ();
 sg13g2_decap_8 FILLER_10_648 ();
 sg13g2_decap_8 FILLER_10_655 ();
 sg13g2_decap_8 FILLER_10_662 ();
 sg13g2_decap_8 FILLER_10_669 ();
 sg13g2_decap_8 FILLER_10_676 ();
 sg13g2_decap_8 FILLER_10_683 ();
 sg13g2_decap_8 FILLER_10_690 ();
 sg13g2_decap_8 FILLER_10_697 ();
 sg13g2_decap_8 FILLER_10_704 ();
 sg13g2_decap_8 FILLER_10_711 ();
 sg13g2_decap_8 FILLER_10_718 ();
 sg13g2_decap_8 FILLER_10_725 ();
 sg13g2_decap_8 FILLER_10_732 ();
 sg13g2_decap_8 FILLER_10_739 ();
 sg13g2_decap_8 FILLER_10_746 ();
 sg13g2_decap_8 FILLER_10_753 ();
 sg13g2_decap_8 FILLER_10_760 ();
 sg13g2_decap_8 FILLER_10_767 ();
 sg13g2_decap_8 FILLER_10_774 ();
 sg13g2_decap_8 FILLER_10_781 ();
 sg13g2_decap_8 FILLER_10_788 ();
 sg13g2_decap_8 FILLER_10_795 ();
 sg13g2_decap_8 FILLER_10_802 ();
 sg13g2_decap_8 FILLER_10_809 ();
 sg13g2_decap_8 FILLER_10_816 ();
 sg13g2_decap_8 FILLER_10_823 ();
 sg13g2_decap_8 FILLER_10_830 ();
 sg13g2_decap_8 FILLER_10_837 ();
 sg13g2_decap_8 FILLER_10_844 ();
 sg13g2_decap_8 FILLER_10_851 ();
 sg13g2_decap_4 FILLER_10_858 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_fill_2 FILLER_11_77 ();
 sg13g2_fill_1 FILLER_11_79 ();
 sg13g2_fill_2 FILLER_11_132 ();
 sg13g2_fill_1 FILLER_11_134 ();
 sg13g2_fill_2 FILLER_11_161 ();
 sg13g2_fill_1 FILLER_11_163 ();
 sg13g2_decap_8 FILLER_11_200 ();
 sg13g2_decap_8 FILLER_11_211 ();
 sg13g2_fill_1 FILLER_11_218 ();
 sg13g2_decap_8 FILLER_11_233 ();
 sg13g2_fill_2 FILLER_11_240 ();
 sg13g2_fill_1 FILLER_11_242 ();
 sg13g2_decap_4 FILLER_11_269 ();
 sg13g2_fill_2 FILLER_11_273 ();
 sg13g2_fill_2 FILLER_11_279 ();
 sg13g2_fill_1 FILLER_11_281 ();
 sg13g2_decap_8 FILLER_11_296 ();
 sg13g2_decap_8 FILLER_11_303 ();
 sg13g2_decap_8 FILLER_11_310 ();
 sg13g2_decap_8 FILLER_11_317 ();
 sg13g2_decap_8 FILLER_11_324 ();
 sg13g2_decap_8 FILLER_11_331 ();
 sg13g2_fill_2 FILLER_11_338 ();
 sg13g2_fill_2 FILLER_11_344 ();
 sg13g2_fill_2 FILLER_11_355 ();
 sg13g2_fill_2 FILLER_11_379 ();
 sg13g2_fill_1 FILLER_11_390 ();
 sg13g2_decap_8 FILLER_11_417 ();
 sg13g2_decap_8 FILLER_11_424 ();
 sg13g2_decap_8 FILLER_11_431 ();
 sg13g2_decap_4 FILLER_11_438 ();
 sg13g2_fill_2 FILLER_11_475 ();
 sg13g2_decap_8 FILLER_11_564 ();
 sg13g2_decap_8 FILLER_11_571 ();
 sg13g2_decap_8 FILLER_11_578 ();
 sg13g2_decap_8 FILLER_11_585 ();
 sg13g2_decap_8 FILLER_11_592 ();
 sg13g2_decap_8 FILLER_11_599 ();
 sg13g2_decap_8 FILLER_11_606 ();
 sg13g2_decap_8 FILLER_11_613 ();
 sg13g2_decap_8 FILLER_11_620 ();
 sg13g2_decap_8 FILLER_11_627 ();
 sg13g2_decap_8 FILLER_11_634 ();
 sg13g2_decap_8 FILLER_11_641 ();
 sg13g2_decap_8 FILLER_11_648 ();
 sg13g2_decap_8 FILLER_11_655 ();
 sg13g2_decap_8 FILLER_11_662 ();
 sg13g2_decap_8 FILLER_11_669 ();
 sg13g2_decap_8 FILLER_11_676 ();
 sg13g2_decap_8 FILLER_11_683 ();
 sg13g2_decap_8 FILLER_11_690 ();
 sg13g2_decap_8 FILLER_11_697 ();
 sg13g2_decap_8 FILLER_11_704 ();
 sg13g2_decap_8 FILLER_11_711 ();
 sg13g2_decap_8 FILLER_11_718 ();
 sg13g2_decap_8 FILLER_11_725 ();
 sg13g2_decap_8 FILLER_11_732 ();
 sg13g2_decap_8 FILLER_11_739 ();
 sg13g2_decap_8 FILLER_11_746 ();
 sg13g2_decap_8 FILLER_11_753 ();
 sg13g2_decap_8 FILLER_11_760 ();
 sg13g2_decap_8 FILLER_11_767 ();
 sg13g2_decap_8 FILLER_11_774 ();
 sg13g2_decap_8 FILLER_11_781 ();
 sg13g2_decap_8 FILLER_11_788 ();
 sg13g2_decap_8 FILLER_11_795 ();
 sg13g2_decap_8 FILLER_11_802 ();
 sg13g2_decap_8 FILLER_11_809 ();
 sg13g2_decap_8 FILLER_11_816 ();
 sg13g2_decap_8 FILLER_11_823 ();
 sg13g2_decap_8 FILLER_11_830 ();
 sg13g2_decap_8 FILLER_11_837 ();
 sg13g2_decap_8 FILLER_11_844 ();
 sg13g2_decap_8 FILLER_11_851 ();
 sg13g2_decap_4 FILLER_11_858 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_4 FILLER_12_56 ();
 sg13g2_fill_2 FILLER_12_60 ();
 sg13g2_fill_1 FILLER_12_88 ();
 sg13g2_decap_8 FILLER_12_107 ();
 sg13g2_decap_8 FILLER_12_114 ();
 sg13g2_fill_2 FILLER_12_147 ();
 sg13g2_fill_2 FILLER_12_184 ();
 sg13g2_fill_1 FILLER_12_247 ();
 sg13g2_decap_4 FILLER_12_257 ();
 sg13g2_decap_8 FILLER_12_313 ();
 sg13g2_decap_8 FILLER_12_320 ();
 sg13g2_fill_2 FILLER_12_327 ();
 sg13g2_fill_1 FILLER_12_329 ();
 sg13g2_decap_4 FILLER_12_356 ();
 sg13g2_fill_1 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_416 ();
 sg13g2_decap_8 FILLER_12_423 ();
 sg13g2_decap_4 FILLER_12_430 ();
 sg13g2_fill_2 FILLER_12_434 ();
 sg13g2_fill_1 FILLER_12_462 ();
 sg13g2_decap_8 FILLER_12_573 ();
 sg13g2_decap_8 FILLER_12_580 ();
 sg13g2_decap_8 FILLER_12_587 ();
 sg13g2_decap_8 FILLER_12_594 ();
 sg13g2_decap_8 FILLER_12_601 ();
 sg13g2_decap_8 FILLER_12_608 ();
 sg13g2_decap_8 FILLER_12_615 ();
 sg13g2_decap_8 FILLER_12_622 ();
 sg13g2_decap_8 FILLER_12_629 ();
 sg13g2_decap_8 FILLER_12_636 ();
 sg13g2_decap_8 FILLER_12_643 ();
 sg13g2_decap_8 FILLER_12_650 ();
 sg13g2_decap_8 FILLER_12_657 ();
 sg13g2_decap_8 FILLER_12_664 ();
 sg13g2_decap_8 FILLER_12_671 ();
 sg13g2_decap_8 FILLER_12_678 ();
 sg13g2_decap_8 FILLER_12_685 ();
 sg13g2_decap_8 FILLER_12_692 ();
 sg13g2_decap_8 FILLER_12_699 ();
 sg13g2_decap_8 FILLER_12_706 ();
 sg13g2_decap_8 FILLER_12_713 ();
 sg13g2_decap_8 FILLER_12_720 ();
 sg13g2_decap_8 FILLER_12_727 ();
 sg13g2_decap_8 FILLER_12_734 ();
 sg13g2_decap_8 FILLER_12_741 ();
 sg13g2_decap_8 FILLER_12_748 ();
 sg13g2_decap_8 FILLER_12_755 ();
 sg13g2_decap_8 FILLER_12_762 ();
 sg13g2_decap_8 FILLER_12_769 ();
 sg13g2_decap_8 FILLER_12_776 ();
 sg13g2_decap_8 FILLER_12_783 ();
 sg13g2_decap_8 FILLER_12_790 ();
 sg13g2_decap_8 FILLER_12_797 ();
 sg13g2_decap_8 FILLER_12_804 ();
 sg13g2_decap_8 FILLER_12_811 ();
 sg13g2_decap_8 FILLER_12_818 ();
 sg13g2_decap_8 FILLER_12_825 ();
 sg13g2_decap_8 FILLER_12_832 ();
 sg13g2_decap_8 FILLER_12_839 ();
 sg13g2_decap_8 FILLER_12_846 ();
 sg13g2_decap_8 FILLER_12_853 ();
 sg13g2_fill_2 FILLER_12_860 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_fill_2 FILLER_13_70 ();
 sg13g2_fill_1 FILLER_13_72 ();
 sg13g2_decap_4 FILLER_13_77 ();
 sg13g2_decap_4 FILLER_13_86 ();
 sg13g2_fill_2 FILLER_13_121 ();
 sg13g2_fill_1 FILLER_13_123 ();
 sg13g2_fill_2 FILLER_13_129 ();
 sg13g2_fill_1 FILLER_13_131 ();
 sg13g2_decap_8 FILLER_13_136 ();
 sg13g2_fill_1 FILLER_13_143 ();
 sg13g2_fill_1 FILLER_13_153 ();
 sg13g2_fill_2 FILLER_13_163 ();
 sg13g2_fill_1 FILLER_13_165 ();
 sg13g2_fill_2 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_208 ();
 sg13g2_decap_8 FILLER_13_215 ();
 sg13g2_fill_1 FILLER_13_222 ();
 sg13g2_fill_2 FILLER_13_231 ();
 sg13g2_decap_4 FILLER_13_242 ();
 sg13g2_fill_1 FILLER_13_246 ();
 sg13g2_fill_2 FILLER_13_252 ();
 sg13g2_decap_4 FILLER_13_258 ();
 sg13g2_fill_2 FILLER_13_276 ();
 sg13g2_fill_1 FILLER_13_278 ();
 sg13g2_fill_2 FILLER_13_319 ();
 sg13g2_fill_1 FILLER_13_354 ();
 sg13g2_decap_4 FILLER_13_424 ();
 sg13g2_fill_1 FILLER_13_428 ();
 sg13g2_fill_1 FILLER_13_455 ();
 sg13g2_fill_1 FILLER_13_464 ();
 sg13g2_fill_2 FILLER_13_500 ();
 sg13g2_fill_1 FILLER_13_502 ();
 sg13g2_fill_1 FILLER_13_560 ();
 sg13g2_decap_8 FILLER_13_587 ();
 sg13g2_decap_8 FILLER_13_594 ();
 sg13g2_decap_8 FILLER_13_601 ();
 sg13g2_decap_8 FILLER_13_608 ();
 sg13g2_fill_2 FILLER_13_615 ();
 sg13g2_decap_8 FILLER_13_625 ();
 sg13g2_decap_8 FILLER_13_632 ();
 sg13g2_decap_8 FILLER_13_639 ();
 sg13g2_decap_8 FILLER_13_646 ();
 sg13g2_decap_8 FILLER_13_653 ();
 sg13g2_decap_8 FILLER_13_660 ();
 sg13g2_decap_8 FILLER_13_667 ();
 sg13g2_decap_8 FILLER_13_674 ();
 sg13g2_decap_8 FILLER_13_681 ();
 sg13g2_decap_8 FILLER_13_688 ();
 sg13g2_decap_8 FILLER_13_695 ();
 sg13g2_decap_8 FILLER_13_702 ();
 sg13g2_decap_8 FILLER_13_709 ();
 sg13g2_decap_8 FILLER_13_716 ();
 sg13g2_decap_8 FILLER_13_723 ();
 sg13g2_decap_8 FILLER_13_730 ();
 sg13g2_decap_8 FILLER_13_737 ();
 sg13g2_decap_8 FILLER_13_744 ();
 sg13g2_decap_8 FILLER_13_751 ();
 sg13g2_decap_8 FILLER_13_758 ();
 sg13g2_decap_8 FILLER_13_765 ();
 sg13g2_decap_8 FILLER_13_772 ();
 sg13g2_decap_8 FILLER_13_779 ();
 sg13g2_decap_8 FILLER_13_786 ();
 sg13g2_decap_8 FILLER_13_793 ();
 sg13g2_decap_8 FILLER_13_800 ();
 sg13g2_decap_8 FILLER_13_807 ();
 sg13g2_decap_8 FILLER_13_814 ();
 sg13g2_decap_8 FILLER_13_821 ();
 sg13g2_decap_8 FILLER_13_828 ();
 sg13g2_decap_8 FILLER_13_835 ();
 sg13g2_decap_8 FILLER_13_842 ();
 sg13g2_decap_8 FILLER_13_849 ();
 sg13g2_decap_4 FILLER_13_856 ();
 sg13g2_fill_2 FILLER_13_860 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_fill_2 FILLER_14_70 ();
 sg13g2_fill_2 FILLER_14_85 ();
 sg13g2_fill_2 FILLER_14_101 ();
 sg13g2_fill_1 FILLER_14_103 ();
 sg13g2_fill_1 FILLER_14_174 ();
 sg13g2_fill_2 FILLER_14_179 ();
 sg13g2_fill_1 FILLER_14_181 ();
 sg13g2_fill_2 FILLER_14_191 ();
 sg13g2_decap_8 FILLER_14_197 ();
 sg13g2_decap_4 FILLER_14_230 ();
 sg13g2_decap_4 FILLER_14_239 ();
 sg13g2_decap_8 FILLER_14_251 ();
 sg13g2_decap_4 FILLER_14_258 ();
 sg13g2_fill_2 FILLER_14_262 ();
 sg13g2_fill_2 FILLER_14_269 ();
 sg13g2_fill_1 FILLER_14_302 ();
 sg13g2_decap_4 FILLER_14_307 ();
 sg13g2_fill_2 FILLER_14_311 ();
 sg13g2_decap_4 FILLER_14_318 ();
 sg13g2_fill_2 FILLER_14_322 ();
 sg13g2_fill_2 FILLER_14_329 ();
 sg13g2_fill_1 FILLER_14_331 ();
 sg13g2_decap_4 FILLER_14_336 ();
 sg13g2_fill_1 FILLER_14_349 ();
 sg13g2_decap_8 FILLER_14_382 ();
 sg13g2_decap_4 FILLER_14_389 ();
 sg13g2_decap_8 FILLER_14_402 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_fill_2 FILLER_14_420 ();
 sg13g2_fill_1 FILLER_14_422 ();
 sg13g2_fill_2 FILLER_14_520 ();
 sg13g2_fill_2 FILLER_14_531 ();
 sg13g2_decap_4 FILLER_14_593 ();
 sg13g2_fill_1 FILLER_14_597 ();
 sg13g2_fill_2 FILLER_14_627 ();
 sg13g2_decap_8 FILLER_14_642 ();
 sg13g2_decap_8 FILLER_14_649 ();
 sg13g2_decap_8 FILLER_14_656 ();
 sg13g2_decap_8 FILLER_14_663 ();
 sg13g2_decap_8 FILLER_14_670 ();
 sg13g2_decap_8 FILLER_14_677 ();
 sg13g2_fill_1 FILLER_14_684 ();
 sg13g2_decap_8 FILLER_14_690 ();
 sg13g2_decap_8 FILLER_14_697 ();
 sg13g2_decap_8 FILLER_14_704 ();
 sg13g2_decap_8 FILLER_14_711 ();
 sg13g2_decap_8 FILLER_14_718 ();
 sg13g2_decap_8 FILLER_14_725 ();
 sg13g2_decap_8 FILLER_14_732 ();
 sg13g2_decap_8 FILLER_14_739 ();
 sg13g2_decap_8 FILLER_14_746 ();
 sg13g2_decap_8 FILLER_14_753 ();
 sg13g2_decap_8 FILLER_14_760 ();
 sg13g2_decap_8 FILLER_14_767 ();
 sg13g2_decap_8 FILLER_14_774 ();
 sg13g2_decap_8 FILLER_14_781 ();
 sg13g2_decap_8 FILLER_14_788 ();
 sg13g2_decap_8 FILLER_14_795 ();
 sg13g2_decap_8 FILLER_14_802 ();
 sg13g2_decap_8 FILLER_14_809 ();
 sg13g2_decap_8 FILLER_14_816 ();
 sg13g2_decap_8 FILLER_14_823 ();
 sg13g2_decap_8 FILLER_14_830 ();
 sg13g2_decap_8 FILLER_14_837 ();
 sg13g2_decap_8 FILLER_14_844 ();
 sg13g2_decap_8 FILLER_14_851 ();
 sg13g2_decap_4 FILLER_14_858 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_4 FILLER_15_56 ();
 sg13g2_fill_1 FILLER_15_127 ();
 sg13g2_decap_8 FILLER_15_132 ();
 sg13g2_fill_2 FILLER_15_139 ();
 sg13g2_fill_2 FILLER_15_162 ();
 sg13g2_decap_8 FILLER_15_220 ();
 sg13g2_decap_4 FILLER_15_227 ();
 sg13g2_fill_1 FILLER_15_257 ();
 sg13g2_decap_8 FILLER_15_345 ();
 sg13g2_fill_2 FILLER_15_352 ();
 sg13g2_fill_1 FILLER_15_358 ();
 sg13g2_decap_8 FILLER_15_419 ();
 sg13g2_decap_8 FILLER_15_426 ();
 sg13g2_fill_1 FILLER_15_433 ();
 sg13g2_fill_1 FILLER_15_438 ();
 sg13g2_fill_2 FILLER_15_498 ();
 sg13g2_fill_2 FILLER_15_588 ();
 sg13g2_fill_1 FILLER_15_590 ();
 sg13g2_decap_8 FILLER_15_647 ();
 sg13g2_decap_8 FILLER_15_654 ();
 sg13g2_decap_8 FILLER_15_661 ();
 sg13g2_fill_2 FILLER_15_677 ();
 sg13g2_fill_1 FILLER_15_679 ();
 sg13g2_fill_2 FILLER_15_685 ();
 sg13g2_fill_2 FILLER_15_700 ();
 sg13g2_fill_1 FILLER_15_702 ();
 sg13g2_decap_8 FILLER_15_712 ();
 sg13g2_decap_8 FILLER_15_719 ();
 sg13g2_decap_8 FILLER_15_726 ();
 sg13g2_decap_8 FILLER_15_733 ();
 sg13g2_decap_8 FILLER_15_740 ();
 sg13g2_decap_8 FILLER_15_747 ();
 sg13g2_decap_8 FILLER_15_754 ();
 sg13g2_decap_8 FILLER_15_761 ();
 sg13g2_decap_8 FILLER_15_768 ();
 sg13g2_decap_8 FILLER_15_775 ();
 sg13g2_decap_8 FILLER_15_782 ();
 sg13g2_decap_8 FILLER_15_789 ();
 sg13g2_decap_8 FILLER_15_796 ();
 sg13g2_decap_8 FILLER_15_803 ();
 sg13g2_decap_8 FILLER_15_810 ();
 sg13g2_decap_8 FILLER_15_817 ();
 sg13g2_decap_8 FILLER_15_824 ();
 sg13g2_decap_8 FILLER_15_831 ();
 sg13g2_decap_8 FILLER_15_838 ();
 sg13g2_decap_8 FILLER_15_845 ();
 sg13g2_decap_8 FILLER_15_852 ();
 sg13g2_fill_2 FILLER_15_859 ();
 sg13g2_fill_1 FILLER_15_861 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_4 FILLER_16_63 ();
 sg13g2_fill_1 FILLER_16_67 ();
 sg13g2_fill_1 FILLER_16_81 ();
 sg13g2_decap_8 FILLER_16_87 ();
 sg13g2_decap_8 FILLER_16_94 ();
 sg13g2_decap_4 FILLER_16_101 ();
 sg13g2_fill_2 FILLER_16_105 ();
 sg13g2_fill_2 FILLER_16_151 ();
 sg13g2_fill_2 FILLER_16_167 ();
 sg13g2_fill_1 FILLER_16_169 ();
 sg13g2_fill_2 FILLER_16_184 ();
 sg13g2_fill_1 FILLER_16_186 ();
 sg13g2_decap_8 FILLER_16_226 ();
 sg13g2_fill_2 FILLER_16_233 ();
 sg13g2_fill_1 FILLER_16_235 ();
 sg13g2_decap_8 FILLER_16_254 ();
 sg13g2_decap_8 FILLER_16_261 ();
 sg13g2_decap_8 FILLER_16_268 ();
 sg13g2_fill_2 FILLER_16_275 ();
 sg13g2_fill_1 FILLER_16_277 ();
 sg13g2_fill_2 FILLER_16_282 ();
 sg13g2_fill_1 FILLER_16_284 ();
 sg13g2_fill_1 FILLER_16_293 ();
 sg13g2_fill_1 FILLER_16_328 ();
 sg13g2_fill_1 FILLER_16_392 ();
 sg13g2_fill_1 FILLER_16_426 ();
 sg13g2_decap_8 FILLER_16_431 ();
 sg13g2_fill_2 FILLER_16_438 ();
 sg13g2_fill_1 FILLER_16_440 ();
 sg13g2_decap_4 FILLER_16_497 ();
 sg13g2_fill_1 FILLER_16_501 ();
 sg13g2_fill_2 FILLER_16_625 ();
 sg13g2_fill_1 FILLER_16_680 ();
 sg13g2_decap_8 FILLER_16_716 ();
 sg13g2_decap_8 FILLER_16_723 ();
 sg13g2_decap_8 FILLER_16_730 ();
 sg13g2_decap_8 FILLER_16_737 ();
 sg13g2_decap_8 FILLER_16_744 ();
 sg13g2_decap_8 FILLER_16_751 ();
 sg13g2_decap_8 FILLER_16_758 ();
 sg13g2_decap_8 FILLER_16_765 ();
 sg13g2_decap_8 FILLER_16_772 ();
 sg13g2_decap_8 FILLER_16_779 ();
 sg13g2_decap_8 FILLER_16_786 ();
 sg13g2_decap_8 FILLER_16_793 ();
 sg13g2_decap_8 FILLER_16_800 ();
 sg13g2_decap_8 FILLER_16_807 ();
 sg13g2_decap_8 FILLER_16_814 ();
 sg13g2_decap_8 FILLER_16_821 ();
 sg13g2_decap_8 FILLER_16_828 ();
 sg13g2_decap_8 FILLER_16_835 ();
 sg13g2_decap_8 FILLER_16_842 ();
 sg13g2_decap_8 FILLER_16_849 ();
 sg13g2_decap_4 FILLER_16_856 ();
 sg13g2_fill_2 FILLER_16_860 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_4 FILLER_17_56 ();
 sg13g2_decap_4 FILLER_17_90 ();
 sg13g2_fill_2 FILLER_17_94 ();
 sg13g2_decap_4 FILLER_17_100 ();
 sg13g2_fill_2 FILLER_17_117 ();
 sg13g2_fill_1 FILLER_17_119 ();
 sg13g2_fill_2 FILLER_17_147 ();
 sg13g2_fill_1 FILLER_17_149 ();
 sg13g2_fill_2 FILLER_17_159 ();
 sg13g2_fill_1 FILLER_17_161 ();
 sg13g2_fill_2 FILLER_17_193 ();
 sg13g2_fill_1 FILLER_17_195 ();
 sg13g2_decap_8 FILLER_17_201 ();
 sg13g2_decap_8 FILLER_17_234 ();
 sg13g2_fill_1 FILLER_17_241 ();
 sg13g2_fill_1 FILLER_17_308 ();
 sg13g2_fill_1 FILLER_17_363 ();
 sg13g2_fill_2 FILLER_17_413 ();
 sg13g2_fill_1 FILLER_17_415 ();
 sg13g2_decap_8 FILLER_17_442 ();
 sg13g2_fill_2 FILLER_17_449 ();
 sg13g2_fill_1 FILLER_17_451 ();
 sg13g2_fill_2 FILLER_17_456 ();
 sg13g2_fill_1 FILLER_17_458 ();
 sg13g2_fill_2 FILLER_17_473 ();
 sg13g2_fill_2 FILLER_17_501 ();
 sg13g2_fill_1 FILLER_17_503 ();
 sg13g2_decap_4 FILLER_17_527 ();
 sg13g2_fill_1 FILLER_17_531 ();
 sg13g2_fill_1 FILLER_17_553 ();
 sg13g2_fill_2 FILLER_17_594 ();
 sg13g2_fill_1 FILLER_17_606 ();
 sg13g2_fill_1 FILLER_17_616 ();
 sg13g2_decap_4 FILLER_17_657 ();
 sg13g2_fill_1 FILLER_17_661 ();
 sg13g2_fill_1 FILLER_17_671 ();
 sg13g2_fill_2 FILLER_17_677 ();
 sg13g2_fill_2 FILLER_17_688 ();
 sg13g2_fill_1 FILLER_17_690 ();
 sg13g2_fill_2 FILLER_17_696 ();
 sg13g2_fill_1 FILLER_17_698 ();
 sg13g2_decap_8 FILLER_17_725 ();
 sg13g2_decap_8 FILLER_17_732 ();
 sg13g2_decap_8 FILLER_17_739 ();
 sg13g2_decap_8 FILLER_17_746 ();
 sg13g2_decap_8 FILLER_17_753 ();
 sg13g2_decap_8 FILLER_17_760 ();
 sg13g2_decap_8 FILLER_17_767 ();
 sg13g2_decap_8 FILLER_17_774 ();
 sg13g2_decap_8 FILLER_17_781 ();
 sg13g2_decap_8 FILLER_17_788 ();
 sg13g2_decap_8 FILLER_17_795 ();
 sg13g2_decap_8 FILLER_17_802 ();
 sg13g2_decap_8 FILLER_17_809 ();
 sg13g2_decap_8 FILLER_17_816 ();
 sg13g2_decap_8 FILLER_17_823 ();
 sg13g2_decap_8 FILLER_17_830 ();
 sg13g2_decap_8 FILLER_17_837 ();
 sg13g2_decap_8 FILLER_17_844 ();
 sg13g2_decap_8 FILLER_17_851 ();
 sg13g2_decap_4 FILLER_17_858 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_4 FILLER_18_63 ();
 sg13g2_fill_1 FILLER_18_67 ();
 sg13g2_fill_2 FILLER_18_129 ();
 sg13g2_fill_2 FILLER_18_172 ();
 sg13g2_fill_1 FILLER_18_177 ();
 sg13g2_decap_4 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_214 ();
 sg13g2_fill_1 FILLER_18_221 ();
 sg13g2_decap_8 FILLER_18_226 ();
 sg13g2_decap_8 FILLER_18_233 ();
 sg13g2_decap_8 FILLER_18_240 ();
 sg13g2_decap_8 FILLER_18_247 ();
 sg13g2_decap_4 FILLER_18_254 ();
 sg13g2_fill_2 FILLER_18_258 ();
 sg13g2_fill_1 FILLER_18_264 ();
 sg13g2_fill_1 FILLER_18_324 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_fill_2 FILLER_18_344 ();
 sg13g2_fill_2 FILLER_18_365 ();
 sg13g2_fill_2 FILLER_18_377 ();
 sg13g2_decap_4 FILLER_18_437 ();
 sg13g2_decap_4 FILLER_18_476 ();
 sg13g2_fill_2 FILLER_18_480 ();
 sg13g2_decap_4 FILLER_18_490 ();
 sg13g2_fill_2 FILLER_18_530 ();
 sg13g2_fill_1 FILLER_18_532 ();
 sg13g2_fill_1 FILLER_18_574 ();
 sg13g2_fill_1 FILLER_18_601 ();
 sg13g2_fill_2 FILLER_18_641 ();
 sg13g2_fill_1 FILLER_18_643 ();
 sg13g2_fill_2 FILLER_18_691 ();
 sg13g2_decap_8 FILLER_18_724 ();
 sg13g2_decap_8 FILLER_18_731 ();
 sg13g2_decap_8 FILLER_18_738 ();
 sg13g2_decap_8 FILLER_18_745 ();
 sg13g2_decap_8 FILLER_18_752 ();
 sg13g2_decap_8 FILLER_18_759 ();
 sg13g2_decap_8 FILLER_18_766 ();
 sg13g2_decap_8 FILLER_18_773 ();
 sg13g2_decap_8 FILLER_18_780 ();
 sg13g2_decap_8 FILLER_18_787 ();
 sg13g2_decap_8 FILLER_18_794 ();
 sg13g2_decap_8 FILLER_18_801 ();
 sg13g2_decap_8 FILLER_18_808 ();
 sg13g2_decap_8 FILLER_18_815 ();
 sg13g2_decap_8 FILLER_18_822 ();
 sg13g2_decap_8 FILLER_18_829 ();
 sg13g2_decap_8 FILLER_18_836 ();
 sg13g2_decap_8 FILLER_18_843 ();
 sg13g2_decap_8 FILLER_18_850 ();
 sg13g2_decap_4 FILLER_18_857 ();
 sg13g2_fill_1 FILLER_18_861 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_4 FILLER_19_77 ();
 sg13g2_fill_2 FILLER_19_81 ();
 sg13g2_fill_1 FILLER_19_97 ();
 sg13g2_fill_2 FILLER_19_105 ();
 sg13g2_decap_4 FILLER_19_111 ();
 sg13g2_decap_4 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_138 ();
 sg13g2_fill_2 FILLER_19_145 ();
 sg13g2_fill_1 FILLER_19_147 ();
 sg13g2_fill_2 FILLER_19_165 ();
 sg13g2_decap_4 FILLER_19_193 ();
 sg13g2_fill_1 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_237 ();
 sg13g2_decap_8 FILLER_19_244 ();
 sg13g2_decap_8 FILLER_19_251 ();
 sg13g2_fill_2 FILLER_19_258 ();
 sg13g2_fill_2 FILLER_19_291 ();
 sg13g2_fill_1 FILLER_19_303 ();
 sg13g2_decap_4 FILLER_19_325 ();
 sg13g2_fill_1 FILLER_19_336 ();
 sg13g2_decap_4 FILLER_19_341 ();
 sg13g2_fill_1 FILLER_19_345 ();
 sg13g2_fill_1 FILLER_19_362 ();
 sg13g2_decap_4 FILLER_19_427 ();
 sg13g2_decap_8 FILLER_19_477 ();
 sg13g2_fill_2 FILLER_19_507 ();
 sg13g2_decap_8 FILLER_19_535 ();
 sg13g2_fill_2 FILLER_19_542 ();
 sg13g2_fill_1 FILLER_19_553 ();
 sg13g2_fill_1 FILLER_19_558 ();
 sg13g2_decap_4 FILLER_19_564 ();
 sg13g2_fill_1 FILLER_19_598 ();
 sg13g2_fill_2 FILLER_19_635 ();
 sg13g2_fill_2 FILLER_19_679 ();
 sg13g2_fill_2 FILLER_19_699 ();
 sg13g2_fill_1 FILLER_19_701 ();
 sg13g2_decap_8 FILLER_19_728 ();
 sg13g2_decap_8 FILLER_19_735 ();
 sg13g2_decap_8 FILLER_19_742 ();
 sg13g2_decap_8 FILLER_19_749 ();
 sg13g2_decap_8 FILLER_19_756 ();
 sg13g2_decap_8 FILLER_19_763 ();
 sg13g2_decap_8 FILLER_19_770 ();
 sg13g2_decap_8 FILLER_19_777 ();
 sg13g2_decap_8 FILLER_19_784 ();
 sg13g2_decap_8 FILLER_19_791 ();
 sg13g2_decap_8 FILLER_19_798 ();
 sg13g2_decap_8 FILLER_19_805 ();
 sg13g2_decap_8 FILLER_19_812 ();
 sg13g2_decap_8 FILLER_19_819 ();
 sg13g2_decap_8 FILLER_19_826 ();
 sg13g2_decap_8 FILLER_19_833 ();
 sg13g2_decap_8 FILLER_19_840 ();
 sg13g2_decap_8 FILLER_19_847 ();
 sg13g2_decap_8 FILLER_19_854 ();
 sg13g2_fill_1 FILLER_19_861 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_fill_2 FILLER_20_70 ();
 sg13g2_fill_1 FILLER_20_72 ();
 sg13g2_fill_1 FILLER_20_107 ();
 sg13g2_fill_2 FILLER_20_138 ();
 sg13g2_fill_1 FILLER_20_246 ();
 sg13g2_fill_2 FILLER_20_273 ();
 sg13g2_fill_2 FILLER_20_302 ();
 sg13g2_fill_2 FILLER_20_324 ();
 sg13g2_fill_1 FILLER_20_359 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_fill_1 FILLER_20_418 ();
 sg13g2_fill_2 FILLER_20_448 ();
 sg13g2_decap_8 FILLER_20_467 ();
 sg13g2_fill_2 FILLER_20_474 ();
 sg13g2_decap_8 FILLER_20_513 ();
 sg13g2_fill_2 FILLER_20_536 ();
 sg13g2_fill_1 FILLER_20_538 ();
 sg13g2_decap_8 FILLER_20_543 ();
 sg13g2_decap_8 FILLER_20_550 ();
 sg13g2_fill_2 FILLER_20_557 ();
 sg13g2_fill_1 FILLER_20_559 ();
 sg13g2_decap_8 FILLER_20_564 ();
 sg13g2_fill_1 FILLER_20_571 ();
 sg13g2_fill_2 FILLER_20_623 ();
 sg13g2_fill_1 FILLER_20_625 ();
 sg13g2_decap_4 FILLER_20_652 ();
 sg13g2_fill_1 FILLER_20_693 ();
 sg13g2_fill_2 FILLER_20_703 ();
 sg13g2_decap_8 FILLER_20_727 ();
 sg13g2_decap_8 FILLER_20_734 ();
 sg13g2_decap_8 FILLER_20_741 ();
 sg13g2_decap_8 FILLER_20_748 ();
 sg13g2_decap_8 FILLER_20_755 ();
 sg13g2_decap_8 FILLER_20_762 ();
 sg13g2_decap_8 FILLER_20_769 ();
 sg13g2_decap_8 FILLER_20_776 ();
 sg13g2_decap_8 FILLER_20_783 ();
 sg13g2_decap_8 FILLER_20_790 ();
 sg13g2_decap_8 FILLER_20_797 ();
 sg13g2_decap_8 FILLER_20_804 ();
 sg13g2_decap_8 FILLER_20_811 ();
 sg13g2_decap_8 FILLER_20_818 ();
 sg13g2_decap_8 FILLER_20_825 ();
 sg13g2_decap_8 FILLER_20_832 ();
 sg13g2_decap_8 FILLER_20_839 ();
 sg13g2_decap_8 FILLER_20_846 ();
 sg13g2_decap_8 FILLER_20_853 ();
 sg13g2_fill_2 FILLER_20_860 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_fill_2 FILLER_21_70 ();
 sg13g2_fill_2 FILLER_21_95 ();
 sg13g2_fill_1 FILLER_21_97 ();
 sg13g2_fill_2 FILLER_21_125 ();
 sg13g2_fill_1 FILLER_21_141 ();
 sg13g2_decap_4 FILLER_21_152 ();
 sg13g2_fill_1 FILLER_21_156 ();
 sg13g2_fill_2 FILLER_21_171 ();
 sg13g2_fill_2 FILLER_21_236 ();
 sg13g2_decap_8 FILLER_21_246 ();
 sg13g2_decap_4 FILLER_21_253 ();
 sg13g2_decap_4 FILLER_21_261 ();
 sg13g2_fill_2 FILLER_21_288 ();
 sg13g2_fill_1 FILLER_21_290 ();
 sg13g2_decap_8 FILLER_21_317 ();
 sg13g2_decap_8 FILLER_21_324 ();
 sg13g2_fill_2 FILLER_21_331 ();
 sg13g2_fill_2 FILLER_21_372 ();
 sg13g2_fill_1 FILLER_21_374 ();
 sg13g2_decap_4 FILLER_21_380 ();
 sg13g2_fill_2 FILLER_21_384 ();
 sg13g2_fill_2 FILLER_21_453 ();
 sg13g2_decap_8 FILLER_21_481 ();
 sg13g2_fill_2 FILLER_21_488 ();
 sg13g2_fill_1 FILLER_21_490 ();
 sg13g2_fill_2 FILLER_21_595 ();
 sg13g2_decap_8 FILLER_21_612 ();
 sg13g2_fill_1 FILLER_21_619 ();
 sg13g2_fill_1 FILLER_21_625 ();
 sg13g2_decap_8 FILLER_21_631 ();
 sg13g2_fill_1 FILLER_21_638 ();
 sg13g2_decap_4 FILLER_21_652 ();
 sg13g2_fill_1 FILLER_21_656 ();
 sg13g2_fill_1 FILLER_21_671 ();
 sg13g2_fill_2 FILLER_21_681 ();
 sg13g2_fill_1 FILLER_21_683 ();
 sg13g2_decap_8 FILLER_21_719 ();
 sg13g2_decap_8 FILLER_21_726 ();
 sg13g2_decap_8 FILLER_21_733 ();
 sg13g2_decap_8 FILLER_21_740 ();
 sg13g2_decap_8 FILLER_21_747 ();
 sg13g2_decap_8 FILLER_21_754 ();
 sg13g2_decap_8 FILLER_21_761 ();
 sg13g2_decap_8 FILLER_21_768 ();
 sg13g2_decap_8 FILLER_21_775 ();
 sg13g2_decap_8 FILLER_21_782 ();
 sg13g2_decap_8 FILLER_21_789 ();
 sg13g2_decap_8 FILLER_21_796 ();
 sg13g2_decap_8 FILLER_21_803 ();
 sg13g2_decap_8 FILLER_21_810 ();
 sg13g2_decap_8 FILLER_21_817 ();
 sg13g2_decap_8 FILLER_21_824 ();
 sg13g2_decap_8 FILLER_21_831 ();
 sg13g2_decap_8 FILLER_21_838 ();
 sg13g2_decap_8 FILLER_21_845 ();
 sg13g2_decap_8 FILLER_21_852 ();
 sg13g2_fill_2 FILLER_21_859 ();
 sg13g2_fill_1 FILLER_21_861 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_fill_1 FILLER_22_94 ();
 sg13g2_fill_2 FILLER_22_104 ();
 sg13g2_fill_1 FILLER_22_117 ();
 sg13g2_fill_2 FILLER_22_128 ();
 sg13g2_fill_1 FILLER_22_130 ();
 sg13g2_fill_2 FILLER_22_174 ();
 sg13g2_fill_1 FILLER_22_176 ();
 sg13g2_fill_2 FILLER_22_200 ();
 sg13g2_fill_1 FILLER_22_202 ();
 sg13g2_fill_1 FILLER_22_275 ();
 sg13g2_fill_1 FILLER_22_299 ();
 sg13g2_decap_8 FILLER_22_310 ();
 sg13g2_decap_4 FILLER_22_317 ();
 sg13g2_fill_1 FILLER_22_325 ();
 sg13g2_decap_4 FILLER_22_352 ();
 sg13g2_fill_1 FILLER_22_356 ();
 sg13g2_decap_8 FILLER_22_366 ();
 sg13g2_decap_4 FILLER_22_373 ();
 sg13g2_fill_1 FILLER_22_377 ();
 sg13g2_fill_2 FILLER_22_391 ();
 sg13g2_decap_8 FILLER_22_456 ();
 sg13g2_fill_2 FILLER_22_463 ();
 sg13g2_fill_1 FILLER_22_465 ();
 sg13g2_decap_8 FILLER_22_470 ();
 sg13g2_decap_8 FILLER_22_481 ();
 sg13g2_decap_8 FILLER_22_488 ();
 sg13g2_decap_4 FILLER_22_495 ();
 sg13g2_fill_2 FILLER_22_595 ();
 sg13g2_fill_1 FILLER_22_597 ();
 sg13g2_fill_2 FILLER_22_610 ();
 sg13g2_decap_8 FILLER_22_642 ();
 sg13g2_fill_2 FILLER_22_687 ();
 sg13g2_fill_1 FILLER_22_689 ();
 sg13g2_fill_1 FILLER_22_703 ();
 sg13g2_decap_8 FILLER_22_708 ();
 sg13g2_decap_8 FILLER_22_715 ();
 sg13g2_decap_8 FILLER_22_722 ();
 sg13g2_decap_8 FILLER_22_729 ();
 sg13g2_decap_8 FILLER_22_736 ();
 sg13g2_decap_8 FILLER_22_743 ();
 sg13g2_decap_8 FILLER_22_750 ();
 sg13g2_decap_8 FILLER_22_757 ();
 sg13g2_decap_8 FILLER_22_764 ();
 sg13g2_decap_8 FILLER_22_771 ();
 sg13g2_decap_8 FILLER_22_778 ();
 sg13g2_decap_8 FILLER_22_785 ();
 sg13g2_decap_8 FILLER_22_792 ();
 sg13g2_decap_8 FILLER_22_799 ();
 sg13g2_decap_8 FILLER_22_806 ();
 sg13g2_decap_8 FILLER_22_813 ();
 sg13g2_decap_8 FILLER_22_820 ();
 sg13g2_decap_8 FILLER_22_827 ();
 sg13g2_decap_8 FILLER_22_834 ();
 sg13g2_decap_8 FILLER_22_841 ();
 sg13g2_decap_8 FILLER_22_848 ();
 sg13g2_decap_8 FILLER_22_855 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_fill_2 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_fill_1 FILLER_23_49 ();
 sg13g2_fill_2 FILLER_23_58 ();
 sg13g2_fill_1 FILLER_23_60 ();
 sg13g2_fill_2 FILLER_23_69 ();
 sg13g2_fill_1 FILLER_23_71 ();
 sg13g2_fill_2 FILLER_23_76 ();
 sg13g2_fill_1 FILLER_23_78 ();
 sg13g2_fill_1 FILLER_23_88 ();
 sg13g2_fill_2 FILLER_23_104 ();
 sg13g2_fill_1 FILLER_23_106 ();
 sg13g2_fill_1 FILLER_23_112 ();
 sg13g2_fill_2 FILLER_23_118 ();
 sg13g2_fill_1 FILLER_23_129 ();
 sg13g2_fill_2 FILLER_23_153 ();
 sg13g2_decap_8 FILLER_23_160 ();
 sg13g2_decap_4 FILLER_23_167 ();
 sg13g2_decap_4 FILLER_23_179 ();
 sg13g2_fill_1 FILLER_23_183 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_fill_1 FILLER_23_218 ();
 sg13g2_fill_2 FILLER_23_232 ();
 sg13g2_decap_8 FILLER_23_247 ();
 sg13g2_decap_4 FILLER_23_254 ();
 sg13g2_fill_2 FILLER_23_258 ();
 sg13g2_decap_8 FILLER_23_264 ();
 sg13g2_fill_1 FILLER_23_271 ();
 sg13g2_fill_2 FILLER_23_283 ();
 sg13g2_fill_2 FILLER_23_321 ();
 sg13g2_fill_1 FILLER_23_345 ();
 sg13g2_fill_1 FILLER_23_410 ();
 sg13g2_fill_2 FILLER_23_437 ();
 sg13g2_fill_1 FILLER_23_439 ();
 sg13g2_decap_8 FILLER_23_458 ();
 sg13g2_fill_1 FILLER_23_465 ();
 sg13g2_fill_1 FILLER_23_515 ();
 sg13g2_fill_1 FILLER_23_529 ();
 sg13g2_fill_1 FILLER_23_587 ();
 sg13g2_decap_4 FILLER_23_613 ();
 sg13g2_fill_2 FILLER_23_617 ();
 sg13g2_fill_1 FILLER_23_627 ();
 sg13g2_decap_4 FILLER_23_701 ();
 sg13g2_fill_2 FILLER_23_705 ();
 sg13g2_decap_8 FILLER_23_726 ();
 sg13g2_decap_8 FILLER_23_733 ();
 sg13g2_decap_8 FILLER_23_740 ();
 sg13g2_decap_8 FILLER_23_747 ();
 sg13g2_decap_8 FILLER_23_754 ();
 sg13g2_decap_8 FILLER_23_761 ();
 sg13g2_decap_8 FILLER_23_768 ();
 sg13g2_decap_8 FILLER_23_775 ();
 sg13g2_decap_8 FILLER_23_782 ();
 sg13g2_decap_8 FILLER_23_789 ();
 sg13g2_decap_8 FILLER_23_796 ();
 sg13g2_decap_8 FILLER_23_803 ();
 sg13g2_decap_8 FILLER_23_810 ();
 sg13g2_decap_8 FILLER_23_817 ();
 sg13g2_decap_8 FILLER_23_824 ();
 sg13g2_decap_8 FILLER_23_831 ();
 sg13g2_decap_8 FILLER_23_838 ();
 sg13g2_decap_8 FILLER_23_845 ();
 sg13g2_decap_8 FILLER_23_852 ();
 sg13g2_fill_2 FILLER_23_859 ();
 sg13g2_fill_1 FILLER_23_861 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_4 FILLER_24_21 ();
 sg13g2_fill_1 FILLER_24_30 ();
 sg13g2_fill_1 FILLER_24_91 ();
 sg13g2_fill_2 FILLER_24_148 ();
 sg13g2_fill_1 FILLER_24_150 ();
 sg13g2_decap_8 FILLER_24_165 ();
 sg13g2_fill_2 FILLER_24_177 ();
 sg13g2_decap_8 FILLER_24_186 ();
 sg13g2_fill_2 FILLER_24_193 ();
 sg13g2_fill_1 FILLER_24_195 ();
 sg13g2_fill_2 FILLER_24_201 ();
 sg13g2_fill_1 FILLER_24_208 ();
 sg13g2_fill_1 FILLER_24_226 ();
 sg13g2_decap_4 FILLER_24_253 ();
 sg13g2_fill_1 FILLER_24_257 ();
 sg13g2_decap_4 FILLER_24_262 ();
 sg13g2_fill_2 FILLER_24_266 ();
 sg13g2_fill_2 FILLER_24_276 ();
 sg13g2_fill_1 FILLER_24_278 ();
 sg13g2_fill_2 FILLER_24_298 ();
 sg13g2_decap_8 FILLER_24_359 ();
 sg13g2_fill_2 FILLER_24_366 ();
 sg13g2_fill_1 FILLER_24_368 ();
 sg13g2_fill_2 FILLER_24_375 ();
 sg13g2_decap_8 FILLER_24_385 ();
 sg13g2_decap_8 FILLER_24_392 ();
 sg13g2_fill_2 FILLER_24_399 ();
 sg13g2_fill_1 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_410 ();
 sg13g2_fill_2 FILLER_24_455 ();
 sg13g2_fill_1 FILLER_24_457 ();
 sg13g2_fill_2 FILLER_24_484 ();
 sg13g2_fill_1 FILLER_24_486 ();
 sg13g2_fill_1 FILLER_24_496 ();
 sg13g2_fill_2 FILLER_24_503 ();
 sg13g2_fill_1 FILLER_24_517 ();
 sg13g2_fill_2 FILLER_24_674 ();
 sg13g2_fill_1 FILLER_24_676 ();
 sg13g2_fill_1 FILLER_24_713 ();
 sg13g2_decap_8 FILLER_24_736 ();
 sg13g2_decap_8 FILLER_24_743 ();
 sg13g2_decap_8 FILLER_24_750 ();
 sg13g2_decap_8 FILLER_24_757 ();
 sg13g2_decap_8 FILLER_24_764 ();
 sg13g2_decap_8 FILLER_24_771 ();
 sg13g2_decap_8 FILLER_24_778 ();
 sg13g2_decap_8 FILLER_24_785 ();
 sg13g2_decap_8 FILLER_24_792 ();
 sg13g2_decap_8 FILLER_24_799 ();
 sg13g2_decap_8 FILLER_24_806 ();
 sg13g2_decap_8 FILLER_24_813 ();
 sg13g2_decap_8 FILLER_24_820 ();
 sg13g2_decap_8 FILLER_24_827 ();
 sg13g2_decap_8 FILLER_24_834 ();
 sg13g2_decap_8 FILLER_24_841 ();
 sg13g2_decap_8 FILLER_24_848 ();
 sg13g2_decap_8 FILLER_24_855 ();
 sg13g2_fill_1 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_30 ();
 sg13g2_fill_2 FILLER_25_43 ();
 sg13g2_fill_1 FILLER_25_55 ();
 sg13g2_fill_2 FILLER_25_65 ();
 sg13g2_fill_2 FILLER_25_77 ();
 sg13g2_fill_2 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_116 ();
 sg13g2_decap_8 FILLER_25_123 ();
 sg13g2_fill_2 FILLER_25_130 ();
 sg13g2_fill_1 FILLER_25_163 ();
 sg13g2_fill_2 FILLER_25_207 ();
 sg13g2_fill_2 FILLER_25_273 ();
 sg13g2_fill_1 FILLER_25_283 ();
 sg13g2_fill_2 FILLER_25_330 ();
 sg13g2_fill_2 FILLER_25_345 ();
 sg13g2_fill_1 FILLER_25_347 ();
 sg13g2_fill_1 FILLER_25_369 ();
 sg13g2_fill_2 FILLER_25_383 ();
 sg13g2_fill_1 FILLER_25_385 ();
 sg13g2_fill_1 FILLER_25_390 ();
 sg13g2_fill_1 FILLER_25_410 ();
 sg13g2_fill_2 FILLER_25_435 ();
 sg13g2_fill_1 FILLER_25_437 ();
 sg13g2_fill_1 FILLER_25_517 ();
 sg13g2_fill_1 FILLER_25_575 ();
 sg13g2_fill_1 FILLER_25_579 ();
 sg13g2_decap_4 FILLER_25_584 ();
 sg13g2_fill_2 FILLER_25_588 ();
 sg13g2_fill_2 FILLER_25_607 ();
 sg13g2_decap_8 FILLER_25_613 ();
 sg13g2_fill_2 FILLER_25_620 ();
 sg13g2_fill_2 FILLER_25_648 ();
 sg13g2_fill_2 FILLER_25_691 ();
 sg13g2_decap_8 FILLER_25_749 ();
 sg13g2_decap_8 FILLER_25_756 ();
 sg13g2_decap_8 FILLER_25_763 ();
 sg13g2_decap_8 FILLER_25_770 ();
 sg13g2_decap_8 FILLER_25_777 ();
 sg13g2_decap_8 FILLER_25_784 ();
 sg13g2_decap_8 FILLER_25_791 ();
 sg13g2_decap_8 FILLER_25_798 ();
 sg13g2_decap_8 FILLER_25_805 ();
 sg13g2_decap_8 FILLER_25_812 ();
 sg13g2_decap_8 FILLER_25_819 ();
 sg13g2_decap_8 FILLER_25_826 ();
 sg13g2_decap_8 FILLER_25_833 ();
 sg13g2_decap_8 FILLER_25_840 ();
 sg13g2_decap_8 FILLER_25_847 ();
 sg13g2_decap_8 FILLER_25_854 ();
 sg13g2_fill_1 FILLER_25_861 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_4 FILLER_26_7 ();
 sg13g2_fill_1 FILLER_26_33 ();
 sg13g2_fill_1 FILLER_26_58 ();
 sg13g2_fill_1 FILLER_26_118 ();
 sg13g2_fill_1 FILLER_26_136 ();
 sg13g2_decap_8 FILLER_26_156 ();
 sg13g2_decap_8 FILLER_26_163 ();
 sg13g2_fill_2 FILLER_26_170 ();
 sg13g2_fill_2 FILLER_26_177 ();
 sg13g2_decap_8 FILLER_26_194 ();
 sg13g2_decap_8 FILLER_26_264 ();
 sg13g2_decap_8 FILLER_26_271 ();
 sg13g2_decap_8 FILLER_26_282 ();
 sg13g2_decap_4 FILLER_26_289 ();
 sg13g2_fill_1 FILLER_26_297 ();
 sg13g2_fill_1 FILLER_26_302 ();
 sg13g2_fill_2 FILLER_26_307 ();
 sg13g2_fill_1 FILLER_26_309 ();
 sg13g2_fill_2 FILLER_26_319 ();
 sg13g2_fill_1 FILLER_26_451 ();
 sg13g2_fill_2 FILLER_26_465 ();
 sg13g2_fill_1 FILLER_26_467 ();
 sg13g2_fill_2 FILLER_26_527 ();
 sg13g2_fill_1 FILLER_26_529 ();
 sg13g2_fill_1 FILLER_26_559 ();
 sg13g2_fill_2 FILLER_26_624 ();
 sg13g2_fill_2 FILLER_26_674 ();
 sg13g2_fill_1 FILLER_26_676 ();
 sg13g2_fill_2 FILLER_26_703 ();
 sg13g2_fill_1 FILLER_26_705 ();
 sg13g2_decap_8 FILLER_26_754 ();
 sg13g2_decap_8 FILLER_26_761 ();
 sg13g2_decap_8 FILLER_26_768 ();
 sg13g2_decap_8 FILLER_26_775 ();
 sg13g2_decap_8 FILLER_26_782 ();
 sg13g2_decap_8 FILLER_26_789 ();
 sg13g2_decap_8 FILLER_26_796 ();
 sg13g2_decap_8 FILLER_26_803 ();
 sg13g2_decap_8 FILLER_26_810 ();
 sg13g2_decap_8 FILLER_26_817 ();
 sg13g2_decap_8 FILLER_26_824 ();
 sg13g2_decap_8 FILLER_26_831 ();
 sg13g2_decap_8 FILLER_26_838 ();
 sg13g2_decap_8 FILLER_26_845 ();
 sg13g2_decap_8 FILLER_26_852 ();
 sg13g2_fill_2 FILLER_26_859 ();
 sg13g2_fill_1 FILLER_26_861 ();
 sg13g2_fill_2 FILLER_27_26 ();
 sg13g2_decap_8 FILLER_27_75 ();
 sg13g2_decap_4 FILLER_27_82 ();
 sg13g2_fill_1 FILLER_27_86 ();
 sg13g2_decap_4 FILLER_27_96 ();
 sg13g2_fill_1 FILLER_27_100 ();
 sg13g2_decap_4 FILLER_27_105 ();
 sg13g2_fill_1 FILLER_27_109 ();
 sg13g2_decap_4 FILLER_27_115 ();
 sg13g2_fill_2 FILLER_27_119 ();
 sg13g2_fill_2 FILLER_27_153 ();
 sg13g2_decap_4 FILLER_27_163 ();
 sg13g2_decap_4 FILLER_27_199 ();
 sg13g2_fill_1 FILLER_27_203 ();
 sg13g2_decap_4 FILLER_27_214 ();
 sg13g2_fill_2 FILLER_27_231 ();
 sg13g2_fill_1 FILLER_27_277 ();
 sg13g2_fill_1 FILLER_27_335 ();
 sg13g2_fill_2 FILLER_27_349 ();
 sg13g2_decap_8 FILLER_27_359 ();
 sg13g2_fill_2 FILLER_27_389 ();
 sg13g2_fill_2 FILLER_27_400 ();
 sg13g2_fill_1 FILLER_27_402 ();
 sg13g2_fill_2 FILLER_27_411 ();
 sg13g2_fill_1 FILLER_27_463 ();
 sg13g2_fill_2 FILLER_27_493 ();
 sg13g2_fill_2 FILLER_27_624 ();
 sg13g2_fill_1 FILLER_27_626 ();
 sg13g2_fill_1 FILLER_27_671 ();
 sg13g2_fill_2 FILLER_27_695 ();
 sg13g2_decap_8 FILLER_27_766 ();
 sg13g2_decap_8 FILLER_27_773 ();
 sg13g2_decap_8 FILLER_27_780 ();
 sg13g2_decap_8 FILLER_27_787 ();
 sg13g2_decap_8 FILLER_27_794 ();
 sg13g2_decap_8 FILLER_27_801 ();
 sg13g2_decap_8 FILLER_27_808 ();
 sg13g2_decap_8 FILLER_27_815 ();
 sg13g2_decap_8 FILLER_27_822 ();
 sg13g2_decap_8 FILLER_27_829 ();
 sg13g2_decap_8 FILLER_27_836 ();
 sg13g2_decap_8 FILLER_27_843 ();
 sg13g2_decap_8 FILLER_27_850 ();
 sg13g2_decap_4 FILLER_27_857 ();
 sg13g2_fill_1 FILLER_27_861 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_4 FILLER_28_7 ();
 sg13g2_fill_1 FILLER_28_15 ();
 sg13g2_fill_1 FILLER_28_37 ();
 sg13g2_fill_2 FILLER_28_46 ();
 sg13g2_fill_2 FILLER_28_76 ();
 sg13g2_decap_4 FILLER_28_116 ();
 sg13g2_decap_4 FILLER_28_125 ();
 sg13g2_fill_2 FILLER_28_129 ();
 sg13g2_fill_1 FILLER_28_134 ();
 sg13g2_decap_8 FILLER_28_143 ();
 sg13g2_decap_4 FILLER_28_150 ();
 sg13g2_fill_1 FILLER_28_154 ();
 sg13g2_decap_4 FILLER_28_163 ();
 sg13g2_fill_2 FILLER_28_167 ();
 sg13g2_decap_4 FILLER_28_174 ();
 sg13g2_fill_2 FILLER_28_184 ();
 sg13g2_fill_1 FILLER_28_195 ();
 sg13g2_decap_8 FILLER_28_201 ();
 sg13g2_fill_1 FILLER_28_208 ();
 sg13g2_fill_2 FILLER_28_219 ();
 sg13g2_fill_2 FILLER_28_264 ();
 sg13g2_decap_8 FILLER_28_275 ();
 sg13g2_fill_2 FILLER_28_300 ();
 sg13g2_fill_1 FILLER_28_302 ();
 sg13g2_fill_1 FILLER_28_317 ();
 sg13g2_decap_8 FILLER_28_344 ();
 sg13g2_fill_2 FILLER_28_355 ();
 sg13g2_fill_1 FILLER_28_392 ();
 sg13g2_fill_1 FILLER_28_412 ();
 sg13g2_fill_1 FILLER_28_434 ();
 sg13g2_decap_8 FILLER_28_460 ();
 sg13g2_fill_2 FILLER_28_467 ();
 sg13g2_fill_1 FILLER_28_469 ();
 sg13g2_fill_2 FILLER_28_560 ();
 sg13g2_fill_2 FILLER_28_638 ();
 sg13g2_fill_1 FILLER_28_699 ();
 sg13g2_fill_1 FILLER_28_711 ();
 sg13g2_fill_2 FILLER_28_738 ();
 sg13g2_decap_8 FILLER_28_775 ();
 sg13g2_decap_8 FILLER_28_782 ();
 sg13g2_decap_8 FILLER_28_789 ();
 sg13g2_decap_8 FILLER_28_796 ();
 sg13g2_decap_8 FILLER_28_803 ();
 sg13g2_decap_8 FILLER_28_810 ();
 sg13g2_decap_8 FILLER_28_817 ();
 sg13g2_decap_8 FILLER_28_824 ();
 sg13g2_decap_8 FILLER_28_831 ();
 sg13g2_decap_8 FILLER_28_838 ();
 sg13g2_decap_8 FILLER_28_845 ();
 sg13g2_decap_8 FILLER_28_852 ();
 sg13g2_fill_2 FILLER_28_859 ();
 sg13g2_fill_1 FILLER_28_861 ();
 sg13g2_fill_1 FILLER_29_26 ();
 sg13g2_decap_8 FILLER_29_53 ();
 sg13g2_decap_8 FILLER_29_60 ();
 sg13g2_fill_1 FILLER_29_67 ();
 sg13g2_fill_1 FILLER_29_78 ();
 sg13g2_decap_4 FILLER_29_83 ();
 sg13g2_fill_1 FILLER_29_87 ();
 sg13g2_fill_2 FILLER_29_93 ();
 sg13g2_decap_8 FILLER_29_113 ();
 sg13g2_fill_2 FILLER_29_143 ();
 sg13g2_fill_1 FILLER_29_145 ();
 sg13g2_fill_1 FILLER_29_164 ();
 sg13g2_fill_2 FILLER_29_183 ();
 sg13g2_fill_1 FILLER_29_185 ();
 sg13g2_decap_4 FILLER_29_214 ();
 sg13g2_fill_1 FILLER_29_282 ();
 sg13g2_fill_1 FILLER_29_306 ();
 sg13g2_fill_2 FILLER_29_326 ();
 sg13g2_decap_8 FILLER_29_353 ();
 sg13g2_fill_1 FILLER_29_360 ();
 sg13g2_fill_2 FILLER_29_374 ();
 sg13g2_fill_2 FILLER_29_423 ();
 sg13g2_fill_1 FILLER_29_425 ();
 sg13g2_fill_2 FILLER_29_445 ();
 sg13g2_decap_8 FILLER_29_473 ();
 sg13g2_fill_2 FILLER_29_480 ();
 sg13g2_fill_1 FILLER_29_482 ();
 sg13g2_fill_1 FILLER_29_519 ();
 sg13g2_decap_4 FILLER_29_617 ();
 sg13g2_fill_2 FILLER_29_621 ();
 sg13g2_fill_1 FILLER_29_678 ();
 sg13g2_fill_1 FILLER_29_709 ();
 sg13g2_fill_1 FILLER_29_736 ();
 sg13g2_fill_2 FILLER_29_755 ();
 sg13g2_fill_1 FILLER_29_757 ();
 sg13g2_decap_8 FILLER_29_784 ();
 sg13g2_decap_8 FILLER_29_791 ();
 sg13g2_decap_8 FILLER_29_798 ();
 sg13g2_decap_8 FILLER_29_805 ();
 sg13g2_decap_8 FILLER_29_812 ();
 sg13g2_decap_8 FILLER_29_819 ();
 sg13g2_decap_8 FILLER_29_826 ();
 sg13g2_decap_8 FILLER_29_833 ();
 sg13g2_decap_8 FILLER_29_840 ();
 sg13g2_decap_8 FILLER_29_847 ();
 sg13g2_decap_8 FILLER_29_854 ();
 sg13g2_fill_1 FILLER_29_861 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_4 FILLER_30_7 ();
 sg13g2_fill_2 FILLER_30_15 ();
 sg13g2_fill_1 FILLER_30_34 ();
 sg13g2_decap_4 FILLER_30_58 ();
 sg13g2_fill_2 FILLER_30_62 ();
 sg13g2_fill_2 FILLER_30_74 ();
 sg13g2_fill_2 FILLER_30_119 ();
 sg13g2_fill_1 FILLER_30_121 ();
 sg13g2_decap_4 FILLER_30_126 ();
 sg13g2_decap_4 FILLER_30_152 ();
 sg13g2_fill_2 FILLER_30_171 ();
 sg13g2_fill_2 FILLER_30_185 ();
 sg13g2_decap_8 FILLER_30_200 ();
 sg13g2_fill_1 FILLER_30_207 ();
 sg13g2_fill_2 FILLER_30_218 ();
 sg13g2_fill_2 FILLER_30_237 ();
 sg13g2_fill_1 FILLER_30_265 ();
 sg13g2_decap_8 FILLER_30_270 ();
 sg13g2_decap_4 FILLER_30_277 ();
 sg13g2_fill_2 FILLER_30_329 ();
 sg13g2_fill_1 FILLER_30_331 ();
 sg13g2_fill_2 FILLER_30_341 ();
 sg13g2_fill_2 FILLER_30_348 ();
 sg13g2_fill_1 FILLER_30_350 ();
 sg13g2_decap_4 FILLER_30_360 ();
 sg13g2_fill_2 FILLER_30_374 ();
 sg13g2_fill_1 FILLER_30_376 ();
 sg13g2_fill_1 FILLER_30_407 ();
 sg13g2_fill_1 FILLER_30_472 ();
 sg13g2_fill_1 FILLER_30_576 ();
 sg13g2_fill_1 FILLER_30_589 ();
 sg13g2_decap_8 FILLER_30_616 ();
 sg13g2_fill_2 FILLER_30_623 ();
 sg13g2_fill_2 FILLER_30_634 ();
 sg13g2_fill_1 FILLER_30_636 ();
 sg13g2_decap_8 FILLER_30_645 ();
 sg13g2_fill_1 FILLER_30_687 ();
 sg13g2_fill_2 FILLER_30_747 ();
 sg13g2_decap_8 FILLER_30_784 ();
 sg13g2_decap_8 FILLER_30_791 ();
 sg13g2_decap_8 FILLER_30_798 ();
 sg13g2_decap_8 FILLER_30_805 ();
 sg13g2_decap_8 FILLER_30_812 ();
 sg13g2_decap_8 FILLER_30_819 ();
 sg13g2_decap_8 FILLER_30_826 ();
 sg13g2_decap_8 FILLER_30_833 ();
 sg13g2_decap_8 FILLER_30_840 ();
 sg13g2_decap_8 FILLER_30_847 ();
 sg13g2_decap_8 FILLER_30_854 ();
 sg13g2_fill_1 FILLER_30_861 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_7 ();
 sg13g2_fill_2 FILLER_31_11 ();
 sg13g2_fill_1 FILLER_31_13 ();
 sg13g2_decap_4 FILLER_31_18 ();
 sg13g2_fill_1 FILLER_31_22 ();
 sg13g2_fill_2 FILLER_31_46 ();
 sg13g2_decap_4 FILLER_31_58 ();
 sg13g2_fill_1 FILLER_31_67 ();
 sg13g2_fill_1 FILLER_31_87 ();
 sg13g2_decap_8 FILLER_31_92 ();
 sg13g2_decap_8 FILLER_31_99 ();
 sg13g2_decap_8 FILLER_31_106 ();
 sg13g2_fill_2 FILLER_31_113 ();
 sg13g2_fill_2 FILLER_31_131 ();
 sg13g2_fill_1 FILLER_31_133 ();
 sg13g2_fill_1 FILLER_31_143 ();
 sg13g2_fill_1 FILLER_31_170 ();
 sg13g2_fill_1 FILLER_31_176 ();
 sg13g2_fill_1 FILLER_31_182 ();
 sg13g2_decap_4 FILLER_31_198 ();
 sg13g2_fill_2 FILLER_31_202 ();
 sg13g2_fill_2 FILLER_31_214 ();
 sg13g2_decap_8 FILLER_31_339 ();
 sg13g2_fill_1 FILLER_31_346 ();
 sg13g2_fill_2 FILLER_31_351 ();
 sg13g2_fill_1 FILLER_31_353 ();
 sg13g2_fill_2 FILLER_31_422 ();
 sg13g2_fill_2 FILLER_31_454 ();
 sg13g2_fill_2 FILLER_31_482 ();
 sg13g2_fill_1 FILLER_31_484 ();
 sg13g2_decap_4 FILLER_31_540 ();
 sg13g2_fill_2 FILLER_31_544 ();
 sg13g2_decap_4 FILLER_31_549 ();
 sg13g2_decap_8 FILLER_31_566 ();
 sg13g2_fill_2 FILLER_31_577 ();
 sg13g2_decap_8 FILLER_31_611 ();
 sg13g2_decap_8 FILLER_31_618 ();
 sg13g2_fill_2 FILLER_31_625 ();
 sg13g2_fill_2 FILLER_31_688 ();
 sg13g2_fill_2 FILLER_31_695 ();
 sg13g2_fill_2 FILLER_31_724 ();
 sg13g2_fill_2 FILLER_31_753 ();
 sg13g2_decap_8 FILLER_31_791 ();
 sg13g2_decap_8 FILLER_31_798 ();
 sg13g2_decap_8 FILLER_31_805 ();
 sg13g2_decap_8 FILLER_31_812 ();
 sg13g2_decap_8 FILLER_31_819 ();
 sg13g2_decap_8 FILLER_31_826 ();
 sg13g2_decap_8 FILLER_31_833 ();
 sg13g2_decap_8 FILLER_31_840 ();
 sg13g2_decap_8 FILLER_31_847 ();
 sg13g2_decap_8 FILLER_31_854 ();
 sg13g2_fill_1 FILLER_31_861 ();
 sg13g2_decap_4 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_44 ();
 sg13g2_decap_8 FILLER_32_51 ();
 sg13g2_decap_8 FILLER_32_58 ();
 sg13g2_fill_2 FILLER_32_65 ();
 sg13g2_decap_4 FILLER_32_77 ();
 sg13g2_fill_2 FILLER_32_81 ();
 sg13g2_decap_4 FILLER_32_86 ();
 sg13g2_fill_2 FILLER_32_90 ();
 sg13g2_decap_4 FILLER_32_125 ();
 sg13g2_fill_1 FILLER_32_139 ();
 sg13g2_decap_4 FILLER_32_151 ();
 sg13g2_decap_8 FILLER_32_159 ();
 sg13g2_decap_8 FILLER_32_166 ();
 sg13g2_fill_1 FILLER_32_173 ();
 sg13g2_fill_2 FILLER_32_198 ();
 sg13g2_fill_1 FILLER_32_200 ();
 sg13g2_decap_8 FILLER_32_205 ();
 sg13g2_fill_2 FILLER_32_212 ();
 sg13g2_fill_2 FILLER_32_217 ();
 sg13g2_fill_1 FILLER_32_219 ();
 sg13g2_decap_8 FILLER_32_258 ();
 sg13g2_fill_1 FILLER_32_265 ();
 sg13g2_fill_2 FILLER_32_278 ();
 sg13g2_fill_1 FILLER_32_280 ();
 sg13g2_decap_4 FILLER_32_321 ();
 sg13g2_fill_2 FILLER_32_329 ();
 sg13g2_fill_1 FILLER_32_331 ();
 sg13g2_decap_4 FILLER_32_353 ();
 sg13g2_fill_1 FILLER_32_357 ();
 sg13g2_decap_4 FILLER_32_379 ();
 sg13g2_fill_2 FILLER_32_383 ();
 sg13g2_fill_2 FILLER_32_389 ();
 sg13g2_fill_1 FILLER_32_391 ();
 sg13g2_decap_4 FILLER_32_401 ();
 sg13g2_fill_2 FILLER_32_405 ();
 sg13g2_fill_2 FILLER_32_432 ();
 sg13g2_decap_8 FILLER_32_452 ();
 sg13g2_decap_4 FILLER_32_459 ();
 sg13g2_fill_1 FILLER_32_463 ();
 sg13g2_decap_8 FILLER_32_486 ();
 sg13g2_fill_2 FILLER_32_493 ();
 sg13g2_fill_1 FILLER_32_513 ();
 sg13g2_fill_2 FILLER_32_534 ();
 sg13g2_decap_8 FILLER_32_540 ();
 sg13g2_fill_1 FILLER_32_547 ();
 sg13g2_fill_1 FILLER_32_583 ();
 sg13g2_decap_8 FILLER_32_626 ();
 sg13g2_decap_4 FILLER_32_633 ();
 sg13g2_fill_1 FILLER_32_641 ();
 sg13g2_fill_2 FILLER_32_650 ();
 sg13g2_fill_2 FILLER_32_717 ();
 sg13g2_fill_1 FILLER_32_719 ();
 sg13g2_decap_8 FILLER_32_790 ();
 sg13g2_decap_8 FILLER_32_797 ();
 sg13g2_decap_8 FILLER_32_804 ();
 sg13g2_decap_8 FILLER_32_811 ();
 sg13g2_decap_8 FILLER_32_818 ();
 sg13g2_decap_8 FILLER_32_825 ();
 sg13g2_decap_8 FILLER_32_832 ();
 sg13g2_decap_8 FILLER_32_839 ();
 sg13g2_decap_8 FILLER_32_846 ();
 sg13g2_decap_8 FILLER_32_853 ();
 sg13g2_fill_2 FILLER_32_860 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_38 ();
 sg13g2_fill_1 FILLER_33_44 ();
 sg13g2_fill_2 FILLER_33_74 ();
 sg13g2_decap_4 FILLER_33_98 ();
 sg13g2_fill_1 FILLER_33_102 ();
 sg13g2_decap_4 FILLER_33_127 ();
 sg13g2_fill_2 FILLER_33_131 ();
 sg13g2_fill_2 FILLER_33_148 ();
 sg13g2_fill_1 FILLER_33_150 ();
 sg13g2_decap_4 FILLER_33_156 ();
 sg13g2_fill_1 FILLER_33_160 ();
 sg13g2_decap_8 FILLER_33_166 ();
 sg13g2_fill_2 FILLER_33_173 ();
 sg13g2_fill_1 FILLER_33_175 ();
 sg13g2_fill_2 FILLER_33_188 ();
 sg13g2_decap_4 FILLER_33_195 ();
 sg13g2_decap_8 FILLER_33_204 ();
 sg13g2_fill_2 FILLER_33_215 ();
 sg13g2_fill_1 FILLER_33_217 ();
 sg13g2_fill_1 FILLER_33_257 ();
 sg13g2_decap_8 FILLER_33_261 ();
 sg13g2_decap_4 FILLER_33_268 ();
 sg13g2_fill_1 FILLER_33_272 ();
 sg13g2_decap_4 FILLER_33_277 ();
 sg13g2_fill_1 FILLER_33_300 ();
 sg13g2_fill_2 FILLER_33_310 ();
 sg13g2_fill_1 FILLER_33_312 ();
 sg13g2_fill_2 FILLER_33_353 ();
 sg13g2_fill_1 FILLER_33_355 ();
 sg13g2_fill_2 FILLER_33_379 ();
 sg13g2_decap_4 FILLER_33_454 ();
 sg13g2_fill_1 FILLER_33_458 ();
 sg13g2_fill_2 FILLER_33_490 ();
 sg13g2_fill_2 FILLER_33_523 ();
 sg13g2_decap_4 FILLER_33_559 ();
 sg13g2_fill_1 FILLER_33_563 ();
 sg13g2_decap_8 FILLER_33_568 ();
 sg13g2_decap_4 FILLER_33_575 ();
 sg13g2_fill_2 FILLER_33_593 ();
 sg13g2_fill_1 FILLER_33_595 ();
 sg13g2_decap_4 FILLER_33_605 ();
 sg13g2_fill_2 FILLER_33_609 ();
 sg13g2_decap_4 FILLER_33_615 ();
 sg13g2_fill_2 FILLER_33_619 ();
 sg13g2_decap_8 FILLER_33_626 ();
 sg13g2_fill_1 FILLER_33_683 ();
 sg13g2_fill_2 FILLER_33_728 ();
 sg13g2_fill_1 FILLER_33_760 ();
 sg13g2_fill_2 FILLER_33_765 ();
 sg13g2_fill_1 FILLER_33_767 ();
 sg13g2_decap_8 FILLER_33_798 ();
 sg13g2_decap_8 FILLER_33_805 ();
 sg13g2_decap_8 FILLER_33_812 ();
 sg13g2_decap_8 FILLER_33_819 ();
 sg13g2_decap_8 FILLER_33_826 ();
 sg13g2_decap_8 FILLER_33_833 ();
 sg13g2_decap_8 FILLER_33_840 ();
 sg13g2_decap_8 FILLER_33_847 ();
 sg13g2_decap_8 FILLER_33_854 ();
 sg13g2_fill_1 FILLER_33_861 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_7 ();
 sg13g2_fill_1 FILLER_34_14 ();
 sg13g2_fill_1 FILLER_34_56 ();
 sg13g2_fill_1 FILLER_34_68 ();
 sg13g2_fill_2 FILLER_34_84 ();
 sg13g2_fill_1 FILLER_34_98 ();
 sg13g2_fill_2 FILLER_34_106 ();
 sg13g2_decap_8 FILLER_34_134 ();
 sg13g2_fill_2 FILLER_34_141 ();
 sg13g2_decap_4 FILLER_34_151 ();
 sg13g2_fill_1 FILLER_34_155 ();
 sg13g2_decap_8 FILLER_34_201 ();
 sg13g2_fill_1 FILLER_34_208 ();
 sg13g2_fill_2 FILLER_34_220 ();
 sg13g2_fill_1 FILLER_34_222 ();
 sg13g2_fill_2 FILLER_34_289 ();
 sg13g2_fill_1 FILLER_34_291 ();
 sg13g2_fill_2 FILLER_34_337 ();
 sg13g2_fill_1 FILLER_34_339 ();
 sg13g2_fill_2 FILLER_34_358 ();
 sg13g2_fill_2 FILLER_34_386 ();
 sg13g2_decap_8 FILLER_34_463 ();
 sg13g2_fill_2 FILLER_34_474 ();
 sg13g2_decap_8 FILLER_34_494 ();
 sg13g2_fill_1 FILLER_34_501 ();
 sg13g2_decap_4 FILLER_34_506 ();
 sg13g2_decap_8 FILLER_34_535 ();
 sg13g2_decap_4 FILLER_34_542 ();
 sg13g2_fill_1 FILLER_34_546 ();
 sg13g2_fill_2 FILLER_34_559 ();
 sg13g2_fill_2 FILLER_34_565 ();
 sg13g2_fill_1 FILLER_34_567 ();
 sg13g2_fill_1 FILLER_34_646 ();
 sg13g2_fill_1 FILLER_34_655 ();
 sg13g2_fill_2 FILLER_34_691 ();
 sg13g2_decap_4 FILLER_34_719 ();
 sg13g2_fill_1 FILLER_34_775 ();
 sg13g2_decap_8 FILLER_34_806 ();
 sg13g2_decap_8 FILLER_34_813 ();
 sg13g2_decap_8 FILLER_34_820 ();
 sg13g2_decap_8 FILLER_34_827 ();
 sg13g2_decap_8 FILLER_34_834 ();
 sg13g2_decap_8 FILLER_34_841 ();
 sg13g2_decap_8 FILLER_34_848 ();
 sg13g2_decap_8 FILLER_34_855 ();
 sg13g2_decap_4 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_45 ();
 sg13g2_fill_2 FILLER_35_51 ();
 sg13g2_fill_1 FILLER_35_53 ();
 sg13g2_fill_2 FILLER_35_77 ();
 sg13g2_fill_2 FILLER_35_113 ();
 sg13g2_decap_4 FILLER_35_136 ();
 sg13g2_fill_1 FILLER_35_140 ();
 sg13g2_decap_4 FILLER_35_146 ();
 sg13g2_fill_1 FILLER_35_150 ();
 sg13g2_fill_2 FILLER_35_156 ();
 sg13g2_fill_1 FILLER_35_158 ();
 sg13g2_decap_4 FILLER_35_175 ();
 sg13g2_fill_1 FILLER_35_205 ();
 sg13g2_fill_2 FILLER_35_244 ();
 sg13g2_decap_4 FILLER_35_277 ();
 sg13g2_fill_1 FILLER_35_281 ();
 sg13g2_fill_2 FILLER_35_295 ();
 sg13g2_fill_1 FILLER_35_332 ();
 sg13g2_decap_8 FILLER_35_354 ();
 sg13g2_decap_8 FILLER_35_361 ();
 sg13g2_fill_1 FILLER_35_368 ();
 sg13g2_decap_8 FILLER_35_377 ();
 sg13g2_fill_2 FILLER_35_396 ();
 sg13g2_fill_2 FILLER_35_470 ();
 sg13g2_fill_1 FILLER_35_472 ();
 sg13g2_fill_1 FILLER_35_481 ();
 sg13g2_fill_2 FILLER_35_487 ();
 sg13g2_fill_1 FILLER_35_507 ();
 sg13g2_fill_2 FILLER_35_534 ();
 sg13g2_decap_8 FILLER_35_540 ();
 sg13g2_fill_2 FILLER_35_547 ();
 sg13g2_decap_8 FILLER_35_584 ();
 sg13g2_fill_1 FILLER_35_591 ();
 sg13g2_fill_2 FILLER_35_634 ();
 sg13g2_fill_1 FILLER_35_645 ();
 sg13g2_fill_2 FILLER_35_659 ();
 sg13g2_decap_4 FILLER_35_704 ();
 sg13g2_fill_1 FILLER_35_708 ();
 sg13g2_fill_1 FILLER_35_723 ();
 sg13g2_fill_1 FILLER_35_729 ();
 sg13g2_fill_2 FILLER_35_767 ();
 sg13g2_decap_8 FILLER_35_810 ();
 sg13g2_decap_8 FILLER_35_817 ();
 sg13g2_decap_8 FILLER_35_824 ();
 sg13g2_decap_8 FILLER_35_831 ();
 sg13g2_decap_8 FILLER_35_838 ();
 sg13g2_decap_8 FILLER_35_845 ();
 sg13g2_decap_8 FILLER_35_852 ();
 sg13g2_fill_2 FILLER_35_859 ();
 sg13g2_fill_1 FILLER_35_861 ();
 sg13g2_fill_2 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_46 ();
 sg13g2_fill_2 FILLER_36_57 ();
 sg13g2_fill_2 FILLER_36_71 ();
 sg13g2_fill_1 FILLER_36_73 ();
 sg13g2_fill_2 FILLER_36_89 ();
 sg13g2_fill_1 FILLER_36_96 ();
 sg13g2_decap_8 FILLER_36_108 ();
 sg13g2_fill_2 FILLER_36_115 ();
 sg13g2_decap_4 FILLER_36_122 ();
 sg13g2_decap_4 FILLER_36_152 ();
 sg13g2_fill_2 FILLER_36_156 ();
 sg13g2_decap_8 FILLER_36_169 ();
 sg13g2_decap_8 FILLER_36_176 ();
 sg13g2_fill_2 FILLER_36_183 ();
 sg13g2_fill_1 FILLER_36_185 ();
 sg13g2_fill_1 FILLER_36_196 ();
 sg13g2_fill_2 FILLER_36_290 ();
 sg13g2_fill_1 FILLER_36_305 ();
 sg13g2_fill_2 FILLER_36_310 ();
 sg13g2_fill_1 FILLER_36_312 ();
 sg13g2_fill_2 FILLER_36_345 ();
 sg13g2_fill_2 FILLER_36_359 ();
 sg13g2_fill_1 FILLER_36_361 ();
 sg13g2_fill_2 FILLER_36_388 ();
 sg13g2_fill_1 FILLER_36_390 ();
 sg13g2_fill_1 FILLER_36_401 ();
 sg13g2_fill_2 FILLER_36_464 ();
 sg13g2_fill_2 FILLER_36_523 ();
 sg13g2_fill_1 FILLER_36_618 ();
 sg13g2_decap_4 FILLER_36_672 ();
 sg13g2_decap_4 FILLER_36_685 ();
 sg13g2_fill_1 FILLER_36_689 ();
 sg13g2_fill_1 FILLER_36_725 ();
 sg13g2_fill_2 FILLER_36_744 ();
 sg13g2_fill_1 FILLER_36_746 ();
 sg13g2_decap_8 FILLER_36_817 ();
 sg13g2_decap_8 FILLER_36_824 ();
 sg13g2_decap_8 FILLER_36_831 ();
 sg13g2_decap_8 FILLER_36_838 ();
 sg13g2_decap_8 FILLER_36_845 ();
 sg13g2_decap_8 FILLER_36_852 ();
 sg13g2_fill_2 FILLER_36_859 ();
 sg13g2_fill_1 FILLER_36_861 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_2 ();
 sg13g2_fill_1 FILLER_37_44 ();
 sg13g2_fill_2 FILLER_37_67 ();
 sg13g2_decap_4 FILLER_37_116 ();
 sg13g2_fill_2 FILLER_37_120 ();
 sg13g2_decap_8 FILLER_37_137 ();
 sg13g2_decap_8 FILLER_37_144 ();
 sg13g2_decap_8 FILLER_37_151 ();
 sg13g2_decap_4 FILLER_37_158 ();
 sg13g2_fill_2 FILLER_37_162 ();
 sg13g2_fill_2 FILLER_37_175 ();
 sg13g2_fill_1 FILLER_37_177 ();
 sg13g2_fill_2 FILLER_37_202 ();
 sg13g2_fill_1 FILLER_37_223 ();
 sg13g2_fill_1 FILLER_37_273 ();
 sg13g2_decap_8 FILLER_37_278 ();
 sg13g2_decap_4 FILLER_37_285 ();
 sg13g2_fill_2 FILLER_37_325 ();
 sg13g2_fill_2 FILLER_37_362 ();
 sg13g2_fill_1 FILLER_37_401 ();
 sg13g2_fill_2 FILLER_37_411 ();
 sg13g2_fill_1 FILLER_37_413 ();
 sg13g2_fill_1 FILLER_37_422 ();
 sg13g2_fill_2 FILLER_37_429 ();
 sg13g2_fill_1 FILLER_37_431 ();
 sg13g2_fill_2 FILLER_37_455 ();
 sg13g2_fill_2 FILLER_37_479 ();
 sg13g2_fill_1 FILLER_37_481 ();
 sg13g2_decap_8 FILLER_37_486 ();
 sg13g2_decap_8 FILLER_37_493 ();
 sg13g2_decap_8 FILLER_37_500 ();
 sg13g2_decap_8 FILLER_37_507 ();
 sg13g2_fill_2 FILLER_37_514 ();
 sg13g2_fill_1 FILLER_37_516 ();
 sg13g2_fill_2 FILLER_37_525 ();
 sg13g2_decap_4 FILLER_37_575 ();
 sg13g2_fill_2 FILLER_37_579 ();
 sg13g2_decap_8 FILLER_37_585 ();
 sg13g2_decap_8 FILLER_37_592 ();
 sg13g2_decap_8 FILLER_37_599 ();
 sg13g2_decap_8 FILLER_37_606 ();
 sg13g2_decap_8 FILLER_37_613 ();
 sg13g2_decap_8 FILLER_37_620 ();
 sg13g2_decap_8 FILLER_37_627 ();
 sg13g2_fill_1 FILLER_37_646 ();
 sg13g2_fill_1 FILLER_37_669 ();
 sg13g2_decap_4 FILLER_37_707 ();
 sg13g2_fill_2 FILLER_37_711 ();
 sg13g2_fill_1 FILLER_37_722 ();
 sg13g2_fill_2 FILLER_37_728 ();
 sg13g2_fill_1 FILLER_37_730 ();
 sg13g2_fill_2 FILLER_37_757 ();
 sg13g2_fill_1 FILLER_37_759 ();
 sg13g2_decap_8 FILLER_37_795 ();
 sg13g2_decap_8 FILLER_37_802 ();
 sg13g2_decap_8 FILLER_37_809 ();
 sg13g2_decap_8 FILLER_37_816 ();
 sg13g2_decap_8 FILLER_37_823 ();
 sg13g2_decap_8 FILLER_37_830 ();
 sg13g2_decap_8 FILLER_37_837 ();
 sg13g2_decap_8 FILLER_37_844 ();
 sg13g2_decap_8 FILLER_37_851 ();
 sg13g2_decap_4 FILLER_37_858 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_38 ();
 sg13g2_fill_2 FILLER_38_45 ();
 sg13g2_fill_1 FILLER_38_52 ();
 sg13g2_decap_8 FILLER_38_61 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_fill_1 FILLER_38_72 ();
 sg13g2_decap_8 FILLER_38_159 ();
 sg13g2_fill_2 FILLER_38_177 ();
 sg13g2_fill_1 FILLER_38_179 ();
 sg13g2_fill_1 FILLER_38_223 ();
 sg13g2_fill_2 FILLER_38_295 ();
 sg13g2_fill_1 FILLER_38_297 ();
 sg13g2_fill_1 FILLER_38_307 ();
 sg13g2_fill_1 FILLER_38_321 ();
 sg13g2_fill_2 FILLER_38_356 ();
 sg13g2_fill_1 FILLER_38_358 ();
 sg13g2_fill_1 FILLER_38_363 ();
 sg13g2_fill_1 FILLER_38_368 ();
 sg13g2_fill_1 FILLER_38_418 ();
 sg13g2_decap_8 FILLER_38_481 ();
 sg13g2_fill_1 FILLER_38_488 ();
 sg13g2_decap_8 FILLER_38_493 ();
 sg13g2_fill_1 FILLER_38_505 ();
 sg13g2_decap_4 FILLER_38_532 ();
 sg13g2_fill_1 FILLER_38_536 ();
 sg13g2_decap_4 FILLER_38_563 ();
 sg13g2_fill_2 FILLER_38_567 ();
 sg13g2_decap_8 FILLER_38_603 ();
 sg13g2_decap_8 FILLER_38_610 ();
 sg13g2_fill_2 FILLER_38_617 ();
 sg13g2_decap_8 FILLER_38_623 ();
 sg13g2_fill_1 FILLER_38_630 ();
 sg13g2_fill_1 FILLER_38_657 ();
 sg13g2_fill_1 FILLER_38_721 ();
 sg13g2_fill_1 FILLER_38_732 ();
 sg13g2_fill_2 FILLER_38_751 ();
 sg13g2_decap_8 FILLER_38_788 ();
 sg13g2_decap_8 FILLER_38_795 ();
 sg13g2_decap_8 FILLER_38_802 ();
 sg13g2_decap_8 FILLER_38_809 ();
 sg13g2_decap_8 FILLER_38_816 ();
 sg13g2_decap_8 FILLER_38_823 ();
 sg13g2_decap_8 FILLER_38_830 ();
 sg13g2_decap_8 FILLER_38_837 ();
 sg13g2_decap_8 FILLER_38_844 ();
 sg13g2_decap_8 FILLER_38_851 ();
 sg13g2_decap_4 FILLER_38_858 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_fill_2 FILLER_39_21 ();
 sg13g2_fill_1 FILLER_39_27 ();
 sg13g2_fill_2 FILLER_39_36 ();
 sg13g2_fill_1 FILLER_39_38 ();
 sg13g2_decap_4 FILLER_39_55 ();
 sg13g2_decap_4 FILLER_39_69 ();
 sg13g2_fill_1 FILLER_39_73 ();
 sg13g2_decap_4 FILLER_39_100 ();
 sg13g2_fill_1 FILLER_39_104 ();
 sg13g2_fill_2 FILLER_39_109 ();
 sg13g2_fill_1 FILLER_39_111 ();
 sg13g2_decap_8 FILLER_39_124 ();
 sg13g2_decap_8 FILLER_39_135 ();
 sg13g2_decap_4 FILLER_39_142 ();
 sg13g2_fill_1 FILLER_39_146 ();
 sg13g2_fill_2 FILLER_39_157 ();
 sg13g2_fill_1 FILLER_39_159 ();
 sg13g2_fill_2 FILLER_39_164 ();
 sg13g2_decap_8 FILLER_39_181 ();
 sg13g2_decap_8 FILLER_39_188 ();
 sg13g2_decap_4 FILLER_39_195 ();
 sg13g2_decap_8 FILLER_39_260 ();
 sg13g2_fill_2 FILLER_39_267 ();
 sg13g2_decap_4 FILLER_39_275 ();
 sg13g2_fill_1 FILLER_39_279 ();
 sg13g2_decap_8 FILLER_39_284 ();
 sg13g2_fill_2 FILLER_39_291 ();
 sg13g2_fill_2 FILLER_39_308 ();
 sg13g2_fill_1 FILLER_39_341 ();
 sg13g2_fill_1 FILLER_39_393 ();
 sg13g2_fill_2 FILLER_39_400 ();
 sg13g2_decap_4 FILLER_39_406 ();
 sg13g2_fill_2 FILLER_39_420 ();
 sg13g2_fill_1 FILLER_39_422 ();
 sg13g2_decap_8 FILLER_39_457 ();
 sg13g2_decap_8 FILLER_39_464 ();
 sg13g2_fill_2 FILLER_39_476 ();
 sg13g2_fill_1 FILLER_39_478 ();
 sg13g2_decap_8 FILLER_39_513 ();
 sg13g2_decap_4 FILLER_39_528 ();
 sg13g2_fill_2 FILLER_39_537 ();
 sg13g2_fill_1 FILLER_39_539 ();
 sg13g2_fill_2 FILLER_39_548 ();
 sg13g2_decap_4 FILLER_39_555 ();
 sg13g2_decap_8 FILLER_39_569 ();
 sg13g2_fill_2 FILLER_39_576 ();
 sg13g2_decap_4 FILLER_39_590 ();
 sg13g2_fill_2 FILLER_39_606 ();
 sg13g2_fill_1 FILLER_39_634 ();
 sg13g2_fill_2 FILLER_39_660 ();
 sg13g2_fill_1 FILLER_39_662 ();
 sg13g2_decap_8 FILLER_39_675 ();
 sg13g2_fill_2 FILLER_39_682 ();
 sg13g2_fill_2 FILLER_39_702 ();
 sg13g2_fill_1 FILLER_39_704 ();
 sg13g2_decap_4 FILLER_39_714 ();
 sg13g2_fill_1 FILLER_39_763 ();
 sg13g2_decap_8 FILLER_39_790 ();
 sg13g2_decap_8 FILLER_39_797 ();
 sg13g2_decap_8 FILLER_39_804 ();
 sg13g2_decap_8 FILLER_39_811 ();
 sg13g2_decap_8 FILLER_39_818 ();
 sg13g2_decap_8 FILLER_39_825 ();
 sg13g2_decap_8 FILLER_39_832 ();
 sg13g2_decap_8 FILLER_39_839 ();
 sg13g2_decap_8 FILLER_39_846 ();
 sg13g2_decap_8 FILLER_39_853 ();
 sg13g2_fill_2 FILLER_39_860 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_67 ();
 sg13g2_decap_8 FILLER_40_74 ();
 sg13g2_decap_4 FILLER_40_81 ();
 sg13g2_fill_1 FILLER_40_89 ();
 sg13g2_fill_2 FILLER_40_99 ();
 sg13g2_decap_4 FILLER_40_116 ();
 sg13g2_decap_8 FILLER_40_135 ();
 sg13g2_fill_2 FILLER_40_142 ();
 sg13g2_fill_2 FILLER_40_153 ();
 sg13g2_fill_2 FILLER_40_169 ();
 sg13g2_fill_1 FILLER_40_171 ();
 sg13g2_fill_2 FILLER_40_202 ();
 sg13g2_fill_1 FILLER_40_204 ();
 sg13g2_fill_2 FILLER_40_218 ();
 sg13g2_fill_1 FILLER_40_224 ();
 sg13g2_decap_8 FILLER_40_279 ();
 sg13g2_decap_8 FILLER_40_286 ();
 sg13g2_fill_1 FILLER_40_301 ();
 sg13g2_fill_2 FILLER_40_306 ();
 sg13g2_decap_4 FILLER_40_315 ();
 sg13g2_fill_1 FILLER_40_319 ();
 sg13g2_decap_4 FILLER_40_324 ();
 sg13g2_fill_1 FILLER_40_328 ();
 sg13g2_fill_2 FILLER_40_364 ();
 sg13g2_fill_1 FILLER_40_366 ();
 sg13g2_fill_2 FILLER_40_388 ();
 sg13g2_fill_1 FILLER_40_390 ();
 sg13g2_decap_8 FILLER_40_415 ();
 sg13g2_fill_1 FILLER_40_448 ();
 sg13g2_fill_2 FILLER_40_454 ();
 sg13g2_fill_1 FILLER_40_472 ();
 sg13g2_decap_8 FILLER_40_485 ();
 sg13g2_decap_4 FILLER_40_492 ();
 sg13g2_decap_8 FILLER_40_508 ();
 sg13g2_decap_4 FILLER_40_515 ();
 sg13g2_fill_2 FILLER_40_519 ();
 sg13g2_decap_4 FILLER_40_540 ();
 sg13g2_decap_4 FILLER_40_552 ();
 sg13g2_fill_2 FILLER_40_576 ();
 sg13g2_fill_1 FILLER_40_578 ();
 sg13g2_fill_2 FILLER_40_587 ();
 sg13g2_fill_1 FILLER_40_589 ();
 sg13g2_fill_1 FILLER_40_595 ();
 sg13g2_decap_8 FILLER_40_621 ();
 sg13g2_fill_2 FILLER_40_628 ();
 sg13g2_decap_8 FILLER_40_638 ();
 sg13g2_decap_4 FILLER_40_651 ();
 sg13g2_fill_2 FILLER_40_663 ();
 sg13g2_decap_8 FILLER_40_681 ();
 sg13g2_decap_8 FILLER_40_708 ();
 sg13g2_decap_8 FILLER_40_715 ();
 sg13g2_decap_8 FILLER_40_722 ();
 sg13g2_decap_4 FILLER_40_733 ();
 sg13g2_fill_2 FILLER_40_737 ();
 sg13g2_fill_1 FILLER_40_743 ();
 sg13g2_decap_8 FILLER_40_779 ();
 sg13g2_decap_8 FILLER_40_786 ();
 sg13g2_decap_8 FILLER_40_793 ();
 sg13g2_decap_8 FILLER_40_800 ();
 sg13g2_decap_8 FILLER_40_807 ();
 sg13g2_decap_8 FILLER_40_814 ();
 sg13g2_decap_8 FILLER_40_821 ();
 sg13g2_decap_8 FILLER_40_828 ();
 sg13g2_decap_8 FILLER_40_835 ();
 sg13g2_decap_8 FILLER_40_842 ();
 sg13g2_decap_8 FILLER_40_849 ();
 sg13g2_decap_4 FILLER_40_856 ();
 sg13g2_fill_2 FILLER_40_860 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_fill_2 FILLER_41_7 ();
 sg13g2_fill_1 FILLER_41_9 ();
 sg13g2_fill_2 FILLER_41_23 ();
 sg13g2_fill_1 FILLER_41_25 ();
 sg13g2_fill_2 FILLER_41_33 ();
 sg13g2_fill_2 FILLER_41_45 ();
 sg13g2_decap_4 FILLER_41_52 ();
 sg13g2_decap_8 FILLER_41_76 ();
 sg13g2_decap_4 FILLER_41_83 ();
 sg13g2_fill_1 FILLER_41_87 ();
 sg13g2_decap_8 FILLER_41_101 ();
 sg13g2_decap_8 FILLER_41_108 ();
 sg13g2_decap_8 FILLER_41_115 ();
 sg13g2_fill_2 FILLER_41_122 ();
 sg13g2_decap_8 FILLER_41_140 ();
 sg13g2_fill_2 FILLER_41_147 ();
 sg13g2_fill_2 FILLER_41_157 ();
 sg13g2_fill_2 FILLER_41_167 ();
 sg13g2_decap_4 FILLER_41_177 ();
 sg13g2_fill_2 FILLER_41_186 ();
 sg13g2_fill_1 FILLER_41_188 ();
 sg13g2_decap_8 FILLER_41_193 ();
 sg13g2_decap_4 FILLER_41_200 ();
 sg13g2_fill_2 FILLER_41_204 ();
 sg13g2_fill_1 FILLER_41_211 ();
 sg13g2_fill_2 FILLER_41_218 ();
 sg13g2_fill_1 FILLER_41_220 ();
 sg13g2_fill_1 FILLER_41_230 ();
 sg13g2_decap_4 FILLER_41_235 ();
 sg13g2_decap_8 FILLER_41_248 ();
 sg13g2_fill_2 FILLER_41_255 ();
 sg13g2_fill_2 FILLER_41_262 ();
 sg13g2_fill_2 FILLER_41_276 ();
 sg13g2_decap_8 FILLER_41_299 ();
 sg13g2_fill_2 FILLER_41_306 ();
 sg13g2_fill_1 FILLER_41_318 ();
 sg13g2_fill_2 FILLER_41_325 ();
 sg13g2_fill_1 FILLER_41_327 ();
 sg13g2_fill_2 FILLER_41_338 ();
 sg13g2_fill_1 FILLER_41_355 ();
 sg13g2_decap_8 FILLER_41_386 ();
 sg13g2_fill_1 FILLER_41_412 ();
 sg13g2_decap_8 FILLER_41_417 ();
 sg13g2_fill_2 FILLER_41_424 ();
 sg13g2_decap_8 FILLER_41_439 ();
 sg13g2_decap_8 FILLER_41_452 ();
 sg13g2_decap_8 FILLER_41_484 ();
 sg13g2_fill_2 FILLER_41_491 ();
 sg13g2_fill_1 FILLER_41_493 ();
 sg13g2_fill_1 FILLER_41_499 ();
 sg13g2_fill_1 FILLER_41_516 ();
 sg13g2_decap_4 FILLER_41_524 ();
 sg13g2_fill_2 FILLER_41_528 ();
 sg13g2_decap_8 FILLER_41_535 ();
 sg13g2_decap_8 FILLER_41_542 ();
 sg13g2_fill_1 FILLER_41_549 ();
 sg13g2_fill_1 FILLER_41_555 ();
 sg13g2_decap_4 FILLER_41_565 ();
 sg13g2_fill_1 FILLER_41_569 ();
 sg13g2_decap_4 FILLER_41_590 ();
 sg13g2_fill_1 FILLER_41_594 ();
 sg13g2_fill_2 FILLER_41_611 ();
 sg13g2_fill_1 FILLER_41_618 ();
 sg13g2_decap_8 FILLER_41_627 ();
 sg13g2_decap_4 FILLER_41_634 ();
 sg13g2_fill_1 FILLER_41_638 ();
 sg13g2_fill_2 FILLER_41_660 ();
 sg13g2_fill_1 FILLER_41_662 ();
 sg13g2_decap_8 FILLER_41_671 ();
 sg13g2_decap_8 FILLER_41_678 ();
 sg13g2_fill_1 FILLER_41_685 ();
 sg13g2_decap_4 FILLER_41_700 ();
 sg13g2_fill_1 FILLER_41_704 ();
 sg13g2_decap_8 FILLER_41_718 ();
 sg13g2_decap_8 FILLER_41_725 ();
 sg13g2_decap_4 FILLER_41_732 ();
 sg13g2_decap_4 FILLER_41_744 ();
 sg13g2_fill_2 FILLER_41_748 ();
 sg13g2_fill_2 FILLER_41_759 ();
 sg13g2_fill_1 FILLER_41_761 ();
 sg13g2_decap_8 FILLER_41_775 ();
 sg13g2_decap_8 FILLER_41_782 ();
 sg13g2_decap_8 FILLER_41_789 ();
 sg13g2_decap_8 FILLER_41_796 ();
 sg13g2_decap_8 FILLER_41_803 ();
 sg13g2_decap_8 FILLER_41_810 ();
 sg13g2_decap_8 FILLER_41_817 ();
 sg13g2_decap_8 FILLER_41_824 ();
 sg13g2_decap_8 FILLER_41_831 ();
 sg13g2_decap_8 FILLER_41_838 ();
 sg13g2_decap_8 FILLER_41_845 ();
 sg13g2_decap_8 FILLER_41_852 ();
 sg13g2_fill_2 FILLER_41_859 ();
 sg13g2_fill_1 FILLER_41_861 ();
 sg13g2_fill_1 FILLER_42_49 ();
 sg13g2_decap_4 FILLER_42_87 ();
 sg13g2_fill_2 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_fill_1 FILLER_42_105 ();
 sg13g2_fill_2 FILLER_42_136 ();
 sg13g2_fill_2 FILLER_42_144 ();
 sg13g2_decap_8 FILLER_42_154 ();
 sg13g2_fill_1 FILLER_42_161 ();
 sg13g2_decap_8 FILLER_42_202 ();
 sg13g2_decap_4 FILLER_42_225 ();
 sg13g2_fill_2 FILLER_42_240 ();
 sg13g2_fill_2 FILLER_42_247 ();
 sg13g2_decap_4 FILLER_42_275 ();
 sg13g2_fill_1 FILLER_42_279 ();
 sg13g2_decap_4 FILLER_42_333 ();
 sg13g2_fill_1 FILLER_42_337 ();
 sg13g2_decap_4 FILLER_42_344 ();
 sg13g2_fill_1 FILLER_42_348 ();
 sg13g2_fill_2 FILLER_42_362 ();
 sg13g2_decap_4 FILLER_42_377 ();
 sg13g2_fill_1 FILLER_42_381 ();
 sg13g2_decap_4 FILLER_42_395 ();
 sg13g2_fill_2 FILLER_42_407 ();
 sg13g2_fill_1 FILLER_42_415 ();
 sg13g2_fill_2 FILLER_42_442 ();
 sg13g2_fill_1 FILLER_42_460 ();
 sg13g2_decap_4 FILLER_42_469 ();
 sg13g2_fill_2 FILLER_42_473 ();
 sg13g2_fill_2 FILLER_42_480 ();
 sg13g2_decap_8 FILLER_42_488 ();
 sg13g2_fill_2 FILLER_42_495 ();
 sg13g2_fill_2 FILLER_42_517 ();
 sg13g2_fill_1 FILLER_42_519 ();
 sg13g2_fill_1 FILLER_42_530 ();
 sg13g2_decap_4 FILLER_42_544 ();
 sg13g2_fill_1 FILLER_42_558 ();
 sg13g2_decap_4 FILLER_42_568 ();
 sg13g2_fill_1 FILLER_42_572 ();
 sg13g2_decap_8 FILLER_42_579 ();
 sg13g2_fill_1 FILLER_42_586 ();
 sg13g2_fill_2 FILLER_42_595 ();
 sg13g2_fill_1 FILLER_42_597 ();
 sg13g2_decap_4 FILLER_42_618 ();
 sg13g2_fill_1 FILLER_42_622 ();
 sg13g2_decap_8 FILLER_42_637 ();
 sg13g2_decap_4 FILLER_42_644 ();
 sg13g2_fill_1 FILLER_42_648 ();
 sg13g2_decap_4 FILLER_42_671 ();
 sg13g2_fill_1 FILLER_42_675 ();
 sg13g2_decap_4 FILLER_42_684 ();
 sg13g2_fill_2 FILLER_42_704 ();
 sg13g2_fill_1 FILLER_42_706 ();
 sg13g2_decap_8 FILLER_42_726 ();
 sg13g2_decap_4 FILLER_42_733 ();
 sg13g2_fill_2 FILLER_42_737 ();
 sg13g2_decap_8 FILLER_42_766 ();
 sg13g2_fill_1 FILLER_42_773 ();
 sg13g2_decap_8 FILLER_42_786 ();
 sg13g2_fill_2 FILLER_42_793 ();
 sg13g2_decap_8 FILLER_42_803 ();
 sg13g2_fill_2 FILLER_42_810 ();
 sg13g2_fill_1 FILLER_42_812 ();
 sg13g2_fill_2 FILLER_42_817 ();
 sg13g2_fill_1 FILLER_42_819 ();
 sg13g2_decap_8 FILLER_42_828 ();
 sg13g2_decap_8 FILLER_42_835 ();
 sg13g2_decap_8 FILLER_42_842 ();
 sg13g2_decap_8 FILLER_42_849 ();
 sg13g2_decap_4 FILLER_42_856 ();
 sg13g2_fill_2 FILLER_42_860 ();
 sg13g2_decap_4 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_43_4 ();
 sg13g2_fill_2 FILLER_43_45 ();
 sg13g2_fill_2 FILLER_43_84 ();
 sg13g2_fill_1 FILLER_43_86 ();
 sg13g2_fill_1 FILLER_43_108 ();
 sg13g2_decap_8 FILLER_43_122 ();
 sg13g2_decap_4 FILLER_43_129 ();
 sg13g2_decap_8 FILLER_43_137 ();
 sg13g2_decap_8 FILLER_43_161 ();
 sg13g2_decap_8 FILLER_43_178 ();
 sg13g2_fill_2 FILLER_43_185 ();
 sg13g2_decap_8 FILLER_43_195 ();
 sg13g2_decap_4 FILLER_43_202 ();
 sg13g2_fill_1 FILLER_43_206 ();
 sg13g2_fill_2 FILLER_43_227 ();
 sg13g2_fill_1 FILLER_43_234 ();
 sg13g2_fill_2 FILLER_43_241 ();
 sg13g2_decap_8 FILLER_43_255 ();
 sg13g2_fill_2 FILLER_43_262 ();
 sg13g2_fill_1 FILLER_43_264 ();
 sg13g2_decap_8 FILLER_43_268 ();
 sg13g2_fill_2 FILLER_43_275 ();
 sg13g2_fill_1 FILLER_43_277 ();
 sg13g2_decap_8 FILLER_43_288 ();
 sg13g2_decap_4 FILLER_43_295 ();
 sg13g2_fill_1 FILLER_43_299 ();
 sg13g2_decap_8 FILLER_43_322 ();
 sg13g2_decap_8 FILLER_43_329 ();
 sg13g2_fill_1 FILLER_43_336 ();
 sg13g2_fill_2 FILLER_43_341 ();
 sg13g2_fill_2 FILLER_43_352 ();
 sg13g2_fill_1 FILLER_43_354 ();
 sg13g2_decap_4 FILLER_43_359 ();
 sg13g2_fill_1 FILLER_43_367 ();
 sg13g2_decap_8 FILLER_43_435 ();
 sg13g2_decap_4 FILLER_43_442 ();
 sg13g2_fill_2 FILLER_43_446 ();
 sg13g2_decap_8 FILLER_43_454 ();
 sg13g2_decap_4 FILLER_43_461 ();
 sg13g2_fill_2 FILLER_43_465 ();
 sg13g2_fill_2 FILLER_43_478 ();
 sg13g2_decap_4 FILLER_43_502 ();
 sg13g2_fill_2 FILLER_43_506 ();
 sg13g2_decap_4 FILLER_43_513 ();
 sg13g2_fill_2 FILLER_43_517 ();
 sg13g2_fill_1 FILLER_43_531 ();
 sg13g2_decap_8 FILLER_43_537 ();
 sg13g2_decap_4 FILLER_43_544 ();
 sg13g2_fill_2 FILLER_43_548 ();
 sg13g2_fill_2 FILLER_43_555 ();
 sg13g2_decap_8 FILLER_43_569 ();
 sg13g2_decap_4 FILLER_43_576 ();
 sg13g2_fill_2 FILLER_43_594 ();
 sg13g2_fill_1 FILLER_43_596 ();
 sg13g2_fill_2 FILLER_43_624 ();
 sg13g2_fill_1 FILLER_43_626 ();
 sg13g2_decap_8 FILLER_43_640 ();
 sg13g2_decap_4 FILLER_43_647 ();
 sg13g2_fill_2 FILLER_43_651 ();
 sg13g2_decap_4 FILLER_43_666 ();
 sg13g2_fill_2 FILLER_43_670 ();
 sg13g2_decap_8 FILLER_43_682 ();
 sg13g2_fill_1 FILLER_43_699 ();
 sg13g2_fill_2 FILLER_43_705 ();
 sg13g2_fill_1 FILLER_43_707 ();
 sg13g2_fill_2 FILLER_43_726 ();
 sg13g2_fill_1 FILLER_43_728 ();
 sg13g2_decap_4 FILLER_43_737 ();
 sg13g2_decap_4 FILLER_43_746 ();
 sg13g2_fill_1 FILLER_43_785 ();
 sg13g2_fill_1 FILLER_43_810 ();
 sg13g2_decap_8 FILLER_43_836 ();
 sg13g2_decap_8 FILLER_43_851 ();
 sg13g2_decap_4 FILLER_43_858 ();
 sg13g2_fill_1 FILLER_44_26 ();
 sg13g2_fill_1 FILLER_44_36 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_fill_1 FILLER_44_63 ();
 sg13g2_fill_1 FILLER_44_72 ();
 sg13g2_fill_2 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_112 ();
 sg13g2_fill_2 FILLER_44_119 ();
 sg13g2_fill_1 FILLER_44_121 ();
 sg13g2_decap_8 FILLER_44_126 ();
 sg13g2_fill_2 FILLER_44_133 ();
 sg13g2_fill_1 FILLER_44_140 ();
 sg13g2_decap_8 FILLER_44_160 ();
 sg13g2_decap_8 FILLER_44_167 ();
 sg13g2_decap_4 FILLER_44_174 ();
 sg13g2_fill_2 FILLER_44_178 ();
 sg13g2_fill_2 FILLER_44_183 ();
 sg13g2_fill_1 FILLER_44_185 ();
 sg13g2_decap_4 FILLER_44_192 ();
 sg13g2_fill_1 FILLER_44_196 ();
 sg13g2_decap_8 FILLER_44_206 ();
 sg13g2_decap_4 FILLER_44_213 ();
 sg13g2_fill_2 FILLER_44_217 ();
 sg13g2_decap_4 FILLER_44_223 ();
 sg13g2_fill_1 FILLER_44_227 ();
 sg13g2_fill_2 FILLER_44_234 ();
 sg13g2_fill_1 FILLER_44_236 ();
 sg13g2_decap_8 FILLER_44_245 ();
 sg13g2_fill_2 FILLER_44_252 ();
 sg13g2_decap_4 FILLER_44_275 ();
 sg13g2_fill_2 FILLER_44_279 ();
 sg13g2_fill_2 FILLER_44_286 ();
 sg13g2_fill_2 FILLER_44_292 ();
 sg13g2_fill_2 FILLER_44_299 ();
 sg13g2_fill_1 FILLER_44_316 ();
 sg13g2_fill_2 FILLER_44_327 ();
 sg13g2_fill_1 FILLER_44_329 ();
 sg13g2_fill_2 FILLER_44_370 ();
 sg13g2_fill_1 FILLER_44_372 ();
 sg13g2_decap_4 FILLER_44_392 ();
 sg13g2_fill_2 FILLER_44_396 ();
 sg13g2_decap_8 FILLER_44_435 ();
 sg13g2_decap_8 FILLER_44_442 ();
 sg13g2_decap_8 FILLER_44_449 ();
 sg13g2_fill_2 FILLER_44_456 ();
 sg13g2_fill_1 FILLER_44_458 ();
 sg13g2_decap_4 FILLER_44_464 ();
 sg13g2_fill_1 FILLER_44_569 ();
 sg13g2_fill_2 FILLER_44_575 ();
 sg13g2_decap_8 FILLER_44_588 ();
 sg13g2_fill_2 FILLER_44_595 ();
 sg13g2_fill_1 FILLER_44_597 ();
 sg13g2_fill_2 FILLER_44_606 ();
 sg13g2_fill_2 FILLER_44_612 ();
 sg13g2_fill_1 FILLER_44_614 ();
 sg13g2_fill_1 FILLER_44_619 ();
 sg13g2_decap_8 FILLER_44_640 ();
 sg13g2_decap_4 FILLER_44_647 ();
 sg13g2_fill_1 FILLER_44_662 ();
 sg13g2_fill_1 FILLER_44_673 ();
 sg13g2_decap_8 FILLER_44_688 ();
 sg13g2_fill_1 FILLER_44_695 ();
 sg13g2_decap_4 FILLER_44_710 ();
 sg13g2_fill_2 FILLER_44_714 ();
 sg13g2_fill_1 FILLER_44_734 ();
 sg13g2_decap_8 FILLER_44_745 ();
 sg13g2_decap_8 FILLER_44_760 ();
 sg13g2_decap_4 FILLER_44_789 ();
 sg13g2_fill_2 FILLER_44_793 ();
 sg13g2_decap_4 FILLER_44_803 ();
 sg13g2_fill_1 FILLER_44_807 ();
 sg13g2_decap_8 FILLER_44_816 ();
 sg13g2_fill_2 FILLER_44_823 ();
 sg13g2_decap_8 FILLER_44_838 ();
 sg13g2_decap_8 FILLER_44_845 ();
 sg13g2_decap_8 FILLER_44_852 ();
 sg13g2_fill_2 FILLER_44_859 ();
 sg13g2_fill_1 FILLER_44_861 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_fill_1 FILLER_45_7 ();
 sg13g2_fill_2 FILLER_45_51 ();
 sg13g2_decap_4 FILLER_45_58 ();
 sg13g2_fill_2 FILLER_45_62 ();
 sg13g2_fill_1 FILLER_45_72 ();
 sg13g2_decap_4 FILLER_45_82 ();
 sg13g2_fill_2 FILLER_45_90 ();
 sg13g2_fill_1 FILLER_45_92 ();
 sg13g2_decap_8 FILLER_45_98 ();
 sg13g2_decap_4 FILLER_45_105 ();
 sg13g2_fill_2 FILLER_45_109 ();
 sg13g2_decap_8 FILLER_45_137 ();
 sg13g2_fill_2 FILLER_45_162 ();
 sg13g2_fill_1 FILLER_45_164 ();
 sg13g2_fill_2 FILLER_45_186 ();
 sg13g2_fill_2 FILLER_45_205 ();
 sg13g2_fill_1 FILLER_45_207 ();
 sg13g2_decap_4 FILLER_45_234 ();
 sg13g2_fill_1 FILLER_45_238 ();
 sg13g2_decap_8 FILLER_45_251 ();
 sg13g2_decap_8 FILLER_45_258 ();
 sg13g2_decap_8 FILLER_45_265 ();
 sg13g2_fill_1 FILLER_45_272 ();
 sg13g2_decap_8 FILLER_45_294 ();
 sg13g2_fill_2 FILLER_45_301 ();
 sg13g2_decap_8 FILLER_45_320 ();
 sg13g2_decap_8 FILLER_45_327 ();
 sg13g2_fill_2 FILLER_45_367 ();
 sg13g2_fill_2 FILLER_45_390 ();
 sg13g2_fill_1 FILLER_45_392 ();
 sg13g2_fill_1 FILLER_45_433 ();
 sg13g2_fill_2 FILLER_45_464 ();
 sg13g2_fill_1 FILLER_45_475 ();
 sg13g2_decap_8 FILLER_45_480 ();
 sg13g2_decap_8 FILLER_45_487 ();
 sg13g2_decap_8 FILLER_45_494 ();
 sg13g2_fill_2 FILLER_45_501 ();
 sg13g2_decap_4 FILLER_45_521 ();
 sg13g2_fill_2 FILLER_45_525 ();
 sg13g2_fill_2 FILLER_45_531 ();
 sg13g2_fill_1 FILLER_45_533 ();
 sg13g2_decap_4 FILLER_45_543 ();
 sg13g2_fill_1 FILLER_45_547 ();
 sg13g2_fill_2 FILLER_45_556 ();
 sg13g2_fill_1 FILLER_45_558 ();
 sg13g2_fill_2 FILLER_45_564 ();
 sg13g2_decap_4 FILLER_45_589 ();
 sg13g2_fill_1 FILLER_45_593 ();
 sg13g2_fill_1 FILLER_45_610 ();
 sg13g2_fill_2 FILLER_45_619 ();
 sg13g2_fill_2 FILLER_45_626 ();
 sg13g2_fill_2 FILLER_45_632 ();
 sg13g2_decap_4 FILLER_45_652 ();
 sg13g2_fill_1 FILLER_45_656 ();
 sg13g2_decap_8 FILLER_45_667 ();
 sg13g2_fill_1 FILLER_45_674 ();
 sg13g2_decap_8 FILLER_45_684 ();
 sg13g2_fill_2 FILLER_45_691 ();
 sg13g2_fill_1 FILLER_45_693 ();
 sg13g2_decap_4 FILLER_45_722 ();
 sg13g2_decap_8 FILLER_45_736 ();
 sg13g2_fill_2 FILLER_45_743 ();
 sg13g2_fill_2 FILLER_45_751 ();
 sg13g2_decap_8 FILLER_45_759 ();
 sg13g2_decap_8 FILLER_45_766 ();
 sg13g2_fill_2 FILLER_45_773 ();
 sg13g2_fill_1 FILLER_45_775 ();
 sg13g2_fill_2 FILLER_45_788 ();
 sg13g2_fill_1 FILLER_45_790 ();
 sg13g2_decap_8 FILLER_45_808 ();
 sg13g2_decap_4 FILLER_45_815 ();
 sg13g2_fill_1 FILLER_45_819 ();
 sg13g2_decap_8 FILLER_45_853 ();
 sg13g2_fill_2 FILLER_45_860 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_4 FILLER_46_7 ();
 sg13g2_decap_4 FILLER_46_15 ();
 sg13g2_fill_2 FILLER_46_19 ();
 sg13g2_fill_2 FILLER_46_30 ();
 sg13g2_fill_1 FILLER_46_32 ();
 sg13g2_decap_8 FILLER_46_52 ();
 sg13g2_fill_2 FILLER_46_111 ();
 sg13g2_fill_1 FILLER_46_113 ();
 sg13g2_decap_4 FILLER_46_151 ();
 sg13g2_decap_8 FILLER_46_160 ();
 sg13g2_decap_4 FILLER_46_167 ();
 sg13g2_fill_2 FILLER_46_171 ();
 sg13g2_fill_2 FILLER_46_182 ();
 sg13g2_fill_1 FILLER_46_184 ();
 sg13g2_fill_2 FILLER_46_216 ();
 sg13g2_fill_2 FILLER_46_227 ();
 sg13g2_decap_8 FILLER_46_233 ();
 sg13g2_decap_8 FILLER_46_240 ();
 sg13g2_fill_2 FILLER_46_247 ();
 sg13g2_decap_8 FILLER_46_270 ();
 sg13g2_decap_8 FILLER_46_277 ();
 sg13g2_fill_2 FILLER_46_284 ();
 sg13g2_decap_4 FILLER_46_290 ();
 sg13g2_fill_1 FILLER_46_294 ();
 sg13g2_fill_2 FILLER_46_303 ();
 sg13g2_decap_8 FILLER_46_319 ();
 sg13g2_decap_4 FILLER_46_326 ();
 sg13g2_fill_2 FILLER_46_334 ();
 sg13g2_fill_1 FILLER_46_336 ();
 sg13g2_fill_2 FILLER_46_346 ();
 sg13g2_fill_2 FILLER_46_399 ();
 sg13g2_fill_1 FILLER_46_410 ();
 sg13g2_decap_8 FILLER_46_419 ();
 sg13g2_decap_8 FILLER_46_426 ();
 sg13g2_fill_2 FILLER_46_433 ();
 sg13g2_fill_1 FILLER_46_435 ();
 sg13g2_fill_2 FILLER_46_441 ();
 sg13g2_fill_1 FILLER_46_443 ();
 sg13g2_decap_4 FILLER_46_454 ();
 sg13g2_fill_1 FILLER_46_468 ();
 sg13g2_fill_1 FILLER_46_480 ();
 sg13g2_decap_4 FILLER_46_485 ();
 sg13g2_fill_1 FILLER_46_504 ();
 sg13g2_decap_8 FILLER_46_524 ();
 sg13g2_decap_4 FILLER_46_531 ();
 sg13g2_decap_8 FILLER_46_560 ();
 sg13g2_decap_8 FILLER_46_567 ();
 sg13g2_decap_4 FILLER_46_585 ();
 sg13g2_fill_2 FILLER_46_589 ();
 sg13g2_decap_4 FILLER_46_599 ();
 sg13g2_decap_8 FILLER_46_609 ();
 sg13g2_decap_8 FILLER_46_616 ();
 sg13g2_decap_4 FILLER_46_641 ();
 sg13g2_fill_1 FILLER_46_690 ();
 sg13g2_fill_2 FILLER_46_697 ();
 sg13g2_decap_4 FILLER_46_704 ();
 sg13g2_fill_2 FILLER_46_708 ();
 sg13g2_fill_2 FILLER_46_719 ();
 sg13g2_fill_1 FILLER_46_721 ();
 sg13g2_fill_1 FILLER_46_727 ();
 sg13g2_fill_2 FILLER_46_738 ();
 sg13g2_fill_1 FILLER_46_740 ();
 sg13g2_decap_4 FILLER_46_754 ();
 sg13g2_fill_2 FILLER_46_772 ();
 sg13g2_fill_2 FILLER_46_782 ();
 sg13g2_fill_1 FILLER_46_784 ();
 sg13g2_decap_8 FILLER_46_791 ();
 sg13g2_fill_1 FILLER_46_819 ();
 sg13g2_decap_4 FILLER_46_824 ();
 sg13g2_fill_1 FILLER_46_828 ();
 sg13g2_decap_8 FILLER_46_833 ();
 sg13g2_decap_8 FILLER_46_840 ();
 sg13g2_decap_8 FILLER_46_847 ();
 sg13g2_decap_8 FILLER_46_854 ();
 sg13g2_fill_1 FILLER_46_861 ();
 sg13g2_fill_2 FILLER_47_56 ();
 sg13g2_fill_1 FILLER_47_58 ();
 sg13g2_fill_2 FILLER_47_82 ();
 sg13g2_fill_1 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_116 ();
 sg13g2_decap_8 FILLER_47_123 ();
 sg13g2_decap_4 FILLER_47_130 ();
 sg13g2_fill_1 FILLER_47_134 ();
 sg13g2_fill_1 FILLER_47_149 ();
 sg13g2_decap_4 FILLER_47_164 ();
 sg13g2_fill_1 FILLER_47_198 ();
 sg13g2_decap_8 FILLER_47_204 ();
 sg13g2_decap_8 FILLER_47_211 ();
 sg13g2_decap_4 FILLER_47_271 ();
 sg13g2_fill_1 FILLER_47_275 ();
 sg13g2_fill_1 FILLER_47_285 ();
 sg13g2_fill_2 FILLER_47_296 ();
 sg13g2_fill_1 FILLER_47_298 ();
 sg13g2_fill_1 FILLER_47_313 ();
 sg13g2_decap_8 FILLER_47_324 ();
 sg13g2_fill_2 FILLER_47_331 ();
 sg13g2_fill_1 FILLER_47_333 ();
 sg13g2_fill_1 FILLER_47_356 ();
 sg13g2_fill_2 FILLER_47_372 ();
 sg13g2_fill_1 FILLER_47_409 ();
 sg13g2_fill_2 FILLER_47_427 ();
 sg13g2_fill_1 FILLER_47_434 ();
 sg13g2_fill_2 FILLER_47_440 ();
 sg13g2_fill_1 FILLER_47_459 ();
 sg13g2_decap_4 FILLER_47_465 ();
 sg13g2_fill_2 FILLER_47_488 ();
 sg13g2_fill_1 FILLER_47_498 ();
 sg13g2_fill_1 FILLER_47_503 ();
 sg13g2_decap_8 FILLER_47_509 ();
 sg13g2_fill_2 FILLER_47_516 ();
 sg13g2_fill_1 FILLER_47_518 ();
 sg13g2_decap_8 FILLER_47_529 ();
 sg13g2_decap_8 FILLER_47_561 ();
 sg13g2_fill_1 FILLER_47_617 ();
 sg13g2_decap_8 FILLER_47_638 ();
 sg13g2_decap_8 FILLER_47_645 ();
 sg13g2_decap_4 FILLER_47_652 ();
 sg13g2_fill_2 FILLER_47_656 ();
 sg13g2_decap_8 FILLER_47_668 ();
 sg13g2_fill_2 FILLER_47_675 ();
 sg13g2_fill_1 FILLER_47_677 ();
 sg13g2_fill_1 FILLER_47_683 ();
 sg13g2_fill_2 FILLER_47_696 ();
 sg13g2_fill_1 FILLER_47_698 ();
 sg13g2_fill_2 FILLER_47_705 ();
 sg13g2_fill_1 FILLER_47_712 ();
 sg13g2_fill_2 FILLER_47_721 ();
 sg13g2_decap_4 FILLER_47_728 ();
 sg13g2_fill_1 FILLER_47_732 ();
 sg13g2_decap_4 FILLER_47_744 ();
 sg13g2_decap_8 FILLER_47_766 ();
 sg13g2_fill_1 FILLER_47_778 ();
 sg13g2_decap_8 FILLER_47_793 ();
 sg13g2_fill_2 FILLER_47_800 ();
 sg13g2_fill_1 FILLER_47_802 ();
 sg13g2_decap_4 FILLER_47_808 ();
 sg13g2_fill_2 FILLER_47_829 ();
 sg13g2_fill_1 FILLER_47_831 ();
 sg13g2_decap_8 FILLER_47_854 ();
 sg13g2_fill_1 FILLER_47_861 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_7 ();
 sg13g2_fill_1 FILLER_48_22 ();
 sg13g2_fill_2 FILLER_48_46 ();
 sg13g2_fill_1 FILLER_48_48 ();
 sg13g2_fill_1 FILLER_48_59 ();
 sg13g2_fill_1 FILLER_48_87 ();
 sg13g2_fill_1 FILLER_48_97 ();
 sg13g2_fill_2 FILLER_48_138 ();
 sg13g2_fill_1 FILLER_48_140 ();
 sg13g2_decap_4 FILLER_48_167 ();
 sg13g2_fill_2 FILLER_48_177 ();
 sg13g2_fill_1 FILLER_48_179 ();
 sg13g2_fill_1 FILLER_48_203 ();
 sg13g2_fill_2 FILLER_48_211 ();
 sg13g2_fill_1 FILLER_48_239 ();
 sg13g2_fill_2 FILLER_48_246 ();
 sg13g2_fill_2 FILLER_48_254 ();
 sg13g2_fill_1 FILLER_48_256 ();
 sg13g2_decap_8 FILLER_48_278 ();
 sg13g2_fill_2 FILLER_48_285 ();
 sg13g2_decap_4 FILLER_48_295 ();
 sg13g2_fill_2 FILLER_48_325 ();
 sg13g2_fill_2 FILLER_48_335 ();
 sg13g2_fill_1 FILLER_48_347 ();
 sg13g2_fill_2 FILLER_48_378 ();
 sg13g2_fill_1 FILLER_48_380 ();
 sg13g2_decap_8 FILLER_48_404 ();
 sg13g2_decap_4 FILLER_48_411 ();
 sg13g2_decap_8 FILLER_48_420 ();
 sg13g2_fill_1 FILLER_48_432 ();
 sg13g2_fill_2 FILLER_48_437 ();
 sg13g2_fill_1 FILLER_48_439 ();
 sg13g2_fill_1 FILLER_48_449 ();
 sg13g2_fill_2 FILLER_48_456 ();
 sg13g2_fill_1 FILLER_48_468 ();
 sg13g2_fill_2 FILLER_48_474 ();
 sg13g2_fill_1 FILLER_48_476 ();
 sg13g2_decap_8 FILLER_48_482 ();
 sg13g2_decap_4 FILLER_48_489 ();
 sg13g2_fill_1 FILLER_48_493 ();
 sg13g2_decap_4 FILLER_48_499 ();
 sg13g2_decap_4 FILLER_48_508 ();
 sg13g2_fill_1 FILLER_48_512 ();
 sg13g2_fill_1 FILLER_48_536 ();
 sg13g2_decap_4 FILLER_48_542 ();
 sg13g2_decap_4 FILLER_48_551 ();
 sg13g2_fill_1 FILLER_48_555 ();
 sg13g2_fill_2 FILLER_48_561 ();
 sg13g2_decap_8 FILLER_48_567 ();
 sg13g2_fill_1 FILLER_48_574 ();
 sg13g2_decap_8 FILLER_48_584 ();
 sg13g2_decap_8 FILLER_48_596 ();
 sg13g2_decap_8 FILLER_48_603 ();
 sg13g2_fill_2 FILLER_48_614 ();
 sg13g2_fill_2 FILLER_48_626 ();
 sg13g2_fill_1 FILLER_48_628 ();
 sg13g2_decap_4 FILLER_48_634 ();
 sg13g2_fill_1 FILLER_48_638 ();
 sg13g2_fill_2 FILLER_48_648 ();
 sg13g2_fill_1 FILLER_48_650 ();
 sg13g2_decap_8 FILLER_48_663 ();
 sg13g2_fill_2 FILLER_48_670 ();
 sg13g2_fill_1 FILLER_48_672 ();
 sg13g2_decap_4 FILLER_48_684 ();
 sg13g2_decap_4 FILLER_48_696 ();
 sg13g2_fill_2 FILLER_48_700 ();
 sg13g2_decap_4 FILLER_48_707 ();
 sg13g2_decap_4 FILLER_48_716 ();
 sg13g2_fill_1 FILLER_48_720 ();
 sg13g2_decap_8 FILLER_48_730 ();
 sg13g2_decap_8 FILLER_48_737 ();
 sg13g2_decap_4 FILLER_48_744 ();
 sg13g2_fill_2 FILLER_48_748 ();
 sg13g2_decap_4 FILLER_48_765 ();
 sg13g2_fill_1 FILLER_48_769 ();
 sg13g2_decap_8 FILLER_48_778 ();
 sg13g2_fill_1 FILLER_48_785 ();
 sg13g2_decap_4 FILLER_48_791 ();
 sg13g2_fill_2 FILLER_48_795 ();
 sg13g2_decap_4 FILLER_48_802 ();
 sg13g2_decap_8 FILLER_48_836 ();
 sg13g2_decap_4 FILLER_48_857 ();
 sg13g2_fill_1 FILLER_48_861 ();
 sg13g2_decap_4 FILLER_49_52 ();
 sg13g2_fill_1 FILLER_49_62 ();
 sg13g2_fill_1 FILLER_49_79 ();
 sg13g2_fill_1 FILLER_49_90 ();
 sg13g2_decap_4 FILLER_49_96 ();
 sg13g2_fill_2 FILLER_49_106 ();
 sg13g2_fill_1 FILLER_49_108 ();
 sg13g2_fill_2 FILLER_49_127 ();
 sg13g2_fill_1 FILLER_49_129 ();
 sg13g2_fill_1 FILLER_49_148 ();
 sg13g2_fill_1 FILLER_49_161 ();
 sg13g2_fill_2 FILLER_49_191 ();
 sg13g2_fill_1 FILLER_49_202 ();
 sg13g2_fill_2 FILLER_49_235 ();
 sg13g2_decap_8 FILLER_49_263 ();
 sg13g2_decap_4 FILLER_49_270 ();
 sg13g2_fill_2 FILLER_49_274 ();
 sg13g2_fill_1 FILLER_49_290 ();
 sg13g2_decap_8 FILLER_49_301 ();
 sg13g2_decap_4 FILLER_49_308 ();
 sg13g2_fill_1 FILLER_49_323 ();
 sg13g2_decap_4 FILLER_49_353 ();
 sg13g2_fill_1 FILLER_49_366 ();
 sg13g2_decap_8 FILLER_49_393 ();
 sg13g2_fill_2 FILLER_49_400 ();
 sg13g2_decap_8 FILLER_49_426 ();
 sg13g2_fill_1 FILLER_49_433 ();
 sg13g2_decap_8 FILLER_49_450 ();
 sg13g2_fill_1 FILLER_49_457 ();
 sg13g2_fill_2 FILLER_49_485 ();
 sg13g2_fill_1 FILLER_49_487 ();
 sg13g2_fill_1 FILLER_49_510 ();
 sg13g2_fill_1 FILLER_49_517 ();
 sg13g2_decap_8 FILLER_49_530 ();
 sg13g2_fill_2 FILLER_49_537 ();
 sg13g2_fill_1 FILLER_49_544 ();
 sg13g2_fill_1 FILLER_49_566 ();
 sg13g2_decap_4 FILLER_49_582 ();
 sg13g2_fill_1 FILLER_49_586 ();
 sg13g2_fill_2 FILLER_49_611 ();
 sg13g2_decap_8 FILLER_49_618 ();
 sg13g2_fill_2 FILLER_49_625 ();
 sg13g2_fill_1 FILLER_49_627 ();
 sg13g2_decap_4 FILLER_49_633 ();
 sg13g2_fill_1 FILLER_49_637 ();
 sg13g2_decap_8 FILLER_49_643 ();
 sg13g2_decap_4 FILLER_49_650 ();
 sg13g2_fill_2 FILLER_49_668 ();
 sg13g2_fill_1 FILLER_49_670 ();
 sg13g2_decap_4 FILLER_49_710 ();
 sg13g2_fill_1 FILLER_49_714 ();
 sg13g2_decap_4 FILLER_49_734 ();
 sg13g2_fill_1 FILLER_49_751 ();
 sg13g2_decap_8 FILLER_49_768 ();
 sg13g2_fill_2 FILLER_49_775 ();
 sg13g2_decap_8 FILLER_49_800 ();
 sg13g2_decap_4 FILLER_49_817 ();
 sg13g2_fill_2 FILLER_49_821 ();
 sg13g2_fill_2 FILLER_49_831 ();
 sg13g2_fill_2 FILLER_49_843 ();
 sg13g2_fill_1 FILLER_49_845 ();
 sg13g2_decap_8 FILLER_49_854 ();
 sg13g2_fill_1 FILLER_49_861 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_4 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_15 ();
 sg13g2_decap_4 FILLER_50_22 ();
 sg13g2_fill_2 FILLER_50_26 ();
 sg13g2_decap_4 FILLER_50_45 ();
 sg13g2_fill_2 FILLER_50_49 ();
 sg13g2_fill_2 FILLER_50_78 ();
 sg13g2_fill_2 FILLER_50_92 ();
 sg13g2_decap_4 FILLER_50_104 ();
 sg13g2_fill_1 FILLER_50_108 ();
 sg13g2_decap_8 FILLER_50_122 ();
 sg13g2_fill_2 FILLER_50_129 ();
 sg13g2_fill_1 FILLER_50_155 ();
 sg13g2_decap_4 FILLER_50_161 ();
 sg13g2_fill_2 FILLER_50_165 ();
 sg13g2_fill_2 FILLER_50_176 ();
 sg13g2_fill_2 FILLER_50_183 ();
 sg13g2_fill_2 FILLER_50_199 ();
 sg13g2_fill_1 FILLER_50_211 ();
 sg13g2_decap_4 FILLER_50_242 ();
 sg13g2_fill_2 FILLER_50_246 ();
 sg13g2_fill_1 FILLER_50_252 ();
 sg13g2_decap_8 FILLER_50_274 ();
 sg13g2_fill_2 FILLER_50_281 ();
 sg13g2_fill_2 FILLER_50_289 ();
 sg13g2_decap_4 FILLER_50_296 ();
 sg13g2_fill_2 FILLER_50_342 ();
 sg13g2_fill_1 FILLER_50_344 ();
 sg13g2_fill_2 FILLER_50_398 ();
 sg13g2_fill_2 FILLER_50_428 ();
 sg13g2_decap_8 FILLER_50_441 ();
 sg13g2_decap_8 FILLER_50_448 ();
 sg13g2_decap_4 FILLER_50_455 ();
 sg13g2_fill_2 FILLER_50_459 ();
 sg13g2_decap_8 FILLER_50_471 ();
 sg13g2_decap_8 FILLER_50_478 ();
 sg13g2_fill_1 FILLER_50_485 ();
 sg13g2_fill_2 FILLER_50_491 ();
 sg13g2_fill_1 FILLER_50_498 ();
 sg13g2_decap_8 FILLER_50_504 ();
 sg13g2_fill_1 FILLER_50_511 ();
 sg13g2_decap_8 FILLER_50_517 ();
 sg13g2_fill_2 FILLER_50_535 ();
 sg13g2_fill_1 FILLER_50_537 ();
 sg13g2_decap_8 FILLER_50_544 ();
 sg13g2_decap_8 FILLER_50_551 ();
 sg13g2_fill_2 FILLER_50_558 ();
 sg13g2_decap_4 FILLER_50_573 ();
 sg13g2_fill_2 FILLER_50_577 ();
 sg13g2_fill_2 FILLER_50_590 ();
 sg13g2_decap_8 FILLER_50_597 ();
 sg13g2_fill_2 FILLER_50_604 ();
 sg13g2_decap_4 FILLER_50_617 ();
 sg13g2_decap_4 FILLER_50_627 ();
 sg13g2_decap_8 FILLER_50_652 ();
 sg13g2_fill_2 FILLER_50_659 ();
 sg13g2_fill_2 FILLER_50_666 ();
 sg13g2_decap_4 FILLER_50_676 ();
 sg13g2_fill_2 FILLER_50_695 ();
 sg13g2_decap_8 FILLER_50_706 ();
 sg13g2_fill_2 FILLER_50_718 ();
 sg13g2_decap_8 FILLER_50_734 ();
 sg13g2_decap_8 FILLER_50_741 ();
 sg13g2_fill_2 FILLER_50_748 ();
 sg13g2_fill_1 FILLER_50_750 ();
 sg13g2_decap_4 FILLER_50_774 ();
 sg13g2_fill_2 FILLER_50_778 ();
 sg13g2_fill_1 FILLER_50_785 ();
 sg13g2_fill_2 FILLER_50_790 ();
 sg13g2_fill_1 FILLER_50_792 ();
 sg13g2_fill_1 FILLER_50_814 ();
 sg13g2_decap_8 FILLER_50_819 ();
 sg13g2_fill_1 FILLER_50_826 ();
 sg13g2_decap_8 FILLER_50_853 ();
 sg13g2_fill_2 FILLER_50_860 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_4 FILLER_51_7 ();
 sg13g2_decap_4 FILLER_51_15 ();
 sg13g2_fill_2 FILLER_51_19 ();
 sg13g2_fill_1 FILLER_51_31 ();
 sg13g2_fill_1 FILLER_51_43 ();
 sg13g2_decap_8 FILLER_51_48 ();
 sg13g2_fill_2 FILLER_51_55 ();
 sg13g2_fill_1 FILLER_51_57 ();
 sg13g2_fill_1 FILLER_51_91 ();
 sg13g2_decap_4 FILLER_51_106 ();
 sg13g2_decap_4 FILLER_51_145 ();
 sg13g2_fill_2 FILLER_51_159 ();
 sg13g2_fill_1 FILLER_51_161 ();
 sg13g2_fill_2 FILLER_51_220 ();
 sg13g2_decap_8 FILLER_51_252 ();
 sg13g2_decap_8 FILLER_51_259 ();
 sg13g2_decap_8 FILLER_51_266 ();
 sg13g2_fill_2 FILLER_51_273 ();
 sg13g2_fill_1 FILLER_51_275 ();
 sg13g2_decap_8 FILLER_51_301 ();
 sg13g2_fill_2 FILLER_51_323 ();
 sg13g2_decap_4 FILLER_51_378 ();
 sg13g2_fill_1 FILLER_51_386 ();
 sg13g2_decap_8 FILLER_51_395 ();
 sg13g2_decap_4 FILLER_51_402 ();
 sg13g2_fill_2 FILLER_51_436 ();
 sg13g2_fill_1 FILLER_51_450 ();
 sg13g2_decap_4 FILLER_51_461 ();
 sg13g2_fill_1 FILLER_51_465 ();
 sg13g2_decap_4 FILLER_51_478 ();
 sg13g2_fill_2 FILLER_51_482 ();
 sg13g2_decap_8 FILLER_51_507 ();
 sg13g2_fill_1 FILLER_51_514 ();
 sg13g2_fill_1 FILLER_51_539 ();
 sg13g2_fill_1 FILLER_51_545 ();
 sg13g2_decap_8 FILLER_51_556 ();
 sg13g2_decap_8 FILLER_51_567 ();
 sg13g2_fill_1 FILLER_51_574 ();
 sg13g2_decap_4 FILLER_51_579 ();
 sg13g2_fill_2 FILLER_51_599 ();
 sg13g2_fill_1 FILLER_51_601 ();
 sg13g2_fill_1 FILLER_51_608 ();
 sg13g2_decap_8 FILLER_51_624 ();
 sg13g2_decap_4 FILLER_51_649 ();
 sg13g2_fill_1 FILLER_51_653 ();
 sg13g2_decap_4 FILLER_51_680 ();
 sg13g2_fill_1 FILLER_51_684 ();
 sg13g2_decap_4 FILLER_51_702 ();
 sg13g2_fill_1 FILLER_51_706 ();
 sg13g2_decap_4 FILLER_51_712 ();
 sg13g2_decap_8 FILLER_51_730 ();
 sg13g2_decap_4 FILLER_51_737 ();
 sg13g2_fill_1 FILLER_51_764 ();
 sg13g2_fill_2 FILLER_51_770 ();
 sg13g2_fill_1 FILLER_51_772 ();
 sg13g2_fill_2 FILLER_51_790 ();
 sg13g2_decap_8 FILLER_51_825 ();
 sg13g2_fill_1 FILLER_51_832 ();
 sg13g2_fill_2 FILLER_51_841 ();
 sg13g2_fill_1 FILLER_51_843 ();
 sg13g2_decap_4 FILLER_51_858 ();
 sg13g2_fill_1 FILLER_52_26 ();
 sg13g2_fill_1 FILLER_52_36 ();
 sg13g2_decap_4 FILLER_52_85 ();
 sg13g2_fill_1 FILLER_52_89 ();
 sg13g2_fill_2 FILLER_52_112 ();
 sg13g2_fill_2 FILLER_52_118 ();
 sg13g2_fill_1 FILLER_52_120 ();
 sg13g2_decap_8 FILLER_52_125 ();
 sg13g2_decap_4 FILLER_52_132 ();
 sg13g2_fill_2 FILLER_52_149 ();
 sg13g2_fill_2 FILLER_52_164 ();
 sg13g2_fill_1 FILLER_52_171 ();
 sg13g2_fill_2 FILLER_52_177 ();
 sg13g2_decap_8 FILLER_52_226 ();
 sg13g2_decap_4 FILLER_52_233 ();
 sg13g2_decap_8 FILLER_52_241 ();
 sg13g2_decap_8 FILLER_52_248 ();
 sg13g2_decap_8 FILLER_52_276 ();
 sg13g2_decap_8 FILLER_52_291 ();
 sg13g2_decap_8 FILLER_52_298 ();
 sg13g2_decap_4 FILLER_52_305 ();
 sg13g2_fill_2 FILLER_52_309 ();
 sg13g2_decap_8 FILLER_52_324 ();
 sg13g2_decap_4 FILLER_52_331 ();
 sg13g2_fill_1 FILLER_52_335 ();
 sg13g2_decap_8 FILLER_52_340 ();
 sg13g2_decap_8 FILLER_52_347 ();
 sg13g2_decap_4 FILLER_52_354 ();
 sg13g2_fill_2 FILLER_52_358 ();
 sg13g2_decap_8 FILLER_52_368 ();
 sg13g2_fill_1 FILLER_52_383 ();
 sg13g2_fill_2 FILLER_52_388 ();
 sg13g2_decap_8 FILLER_52_395 ();
 sg13g2_decap_4 FILLER_52_402 ();
 sg13g2_fill_1 FILLER_52_406 ();
 sg13g2_decap_8 FILLER_52_416 ();
 sg13g2_fill_1 FILLER_52_423 ();
 sg13g2_decap_4 FILLER_52_443 ();
 sg13g2_fill_2 FILLER_52_447 ();
 sg13g2_fill_1 FILLER_52_455 ();
 sg13g2_fill_2 FILLER_52_471 ();
 sg13g2_fill_1 FILLER_52_473 ();
 sg13g2_fill_1 FILLER_52_492 ();
 sg13g2_decap_8 FILLER_52_499 ();
 sg13g2_fill_1 FILLER_52_506 ();
 sg13g2_fill_1 FILLER_52_522 ();
 sg13g2_fill_2 FILLER_52_529 ();
 sg13g2_fill_1 FILLER_52_531 ();
 sg13g2_fill_1 FILLER_52_537 ();
 sg13g2_decap_4 FILLER_52_541 ();
 sg13g2_decap_4 FILLER_52_574 ();
 sg13g2_fill_1 FILLER_52_578 ();
 sg13g2_fill_1 FILLER_52_587 ();
 sg13g2_decap_4 FILLER_52_598 ();
 sg13g2_fill_2 FILLER_52_602 ();
 sg13g2_decap_8 FILLER_52_616 ();
 sg13g2_fill_1 FILLER_52_637 ();
 sg13g2_decap_8 FILLER_52_643 ();
 sg13g2_decap_8 FILLER_52_650 ();
 sg13g2_decap_8 FILLER_52_657 ();
 sg13g2_fill_2 FILLER_52_664 ();
 sg13g2_decap_4 FILLER_52_673 ();
 sg13g2_fill_2 FILLER_52_677 ();
 sg13g2_decap_8 FILLER_52_694 ();
 sg13g2_decap_8 FILLER_52_707 ();
 sg13g2_fill_2 FILLER_52_714 ();
 sg13g2_decap_4 FILLER_52_738 ();
 sg13g2_fill_2 FILLER_52_742 ();
 sg13g2_decap_8 FILLER_52_768 ();
 sg13g2_decap_8 FILLER_52_775 ();
 sg13g2_decap_4 FILLER_52_782 ();
 sg13g2_fill_2 FILLER_52_786 ();
 sg13g2_fill_1 FILLER_52_798 ();
 sg13g2_decap_8 FILLER_52_803 ();
 sg13g2_decap_8 FILLER_52_810 ();
 sg13g2_decap_8 FILLER_52_817 ();
 sg13g2_decap_4 FILLER_52_824 ();
 sg13g2_decap_4 FILLER_52_856 ();
 sg13g2_fill_2 FILLER_52_860 ();
 sg13g2_decap_4 FILLER_53_0 ();
 sg13g2_fill_1 FILLER_53_4 ();
 sg13g2_fill_2 FILLER_53_24 ();
 sg13g2_fill_1 FILLER_53_26 ();
 sg13g2_fill_2 FILLER_53_39 ();
 sg13g2_fill_1 FILLER_53_67 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_fill_1 FILLER_53_91 ();
 sg13g2_fill_2 FILLER_53_97 ();
 sg13g2_fill_1 FILLER_53_99 ();
 sg13g2_fill_2 FILLER_53_113 ();
 sg13g2_fill_1 FILLER_53_141 ();
 sg13g2_fill_2 FILLER_53_147 ();
 sg13g2_fill_1 FILLER_53_149 ();
 sg13g2_fill_2 FILLER_53_155 ();
 sg13g2_fill_1 FILLER_53_161 ();
 sg13g2_fill_2 FILLER_53_171 ();
 sg13g2_fill_1 FILLER_53_173 ();
 sg13g2_fill_2 FILLER_53_184 ();
 sg13g2_fill_1 FILLER_53_186 ();
 sg13g2_decap_4 FILLER_53_245 ();
 sg13g2_decap_4 FILLER_53_270 ();
 sg13g2_fill_2 FILLER_53_274 ();
 sg13g2_fill_1 FILLER_53_299 ();
 sg13g2_decap_8 FILLER_53_329 ();
 sg13g2_fill_1 FILLER_53_336 ();
 sg13g2_fill_2 FILLER_53_341 ();
 sg13g2_decap_4 FILLER_53_404 ();
 sg13g2_fill_2 FILLER_53_408 ();
 sg13g2_decap_8 FILLER_53_420 ();
 sg13g2_fill_2 FILLER_53_427 ();
 sg13g2_fill_2 FILLER_53_435 ();
 sg13g2_fill_1 FILLER_53_437 ();
 sg13g2_fill_1 FILLER_53_453 ();
 sg13g2_decap_8 FILLER_53_479 ();
 sg13g2_decap_8 FILLER_53_486 ();
 sg13g2_decap_8 FILLER_53_493 ();
 sg13g2_decap_4 FILLER_53_500 ();
 sg13g2_fill_1 FILLER_53_504 ();
 sg13g2_fill_2 FILLER_53_510 ();
 sg13g2_decap_4 FILLER_53_518 ();
 sg13g2_fill_1 FILLER_53_522 ();
 sg13g2_decap_8 FILLER_53_552 ();
 sg13g2_fill_2 FILLER_53_559 ();
 sg13g2_fill_1 FILLER_53_561 ();
 sg13g2_decap_4 FILLER_53_573 ();
 sg13g2_fill_1 FILLER_53_577 ();
 sg13g2_fill_2 FILLER_53_599 ();
 sg13g2_fill_1 FILLER_53_601 ();
 sg13g2_fill_2 FILLER_53_617 ();
 sg13g2_fill_2 FILLER_53_624 ();
 sg13g2_fill_2 FILLER_53_631 ();
 sg13g2_decap_8 FILLER_53_642 ();
 sg13g2_fill_2 FILLER_53_649 ();
 sg13g2_fill_1 FILLER_53_651 ();
 sg13g2_fill_1 FILLER_53_656 ();
 sg13g2_fill_2 FILLER_53_677 ();
 sg13g2_fill_2 FILLER_53_689 ();
 sg13g2_fill_2 FILLER_53_702 ();
 sg13g2_decap_8 FILLER_53_709 ();
 sg13g2_fill_1 FILLER_53_743 ();
 sg13g2_fill_1 FILLER_53_752 ();
 sg13g2_decap_8 FILLER_53_763 ();
 sg13g2_fill_2 FILLER_53_796 ();
 sg13g2_fill_1 FILLER_53_798 ();
 sg13g2_fill_2 FILLER_53_804 ();
 sg13g2_fill_1 FILLER_53_806 ();
 sg13g2_decap_4 FILLER_53_812 ();
 sg13g2_fill_1 FILLER_53_816 ();
 sg13g2_fill_2 FILLER_53_847 ();
 sg13g2_fill_1 FILLER_53_849 ();
 sg13g2_decap_4 FILLER_53_858 ();
 sg13g2_fill_1 FILLER_54_39 ();
 sg13g2_fill_1 FILLER_54_54 ();
 sg13g2_decap_4 FILLER_54_85 ();
 sg13g2_fill_1 FILLER_54_99 ();
 sg13g2_fill_2 FILLER_54_119 ();
 sg13g2_fill_2 FILLER_54_134 ();
 sg13g2_fill_1 FILLER_54_156 ();
 sg13g2_decap_8 FILLER_54_188 ();
 sg13g2_decap_8 FILLER_54_203 ();
 sg13g2_fill_1 FILLER_54_210 ();
 sg13g2_fill_1 FILLER_54_215 ();
 sg13g2_decap_4 FILLER_54_225 ();
 sg13g2_fill_1 FILLER_54_229 ();
 sg13g2_decap_8 FILLER_54_238 ();
 sg13g2_decap_4 FILLER_54_245 ();
 sg13g2_fill_2 FILLER_54_249 ();
 sg13g2_fill_1 FILLER_54_265 ();
 sg13g2_decap_8 FILLER_54_353 ();
 sg13g2_fill_1 FILLER_54_365 ();
 sg13g2_fill_2 FILLER_54_375 ();
 sg13g2_fill_1 FILLER_54_377 ();
 sg13g2_decap_4 FILLER_54_401 ();
 sg13g2_fill_1 FILLER_54_405 ();
 sg13g2_fill_2 FILLER_54_414 ();
 sg13g2_decap_8 FILLER_54_427 ();
 sg13g2_fill_2 FILLER_54_434 ();
 sg13g2_decap_8 FILLER_54_444 ();
 sg13g2_decap_8 FILLER_54_459 ();
 sg13g2_fill_1 FILLER_54_466 ();
 sg13g2_fill_2 FILLER_54_472 ();
 sg13g2_decap_4 FILLER_54_489 ();
 sg13g2_fill_1 FILLER_54_493 ();
 sg13g2_decap_4 FILLER_54_504 ();
 sg13g2_decap_8 FILLER_54_521 ();
 sg13g2_decap_4 FILLER_54_528 ();
 sg13g2_fill_2 FILLER_54_532 ();
 sg13g2_decap_4 FILLER_54_552 ();
 sg13g2_fill_2 FILLER_54_556 ();
 sg13g2_fill_2 FILLER_54_578 ();
 sg13g2_fill_1 FILLER_54_580 ();
 sg13g2_decap_8 FILLER_54_589 ();
 sg13g2_fill_2 FILLER_54_600 ();
 sg13g2_fill_1 FILLER_54_602 ();
 sg13g2_decap_8 FILLER_54_608 ();
 sg13g2_decap_4 FILLER_54_615 ();
 sg13g2_fill_1 FILLER_54_638 ();
 sg13g2_decap_8 FILLER_54_658 ();
 sg13g2_decap_8 FILLER_54_665 ();
 sg13g2_decap_4 FILLER_54_672 ();
 sg13g2_fill_1 FILLER_54_676 ();
 sg13g2_fill_1 FILLER_54_687 ();
 sg13g2_fill_2 FILLER_54_693 ();
 sg13g2_fill_1 FILLER_54_695 ();
 sg13g2_fill_2 FILLER_54_706 ();
 sg13g2_fill_2 FILLER_54_721 ();
 sg13g2_decap_8 FILLER_54_728 ();
 sg13g2_decap_4 FILLER_54_735 ();
 sg13g2_fill_2 FILLER_54_773 ();
 sg13g2_decap_8 FILLER_54_793 ();
 sg13g2_decap_8 FILLER_54_800 ();
 sg13g2_fill_2 FILLER_54_807 ();
 sg13g2_decap_4 FILLER_54_818 ();
 sg13g2_fill_1 FILLER_54_832 ();
 sg13g2_decap_8 FILLER_54_843 ();
 sg13g2_decap_8 FILLER_54_850 ();
 sg13g2_decap_4 FILLER_54_857 ();
 sg13g2_fill_1 FILLER_54_861 ();
 sg13g2_fill_1 FILLER_55_23 ();
 sg13g2_fill_1 FILLER_55_43 ();
 sg13g2_fill_2 FILLER_55_49 ();
 sg13g2_fill_1 FILLER_55_61 ();
 sg13g2_fill_2 FILLER_55_81 ();
 sg13g2_fill_2 FILLER_55_98 ();
 sg13g2_fill_2 FILLER_55_156 ();
 sg13g2_fill_1 FILLER_55_158 ();
 sg13g2_decap_4 FILLER_55_163 ();
 sg13g2_fill_2 FILLER_55_167 ();
 sg13g2_fill_1 FILLER_55_184 ();
 sg13g2_fill_1 FILLER_55_196 ();
 sg13g2_decap_4 FILLER_55_210 ();
 sg13g2_fill_2 FILLER_55_214 ();
 sg13g2_decap_8 FILLER_55_242 ();
 sg13g2_fill_2 FILLER_55_249 ();
 sg13g2_decap_8 FILLER_55_269 ();
 sg13g2_decap_8 FILLER_55_288 ();
 sg13g2_decap_8 FILLER_55_295 ();
 sg13g2_fill_2 FILLER_55_315 ();
 sg13g2_fill_1 FILLER_55_317 ();
 sg13g2_fill_1 FILLER_55_395 ();
 sg13g2_fill_2 FILLER_55_418 ();
 sg13g2_decap_8 FILLER_55_430 ();
 sg13g2_fill_1 FILLER_55_437 ();
 sg13g2_fill_2 FILLER_55_448 ();
 sg13g2_fill_1 FILLER_55_455 ();
 sg13g2_decap_8 FILLER_55_466 ();
 sg13g2_fill_2 FILLER_55_473 ();
 sg13g2_fill_1 FILLER_55_475 ();
 sg13g2_decap_4 FILLER_55_485 ();
 sg13g2_fill_1 FILLER_55_489 ();
 sg13g2_fill_2 FILLER_55_500 ();
 sg13g2_fill_2 FILLER_55_529 ();
 sg13g2_fill_1 FILLER_55_531 ();
 sg13g2_fill_2 FILLER_55_538 ();
 sg13g2_fill_1 FILLER_55_540 ();
 sg13g2_decap_8 FILLER_55_576 ();
 sg13g2_decap_4 FILLER_55_583 ();
 sg13g2_decap_4 FILLER_55_608 ();
 sg13g2_fill_2 FILLER_55_616 ();
 sg13g2_fill_1 FILLER_55_618 ();
 sg13g2_fill_2 FILLER_55_625 ();
 sg13g2_fill_1 FILLER_55_627 ();
 sg13g2_decap_8 FILLER_55_646 ();
 sg13g2_decap_4 FILLER_55_653 ();
 sg13g2_fill_1 FILLER_55_657 ();
 sg13g2_fill_2 FILLER_55_674 ();
 sg13g2_fill_1 FILLER_55_676 ();
 sg13g2_fill_1 FILLER_55_697 ();
 sg13g2_decap_4 FILLER_55_703 ();
 sg13g2_fill_1 FILLER_55_707 ();
 sg13g2_fill_1 FILLER_55_718 ();
 sg13g2_decap_8 FILLER_55_724 ();
 sg13g2_decap_8 FILLER_55_731 ();
 sg13g2_fill_1 FILLER_55_738 ();
 sg13g2_decap_8 FILLER_55_749 ();
 sg13g2_fill_1 FILLER_55_756 ();
 sg13g2_decap_8 FILLER_55_770 ();
 sg13g2_fill_2 FILLER_55_777 ();
 sg13g2_fill_2 FILLER_55_784 ();
 sg13g2_decap_4 FILLER_55_791 ();
 sg13g2_fill_2 FILLER_55_795 ();
 sg13g2_fill_2 FILLER_55_808 ();
 sg13g2_fill_2 FILLER_55_815 ();
 sg13g2_decap_4 FILLER_55_826 ();
 sg13g2_fill_1 FILLER_55_861 ();
 sg13g2_decap_4 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_4 ();
 sg13g2_fill_1 FILLER_56_37 ();
 sg13g2_fill_2 FILLER_56_58 ();
 sg13g2_fill_2 FILLER_56_70 ();
 sg13g2_fill_1 FILLER_56_72 ();
 sg13g2_fill_1 FILLER_56_103 ();
 sg13g2_fill_2 FILLER_56_164 ();
 sg13g2_fill_1 FILLER_56_166 ();
 sg13g2_decap_4 FILLER_56_177 ();
 sg13g2_fill_1 FILLER_56_191 ();
 sg13g2_decap_4 FILLER_56_197 ();
 sg13g2_fill_2 FILLER_56_201 ();
 sg13g2_fill_2 FILLER_56_210 ();
 sg13g2_decap_8 FILLER_56_243 ();
 sg13g2_fill_2 FILLER_56_254 ();
 sg13g2_fill_1 FILLER_56_256 ();
 sg13g2_decap_4 FILLER_56_262 ();
 sg13g2_fill_1 FILLER_56_266 ();
 sg13g2_fill_2 FILLER_56_317 ();
 sg13g2_decap_8 FILLER_56_359 ();
 sg13g2_decap_8 FILLER_56_366 ();
 sg13g2_decap_4 FILLER_56_373 ();
 sg13g2_decap_4 FILLER_56_385 ();
 sg13g2_decap_8 FILLER_56_393 ();
 sg13g2_decap_4 FILLER_56_403 ();
 sg13g2_fill_1 FILLER_56_407 ();
 sg13g2_decap_8 FILLER_56_425 ();
 sg13g2_fill_1 FILLER_56_432 ();
 sg13g2_fill_2 FILLER_56_451 ();
 sg13g2_fill_1 FILLER_56_453 ();
 sg13g2_fill_2 FILLER_56_472 ();
 sg13g2_decap_8 FILLER_56_503 ();
 sg13g2_fill_2 FILLER_56_510 ();
 sg13g2_fill_1 FILLER_56_512 ();
 sg13g2_decap_8 FILLER_56_522 ();
 sg13g2_fill_1 FILLER_56_529 ();
 sg13g2_fill_1 FILLER_56_534 ();
 sg13g2_fill_2 FILLER_56_541 ();
 sg13g2_decap_8 FILLER_56_553 ();
 sg13g2_decap_8 FILLER_56_568 ();
 sg13g2_fill_2 FILLER_56_575 ();
 sg13g2_fill_1 FILLER_56_577 ();
 sg13g2_fill_1 FILLER_56_582 ();
 sg13g2_decap_8 FILLER_56_602 ();
 sg13g2_fill_2 FILLER_56_609 ();
 sg13g2_fill_2 FILLER_56_617 ();
 sg13g2_fill_1 FILLER_56_619 ();
 sg13g2_decap_8 FILLER_56_625 ();
 sg13g2_decap_8 FILLER_56_632 ();
 sg13g2_decap_8 FILLER_56_649 ();
 sg13g2_fill_1 FILLER_56_656 ();
 sg13g2_fill_1 FILLER_56_669 ();
 sg13g2_decap_8 FILLER_56_675 ();
 sg13g2_decap_8 FILLER_56_682 ();
 sg13g2_fill_2 FILLER_56_706 ();
 sg13g2_decap_4 FILLER_56_715 ();
 sg13g2_fill_1 FILLER_56_737 ();
 sg13g2_decap_8 FILLER_56_748 ();
 sg13g2_fill_2 FILLER_56_755 ();
 sg13g2_fill_1 FILLER_56_757 ();
 sg13g2_decap_8 FILLER_56_766 ();
 sg13g2_fill_2 FILLER_56_773 ();
 sg13g2_fill_2 FILLER_56_793 ();
 sg13g2_fill_2 FILLER_56_814 ();
 sg13g2_fill_2 FILLER_56_830 ();
 sg13g2_fill_1 FILLER_56_832 ();
 sg13g2_decap_8 FILLER_56_852 ();
 sg13g2_fill_2 FILLER_56_859 ();
 sg13g2_fill_1 FILLER_56_861 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_7 ();
 sg13g2_fill_1 FILLER_57_9 ();
 sg13g2_fill_1 FILLER_57_33 ();
 sg13g2_fill_1 FILLER_57_45 ();
 sg13g2_fill_1 FILLER_57_56 ();
 sg13g2_fill_2 FILLER_57_86 ();
 sg13g2_decap_8 FILLER_57_104 ();
 sg13g2_fill_2 FILLER_57_111 ();
 sg13g2_fill_1 FILLER_57_113 ();
 sg13g2_fill_2 FILLER_57_140 ();
 sg13g2_fill_2 FILLER_57_150 ();
 sg13g2_fill_2 FILLER_57_164 ();
 sg13g2_fill_1 FILLER_57_181 ();
 sg13g2_fill_1 FILLER_57_222 ();
 sg13g2_decap_4 FILLER_57_239 ();
 sg13g2_fill_2 FILLER_57_243 ();
 sg13g2_fill_1 FILLER_57_266 ();
 sg13g2_fill_1 FILLER_57_276 ();
 sg13g2_fill_1 FILLER_57_298 ();
 sg13g2_fill_1 FILLER_57_315 ();
 sg13g2_fill_1 FILLER_57_348 ();
 sg13g2_decap_8 FILLER_57_353 ();
 sg13g2_fill_2 FILLER_57_372 ();
 sg13g2_fill_1 FILLER_57_379 ();
 sg13g2_fill_1 FILLER_57_392 ();
 sg13g2_fill_2 FILLER_57_428 ();
 sg13g2_decap_4 FILLER_57_449 ();
 sg13g2_decap_4 FILLER_57_459 ();
 sg13g2_decap_4 FILLER_57_472 ();
 sg13g2_fill_2 FILLER_57_476 ();
 sg13g2_decap_8 FILLER_57_494 ();
 sg13g2_fill_2 FILLER_57_501 ();
 sg13g2_fill_2 FILLER_57_511 ();
 sg13g2_decap_4 FILLER_57_518 ();
 sg13g2_fill_2 FILLER_57_522 ();
 sg13g2_decap_8 FILLER_57_530 ();
 sg13g2_decap_4 FILLER_57_537 ();
 sg13g2_decap_4 FILLER_57_566 ();
 sg13g2_fill_2 FILLER_57_570 ();
 sg13g2_fill_1 FILLER_57_581 ();
 sg13g2_decap_4 FILLER_57_598 ();
 sg13g2_fill_1 FILLER_57_602 ();
 sg13g2_fill_2 FILLER_57_622 ();
 sg13g2_fill_2 FILLER_57_637 ();
 sg13g2_fill_2 FILLER_57_656 ();
 sg13g2_fill_1 FILLER_57_658 ();
 sg13g2_decap_8 FILLER_57_674 ();
 sg13g2_decap_8 FILLER_57_681 ();
 sg13g2_fill_1 FILLER_57_688 ();
 sg13g2_decap_8 FILLER_57_709 ();
 sg13g2_decap_4 FILLER_57_716 ();
 sg13g2_fill_1 FILLER_57_720 ();
 sg13g2_fill_2 FILLER_57_737 ();
 sg13g2_fill_2 FILLER_57_758 ();
 sg13g2_fill_1 FILLER_57_760 ();
 sg13g2_fill_2 FILLER_57_769 ();
 sg13g2_fill_1 FILLER_57_771 ();
 sg13g2_fill_2 FILLER_57_777 ();
 sg13g2_fill_1 FILLER_57_779 ();
 sg13g2_decap_8 FILLER_57_789 ();
 sg13g2_fill_1 FILLER_57_817 ();
 sg13g2_fill_1 FILLER_57_823 ();
 sg13g2_fill_1 FILLER_57_829 ();
 sg13g2_fill_1 FILLER_57_835 ();
 sg13g2_fill_1 FILLER_57_845 ();
 sg13g2_decap_8 FILLER_57_855 ();
 sg13g2_decap_4 FILLER_58_0 ();
 sg13g2_fill_2 FILLER_58_41 ();
 sg13g2_fill_2 FILLER_58_61 ();
 sg13g2_decap_8 FILLER_58_113 ();
 sg13g2_decap_4 FILLER_58_120 ();
 sg13g2_fill_1 FILLER_58_124 ();
 sg13g2_fill_2 FILLER_58_129 ();
 sg13g2_fill_1 FILLER_58_131 ();
 sg13g2_decap_8 FILLER_58_142 ();
 sg13g2_decap_8 FILLER_58_149 ();
 sg13g2_decap_8 FILLER_58_156 ();
 sg13g2_fill_2 FILLER_58_167 ();
 sg13g2_fill_2 FILLER_58_179 ();
 sg13g2_decap_8 FILLER_58_187 ();
 sg13g2_decap_4 FILLER_58_194 ();
 sg13g2_fill_2 FILLER_58_198 ();
 sg13g2_fill_2 FILLER_58_226 ();
 sg13g2_fill_1 FILLER_58_228 ();
 sg13g2_fill_1 FILLER_58_254 ();
 sg13g2_decap_8 FILLER_58_261 ();
 sg13g2_fill_2 FILLER_58_268 ();
 sg13g2_fill_1 FILLER_58_302 ();
 sg13g2_fill_1 FILLER_58_328 ();
 sg13g2_fill_2 FILLER_58_350 ();
 sg13g2_decap_4 FILLER_58_378 ();
 sg13g2_fill_1 FILLER_58_401 ();
 sg13g2_fill_1 FILLER_58_411 ();
 sg13g2_fill_2 FILLER_58_417 ();
 sg13g2_fill_2 FILLER_58_423 ();
 sg13g2_fill_1 FILLER_58_425 ();
 sg13g2_decap_8 FILLER_58_430 ();
 sg13g2_decap_8 FILLER_58_437 ();
 sg13g2_decap_4 FILLER_58_449 ();
 sg13g2_fill_2 FILLER_58_459 ();
 sg13g2_fill_2 FILLER_58_466 ();
 sg13g2_fill_2 FILLER_58_480 ();
 sg13g2_fill_1 FILLER_58_502 ();
 sg13g2_fill_2 FILLER_58_507 ();
 sg13g2_fill_1 FILLER_58_509 ();
 sg13g2_fill_1 FILLER_58_515 ();
 sg13g2_fill_1 FILLER_58_530 ();
 sg13g2_decap_8 FILLER_58_542 ();
 sg13g2_fill_2 FILLER_58_549 ();
 sg13g2_fill_1 FILLER_58_551 ();
 sg13g2_decap_8 FILLER_58_560 ();
 sg13g2_fill_2 FILLER_58_567 ();
 sg13g2_decap_4 FILLER_58_574 ();
 sg13g2_fill_2 FILLER_58_578 ();
 sg13g2_decap_4 FILLER_58_588 ();
 sg13g2_fill_1 FILLER_58_592 ();
 sg13g2_fill_2 FILLER_58_598 ();
 sg13g2_fill_1 FILLER_58_600 ();
 sg13g2_decap_8 FILLER_58_620 ();
 sg13g2_decap_8 FILLER_58_627 ();
 sg13g2_decap_4 FILLER_58_634 ();
 sg13g2_fill_1 FILLER_58_638 ();
 sg13g2_decap_4 FILLER_58_659 ();
 sg13g2_fill_1 FILLER_58_663 ();
 sg13g2_fill_2 FILLER_58_669 ();
 sg13g2_decap_8 FILLER_58_682 ();
 sg13g2_fill_2 FILLER_58_689 ();
 sg13g2_decap_4 FILLER_58_697 ();
 sg13g2_fill_2 FILLER_58_701 ();
 sg13g2_decap_8 FILLER_58_708 ();
 sg13g2_fill_1 FILLER_58_715 ();
 sg13g2_decap_4 FILLER_58_731 ();
 sg13g2_decap_4 FILLER_58_744 ();
 sg13g2_fill_2 FILLER_58_771 ();
 sg13g2_fill_1 FILLER_58_773 ();
 sg13g2_decap_4 FILLER_58_782 ();
 sg13g2_fill_1 FILLER_58_792 ();
 sg13g2_decap_8 FILLER_58_806 ();
 sg13g2_decap_4 FILLER_58_813 ();
 sg13g2_fill_2 FILLER_58_817 ();
 sg13g2_fill_2 FILLER_58_825 ();
 sg13g2_fill_1 FILLER_58_827 ();
 sg13g2_decap_4 FILLER_58_858 ();
 sg13g2_fill_2 FILLER_59_61 ();
 sg13g2_fill_2 FILLER_59_95 ();
 sg13g2_fill_1 FILLER_59_97 ();
 sg13g2_fill_1 FILLER_59_224 ();
 sg13g2_fill_2 FILLER_59_231 ();
 sg13g2_fill_2 FILLER_59_261 ();
 sg13g2_fill_1 FILLER_59_263 ();
 sg13g2_fill_2 FILLER_59_273 ();
 sg13g2_fill_2 FILLER_59_343 ();
 sg13g2_fill_2 FILLER_59_364 ();
 sg13g2_fill_1 FILLER_59_397 ();
 sg13g2_decap_8 FILLER_59_411 ();
 sg13g2_fill_2 FILLER_59_418 ();
 sg13g2_fill_1 FILLER_59_439 ();
 sg13g2_decap_8 FILLER_59_450 ();
 sg13g2_fill_2 FILLER_59_457 ();
 sg13g2_fill_2 FILLER_59_474 ();
 sg13g2_fill_1 FILLER_59_476 ();
 sg13g2_fill_1 FILLER_59_482 ();
 sg13g2_decap_8 FILLER_59_493 ();
 sg13g2_fill_2 FILLER_59_500 ();
 sg13g2_fill_1 FILLER_59_502 ();
 sg13g2_fill_2 FILLER_59_511 ();
 sg13g2_decap_8 FILLER_59_523 ();
 sg13g2_decap_4 FILLER_59_530 ();
 sg13g2_fill_1 FILLER_59_534 ();
 sg13g2_decap_4 FILLER_59_551 ();
 sg13g2_fill_2 FILLER_59_606 ();
 sg13g2_fill_1 FILLER_59_608 ();
 sg13g2_decap_4 FILLER_59_614 ();
 sg13g2_fill_1 FILLER_59_618 ();
 sg13g2_decap_8 FILLER_59_628 ();
 sg13g2_decap_4 FILLER_59_640 ();
 sg13g2_decap_4 FILLER_59_649 ();
 sg13g2_fill_1 FILLER_59_653 ();
 sg13g2_decap_8 FILLER_59_670 ();
 sg13g2_fill_2 FILLER_59_683 ();
 sg13g2_fill_2 FILLER_59_705 ();
 sg13g2_fill_1 FILLER_59_711 ();
 sg13g2_decap_4 FILLER_59_716 ();
 sg13g2_fill_2 FILLER_59_732 ();
 sg13g2_decap_8 FILLER_59_740 ();
 sg13g2_decap_4 FILLER_59_747 ();
 sg13g2_fill_1 FILLER_59_751 ();
 sg13g2_decap_8 FILLER_59_759 ();
 sg13g2_decap_8 FILLER_59_766 ();
 sg13g2_fill_2 FILLER_59_791 ();
 sg13g2_fill_1 FILLER_59_793 ();
 sg13g2_decap_8 FILLER_59_798 ();
 sg13g2_decap_8 FILLER_59_818 ();
 sg13g2_fill_2 FILLER_59_825 ();
 sg13g2_decap_8 FILLER_59_836 ();
 sg13g2_decap_4 FILLER_59_843 ();
 sg13g2_fill_2 FILLER_59_847 ();
 sg13g2_decap_4 FILLER_59_857 ();
 sg13g2_fill_1 FILLER_59_861 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_7 ();
 sg13g2_fill_1 FILLER_60_9 ();
 sg13g2_fill_2 FILLER_60_21 ();
 sg13g2_fill_2 FILLER_60_38 ();
 sg13g2_fill_1 FILLER_60_40 ();
 sg13g2_fill_2 FILLER_60_63 ();
 sg13g2_decap_4 FILLER_60_87 ();
 sg13g2_fill_2 FILLER_60_108 ();
 sg13g2_fill_1 FILLER_60_110 ();
 sg13g2_decap_8 FILLER_60_125 ();
 sg13g2_fill_2 FILLER_60_132 ();
 sg13g2_fill_1 FILLER_60_134 ();
 sg13g2_decap_8 FILLER_60_147 ();
 sg13g2_decap_4 FILLER_60_180 ();
 sg13g2_fill_2 FILLER_60_184 ();
 sg13g2_fill_2 FILLER_60_191 ();
 sg13g2_decap_8 FILLER_60_325 ();
 sg13g2_decap_8 FILLER_60_332 ();
 sg13g2_fill_1 FILLER_60_339 ();
 sg13g2_decap_4 FILLER_60_362 ();
 sg13g2_fill_2 FILLER_60_375 ();
 sg13g2_fill_2 FILLER_60_393 ();
 sg13g2_decap_4 FILLER_60_414 ();
 sg13g2_decap_4 FILLER_60_431 ();
 sg13g2_fill_2 FILLER_60_435 ();
 sg13g2_fill_2 FILLER_60_450 ();
 sg13g2_fill_1 FILLER_60_452 ();
 sg13g2_decap_8 FILLER_60_471 ();
 sg13g2_fill_2 FILLER_60_478 ();
 sg13g2_fill_1 FILLER_60_480 ();
 sg13g2_decap_8 FILLER_60_487 ();
 sg13g2_fill_1 FILLER_60_494 ();
 sg13g2_fill_2 FILLER_60_501 ();
 sg13g2_fill_1 FILLER_60_513 ();
 sg13g2_fill_1 FILLER_60_524 ();
 sg13g2_decap_4 FILLER_60_539 ();
 sg13g2_fill_2 FILLER_60_543 ();
 sg13g2_decap_4 FILLER_60_550 ();
 sg13g2_fill_2 FILLER_60_554 ();
 sg13g2_fill_1 FILLER_60_576 ();
 sg13g2_decap_4 FILLER_60_583 ();
 sg13g2_fill_1 FILLER_60_587 ();
 sg13g2_fill_1 FILLER_60_601 ();
 sg13g2_fill_2 FILLER_60_615 ();
 sg13g2_fill_1 FILLER_60_617 ();
 sg13g2_fill_1 FILLER_60_629 ();
 sg13g2_fill_1 FILLER_60_636 ();
 sg13g2_fill_2 FILLER_60_646 ();
 sg13g2_fill_1 FILLER_60_648 ();
 sg13g2_decap_4 FILLER_60_654 ();
 sg13g2_decap_8 FILLER_60_676 ();
 sg13g2_fill_1 FILLER_60_688 ();
 sg13g2_decap_8 FILLER_60_704 ();
 sg13g2_decap_4 FILLER_60_711 ();
 sg13g2_fill_2 FILLER_60_715 ();
 sg13g2_fill_1 FILLER_60_727 ();
 sg13g2_decap_4 FILLER_60_734 ();
 sg13g2_decap_8 FILLER_60_743 ();
 sg13g2_fill_2 FILLER_60_750 ();
 sg13g2_fill_2 FILLER_60_757 ();
 sg13g2_fill_1 FILLER_60_759 ();
 sg13g2_decap_4 FILLER_60_784 ();
 sg13g2_fill_1 FILLER_60_788 ();
 sg13g2_decap_4 FILLER_60_793 ();
 sg13g2_fill_1 FILLER_60_797 ();
 sg13g2_decap_4 FILLER_60_816 ();
 sg13g2_fill_2 FILLER_60_820 ();
 sg13g2_fill_2 FILLER_60_826 ();
 sg13g2_fill_2 FILLER_60_848 ();
 sg13g2_decap_8 FILLER_60_855 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_4 FILLER_61_29 ();
 sg13g2_fill_1 FILLER_61_33 ();
 sg13g2_fill_2 FILLER_61_45 ();
 sg13g2_fill_1 FILLER_61_47 ();
 sg13g2_decap_8 FILLER_61_64 ();
 sg13g2_decap_4 FILLER_61_71 ();
 sg13g2_fill_2 FILLER_61_75 ();
 sg13g2_fill_1 FILLER_61_91 ();
 sg13g2_decap_4 FILLER_61_98 ();
 sg13g2_fill_2 FILLER_61_102 ();
 sg13g2_decap_8 FILLER_61_123 ();
 sg13g2_fill_2 FILLER_61_130 ();
 sg13g2_fill_1 FILLER_61_132 ();
 sg13g2_decap_8 FILLER_61_153 ();
 sg13g2_decap_4 FILLER_61_160 ();
 sg13g2_fill_2 FILLER_61_164 ();
 sg13g2_fill_2 FILLER_61_174 ();
 sg13g2_fill_1 FILLER_61_176 ();
 sg13g2_fill_1 FILLER_61_249 ();
 sg13g2_fill_1 FILLER_61_259 ();
 sg13g2_fill_1 FILLER_61_278 ();
 sg13g2_fill_1 FILLER_61_288 ();
 sg13g2_fill_2 FILLER_61_304 ();
 sg13g2_fill_1 FILLER_61_315 ();
 sg13g2_fill_2 FILLER_61_322 ();
 sg13g2_fill_2 FILLER_61_339 ();
 sg13g2_fill_1 FILLER_61_341 ();
 sg13g2_decap_4 FILLER_61_350 ();
 sg13g2_decap_4 FILLER_61_364 ();
 sg13g2_fill_2 FILLER_61_393 ();
 sg13g2_fill_1 FILLER_61_404 ();
 sg13g2_decap_8 FILLER_61_410 ();
 sg13g2_decap_8 FILLER_61_417 ();
 sg13g2_decap_8 FILLER_61_424 ();
 sg13g2_decap_4 FILLER_61_431 ();
 sg13g2_decap_8 FILLER_61_450 ();
 sg13g2_fill_1 FILLER_61_457 ();
 sg13g2_fill_2 FILLER_61_472 ();
 sg13g2_fill_1 FILLER_61_474 ();
 sg13g2_fill_2 FILLER_61_481 ();
 sg13g2_fill_2 FILLER_61_503 ();
 sg13g2_fill_1 FILLER_61_505 ();
 sg13g2_fill_1 FILLER_61_514 ();
 sg13g2_decap_8 FILLER_61_520 ();
 sg13g2_decap_8 FILLER_61_527 ();
 sg13g2_decap_8 FILLER_61_534 ();
 sg13g2_decap_4 FILLER_61_541 ();
 sg13g2_fill_2 FILLER_61_557 ();
 sg13g2_decap_4 FILLER_61_565 ();
 sg13g2_fill_2 FILLER_61_569 ();
 sg13g2_decap_8 FILLER_61_577 ();
 sg13g2_decap_4 FILLER_61_584 ();
 sg13g2_decap_4 FILLER_61_603 ();
 sg13g2_fill_2 FILLER_61_615 ();
 sg13g2_decap_8 FILLER_61_628 ();
 sg13g2_decap_8 FILLER_61_635 ();
 sg13g2_fill_1 FILLER_61_642 ();
 sg13g2_fill_1 FILLER_61_648 ();
 sg13g2_fill_2 FILLER_61_658 ();
 sg13g2_fill_1 FILLER_61_660 ();
 sg13g2_decap_4 FILLER_61_666 ();
 sg13g2_fill_2 FILLER_61_670 ();
 sg13g2_fill_2 FILLER_61_700 ();
 sg13g2_decap_4 FILLER_61_712 ();
 sg13g2_decap_4 FILLER_61_737 ();
 sg13g2_fill_1 FILLER_61_741 ();
 sg13g2_decap_8 FILLER_61_764 ();
 sg13g2_decap_4 FILLER_61_771 ();
 sg13g2_fill_2 FILLER_61_780 ();
 sg13g2_fill_2 FILLER_61_801 ();
 sg13g2_fill_1 FILLER_61_803 ();
 sg13g2_fill_2 FILLER_61_810 ();
 sg13g2_fill_1 FILLER_61_812 ();
 sg13g2_decap_8 FILLER_61_819 ();
 sg13g2_fill_2 FILLER_61_826 ();
 sg13g2_decap_8 FILLER_61_852 ();
 sg13g2_fill_2 FILLER_61_859 ();
 sg13g2_fill_1 FILLER_61_861 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_4 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_29 ();
 sg13g2_decap_8 FILLER_62_36 ();
 sg13g2_decap_8 FILLER_62_43 ();
 sg13g2_fill_2 FILLER_62_63 ();
 sg13g2_fill_1 FILLER_62_65 ();
 sg13g2_decap_4 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_91 ();
 sg13g2_fill_1 FILLER_62_98 ();
 sg13g2_fill_2 FILLER_62_107 ();
 sg13g2_fill_1 FILLER_62_109 ();
 sg13g2_decap_8 FILLER_62_114 ();
 sg13g2_decap_8 FILLER_62_121 ();
 sg13g2_fill_2 FILLER_62_128 ();
 sg13g2_decap_8 FILLER_62_138 ();
 sg13g2_fill_2 FILLER_62_145 ();
 sg13g2_decap_8 FILLER_62_181 ();
 sg13g2_decap_4 FILLER_62_188 ();
 sg13g2_fill_1 FILLER_62_192 ();
 sg13g2_decap_8 FILLER_62_197 ();
 sg13g2_decap_4 FILLER_62_204 ();
 sg13g2_fill_1 FILLER_62_208 ();
 sg13g2_fill_1 FILLER_62_213 ();
 sg13g2_fill_2 FILLER_62_255 ();
 sg13g2_fill_1 FILLER_62_283 ();
 sg13g2_decap_4 FILLER_62_336 ();
 sg13g2_fill_1 FILLER_62_340 ();
 sg13g2_fill_2 FILLER_62_346 ();
 sg13g2_fill_1 FILLER_62_348 ();
 sg13g2_fill_1 FILLER_62_380 ();
 sg13g2_decap_8 FILLER_62_391 ();
 sg13g2_decap_8 FILLER_62_398 ();
 sg13g2_decap_4 FILLER_62_422 ();
 sg13g2_fill_2 FILLER_62_426 ();
 sg13g2_fill_2 FILLER_62_442 ();
 sg13g2_fill_1 FILLER_62_444 ();
 sg13g2_fill_2 FILLER_62_450 ();
 sg13g2_fill_1 FILLER_62_460 ();
 sg13g2_decap_8 FILLER_62_466 ();
 sg13g2_decap_8 FILLER_62_473 ();
 sg13g2_decap_4 FILLER_62_480 ();
 sg13g2_fill_1 FILLER_62_484 ();
 sg13g2_decap_8 FILLER_62_491 ();
 sg13g2_fill_1 FILLER_62_498 ();
 sg13g2_fill_2 FILLER_62_508 ();
 sg13g2_fill_1 FILLER_62_526 ();
 sg13g2_fill_2 FILLER_62_549 ();
 sg13g2_fill_1 FILLER_62_551 ();
 sg13g2_fill_1 FILLER_62_563 ();
 sg13g2_decap_4 FILLER_62_586 ();
 sg13g2_fill_2 FILLER_62_603 ();
 sg13g2_fill_1 FILLER_62_605 ();
 sg13g2_fill_2 FILLER_62_613 ();
 sg13g2_decap_4 FILLER_62_626 ();
 sg13g2_fill_2 FILLER_62_630 ();
 sg13g2_decap_4 FILLER_62_636 ();
 sg13g2_fill_2 FILLER_62_640 ();
 sg13g2_decap_4 FILLER_62_656 ();
 sg13g2_fill_2 FILLER_62_660 ();
 sg13g2_fill_2 FILLER_62_668 ();
 sg13g2_fill_1 FILLER_62_670 ();
 sg13g2_decap_8 FILLER_62_680 ();
 sg13g2_decap_4 FILLER_62_687 ();
 sg13g2_decap_8 FILLER_62_696 ();
 sg13g2_decap_4 FILLER_62_715 ();
 sg13g2_fill_2 FILLER_62_719 ();
 sg13g2_decap_8 FILLER_62_736 ();
 sg13g2_fill_2 FILLER_62_743 ();
 sg13g2_fill_2 FILLER_62_750 ();
 sg13g2_fill_1 FILLER_62_752 ();
 sg13g2_decap_8 FILLER_62_759 ();
 sg13g2_fill_2 FILLER_62_766 ();
 sg13g2_decap_8 FILLER_62_789 ();
 sg13g2_decap_4 FILLER_62_796 ();
 sg13g2_fill_2 FILLER_62_800 ();
 sg13g2_fill_1 FILLER_62_849 ();
 sg13g2_decap_4 FILLER_62_858 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_4 FILLER_63_7 ();
 sg13g2_fill_2 FILLER_63_11 ();
 sg13g2_decap_4 FILLER_63_28 ();
 sg13g2_fill_2 FILLER_63_32 ();
 sg13g2_decap_8 FILLER_63_39 ();
 sg13g2_decap_4 FILLER_63_63 ();
 sg13g2_fill_1 FILLER_63_67 ();
 sg13g2_fill_2 FILLER_63_93 ();
 sg13g2_fill_2 FILLER_63_115 ();
 sg13g2_fill_1 FILLER_63_117 ();
 sg13g2_decap_8 FILLER_63_146 ();
 sg13g2_decap_4 FILLER_63_153 ();
 sg13g2_fill_1 FILLER_63_170 ();
 sg13g2_fill_1 FILLER_63_181 ();
 sg13g2_fill_2 FILLER_63_213 ();
 sg13g2_decap_8 FILLER_63_218 ();
 sg13g2_decap_4 FILLER_63_225 ();
 sg13g2_fill_2 FILLER_63_236 ();
 sg13g2_fill_2 FILLER_63_259 ();
 sg13g2_fill_2 FILLER_63_307 ();
 sg13g2_fill_1 FILLER_63_309 ();
 sg13g2_fill_2 FILLER_63_362 ();
 sg13g2_fill_1 FILLER_63_364 ();
 sg13g2_decap_8 FILLER_63_369 ();
 sg13g2_fill_1 FILLER_63_376 ();
 sg13g2_decap_4 FILLER_63_381 ();
 sg13g2_fill_1 FILLER_63_385 ();
 sg13g2_decap_8 FILLER_63_412 ();
 sg13g2_decap_8 FILLER_63_419 ();
 sg13g2_decap_4 FILLER_63_426 ();
 sg13g2_decap_8 FILLER_63_450 ();
 sg13g2_decap_8 FILLER_63_501 ();
 sg13g2_fill_1 FILLER_63_508 ();
 sg13g2_fill_2 FILLER_63_523 ();
 sg13g2_fill_1 FILLER_63_525 ();
 sg13g2_decap_4 FILLER_63_532 ();
 sg13g2_fill_2 FILLER_63_547 ();
 sg13g2_fill_1 FILLER_63_549 ();
 sg13g2_decap_4 FILLER_63_559 ();
 sg13g2_fill_1 FILLER_63_569 ();
 sg13g2_decap_8 FILLER_63_575 ();
 sg13g2_fill_2 FILLER_63_582 ();
 sg13g2_fill_1 FILLER_63_584 ();
 sg13g2_decap_4 FILLER_63_598 ();
 sg13g2_fill_2 FILLER_63_602 ();
 sg13g2_decap_8 FILLER_63_630 ();
 sg13g2_decap_8 FILLER_63_657 ();
 sg13g2_fill_2 FILLER_63_664 ();
 sg13g2_fill_1 FILLER_63_666 ();
 sg13g2_decap_4 FILLER_63_684 ();
 sg13g2_decap_8 FILLER_63_711 ();
 sg13g2_decap_8 FILLER_63_718 ();
 sg13g2_fill_2 FILLER_63_730 ();
 sg13g2_fill_1 FILLER_63_732 ();
 sg13g2_fill_1 FILLER_63_768 ();
 sg13g2_decap_4 FILLER_63_791 ();
 sg13g2_fill_2 FILLER_63_795 ();
 sg13g2_decap_8 FILLER_63_813 ();
 sg13g2_decap_4 FILLER_63_820 ();
 sg13g2_fill_1 FILLER_63_824 ();
 sg13g2_fill_2 FILLER_63_842 ();
 sg13g2_fill_1 FILLER_63_844 ();
 sg13g2_decap_4 FILLER_63_858 ();
 sg13g2_fill_2 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_fill_2 FILLER_64_42 ();
 sg13g2_fill_1 FILLER_64_44 ();
 sg13g2_decap_4 FILLER_64_65 ();
 sg13g2_fill_1 FILLER_64_69 ();
 sg13g2_fill_2 FILLER_64_75 ();
 sg13g2_fill_2 FILLER_64_83 ();
 sg13g2_decap_4 FILLER_64_90 ();
 sg13g2_fill_2 FILLER_64_117 ();
 sg13g2_fill_1 FILLER_64_119 ();
 sg13g2_decap_8 FILLER_64_135 ();
 sg13g2_fill_2 FILLER_64_173 ();
 sg13g2_fill_2 FILLER_64_185 ();
 sg13g2_fill_2 FILLER_64_196 ();
 sg13g2_decap_8 FILLER_64_202 ();
 sg13g2_fill_2 FILLER_64_209 ();
 sg13g2_fill_2 FILLER_64_219 ();
 sg13g2_fill_1 FILLER_64_247 ();
 sg13g2_decap_4 FILLER_64_253 ();
 sg13g2_fill_1 FILLER_64_257 ();
 sg13g2_fill_1 FILLER_64_265 ();
 sg13g2_decap_4 FILLER_64_303 ();
 sg13g2_fill_1 FILLER_64_307 ();
 sg13g2_fill_1 FILLER_64_340 ();
 sg13g2_fill_1 FILLER_64_346 ();
 sg13g2_decap_8 FILLER_64_351 ();
 sg13g2_decap_8 FILLER_64_358 ();
 sg13g2_decap_8 FILLER_64_424 ();
 sg13g2_fill_1 FILLER_64_431 ();
 sg13g2_fill_2 FILLER_64_457 ();
 sg13g2_decap_8 FILLER_64_475 ();
 sg13g2_decap_8 FILLER_64_496 ();
 sg13g2_fill_2 FILLER_64_503 ();
 sg13g2_fill_1 FILLER_64_505 ();
 sg13g2_fill_2 FILLER_64_524 ();
 sg13g2_decap_8 FILLER_64_536 ();
 sg13g2_fill_2 FILLER_64_558 ();
 sg13g2_fill_1 FILLER_64_560 ();
 sg13g2_decap_8 FILLER_64_577 ();
 sg13g2_fill_2 FILLER_64_584 ();
 sg13g2_fill_1 FILLER_64_586 ();
 sg13g2_decap_4 FILLER_64_608 ();
 sg13g2_fill_1 FILLER_64_612 ();
 sg13g2_fill_2 FILLER_64_618 ();
 sg13g2_decap_8 FILLER_64_623 ();
 sg13g2_decap_4 FILLER_64_636 ();
 sg13g2_decap_8 FILLER_64_650 ();
 sg13g2_decap_4 FILLER_64_657 ();
 sg13g2_decap_8 FILLER_64_679 ();
 sg13g2_decap_8 FILLER_64_686 ();
 sg13g2_fill_1 FILLER_64_693 ();
 sg13g2_decap_8 FILLER_64_702 ();
 sg13g2_fill_2 FILLER_64_709 ();
 sg13g2_fill_1 FILLER_64_711 ();
 sg13g2_fill_2 FILLER_64_742 ();
 sg13g2_fill_1 FILLER_64_744 ();
 sg13g2_fill_2 FILLER_64_767 ();
 sg13g2_decap_8 FILLER_64_779 ();
 sg13g2_decap_4 FILLER_64_786 ();
 sg13g2_decap_4 FILLER_64_795 ();
 sg13g2_decap_8 FILLER_64_819 ();
 sg13g2_decap_4 FILLER_64_826 ();
 sg13g2_decap_8 FILLER_64_847 ();
 sg13g2_decap_8 FILLER_64_854 ();
 sg13g2_fill_1 FILLER_64_861 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_4 FILLER_65_7 ();
 sg13g2_fill_1 FILLER_65_11 ();
 sg13g2_decap_8 FILLER_65_37 ();
 sg13g2_decap_4 FILLER_65_64 ();
 sg13g2_fill_2 FILLER_65_68 ();
 sg13g2_decap_8 FILLER_65_90 ();
 sg13g2_fill_1 FILLER_65_101 ();
 sg13g2_decap_8 FILLER_65_113 ();
 sg13g2_decap_8 FILLER_65_120 ();
 sg13g2_decap_8 FILLER_65_141 ();
 sg13g2_decap_4 FILLER_65_148 ();
 sg13g2_fill_1 FILLER_65_157 ();
 sg13g2_decap_4 FILLER_65_162 ();
 sg13g2_fill_1 FILLER_65_166 ();
 sg13g2_fill_2 FILLER_65_176 ();
 sg13g2_decap_4 FILLER_65_186 ();
 sg13g2_decap_8 FILLER_65_194 ();
 sg13g2_decap_8 FILLER_65_201 ();
 sg13g2_fill_2 FILLER_65_208 ();
 sg13g2_fill_1 FILLER_65_210 ();
 sg13g2_fill_2 FILLER_65_237 ();
 sg13g2_fill_1 FILLER_65_239 ();
 sg13g2_decap_8 FILLER_65_244 ();
 sg13g2_decap_4 FILLER_65_251 ();
 sg13g2_fill_1 FILLER_65_255 ();
 sg13g2_fill_1 FILLER_65_292 ();
 sg13g2_decap_4 FILLER_65_335 ();
 sg13g2_decap_4 FILLER_65_370 ();
 sg13g2_fill_2 FILLER_65_383 ();
 sg13g2_fill_2 FILLER_65_394 ();
 sg13g2_fill_1 FILLER_65_401 ();
 sg13g2_decap_4 FILLER_65_417 ();
 sg13g2_decap_8 FILLER_65_429 ();
 sg13g2_decap_8 FILLER_65_436 ();
 sg13g2_fill_2 FILLER_65_443 ();
 sg13g2_fill_1 FILLER_65_445 ();
 sg13g2_fill_2 FILLER_65_451 ();
 sg13g2_fill_1 FILLER_65_453 ();
 sg13g2_decap_8 FILLER_65_468 ();
 sg13g2_decap_8 FILLER_65_475 ();
 sg13g2_fill_1 FILLER_65_486 ();
 sg13g2_decap_8 FILLER_65_497 ();
 sg13g2_fill_2 FILLER_65_504 ();
 sg13g2_decap_8 FILLER_65_519 ();
 sg13g2_decap_8 FILLER_65_526 ();
 sg13g2_decap_8 FILLER_65_541 ();
 sg13g2_decap_8 FILLER_65_548 ();
 sg13g2_fill_1 FILLER_65_555 ();
 sg13g2_decap_8 FILLER_65_575 ();
 sg13g2_fill_1 FILLER_65_582 ();
 sg13g2_fill_2 FILLER_65_588 ();
 sg13g2_fill_1 FILLER_65_590 ();
 sg13g2_decap_8 FILLER_65_601 ();
 sg13g2_decap_8 FILLER_65_608 ();
 sg13g2_fill_1 FILLER_65_615 ();
 sg13g2_decap_4 FILLER_65_632 ();
 sg13g2_fill_1 FILLER_65_641 ();
 sg13g2_decap_4 FILLER_65_664 ();
 sg13g2_fill_2 FILLER_65_673 ();
 sg13g2_fill_2 FILLER_65_693 ();
 sg13g2_fill_1 FILLER_65_701 ();
 sg13g2_fill_1 FILLER_65_712 ();
 sg13g2_decap_8 FILLER_65_719 ();
 sg13g2_decap_8 FILLER_65_739 ();
 sg13g2_fill_2 FILLER_65_746 ();
 sg13g2_fill_1 FILLER_65_748 ();
 sg13g2_fill_1 FILLER_65_768 ();
 sg13g2_fill_2 FILLER_65_773 ();
 sg13g2_decap_4 FILLER_65_780 ();
 sg13g2_fill_2 FILLER_65_784 ();
 sg13g2_decap_8 FILLER_65_799 ();
 sg13g2_fill_2 FILLER_65_811 ();
 sg13g2_fill_1 FILLER_65_813 ();
 sg13g2_decap_8 FILLER_65_855 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_4 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_54 ();
 sg13g2_decap_8 FILLER_66_61 ();
 sg13g2_decap_8 FILLER_66_68 ();
 sg13g2_decap_4 FILLER_66_75 ();
 sg13g2_decap_8 FILLER_66_99 ();
 sg13g2_decap_4 FILLER_66_106 ();
 sg13g2_fill_2 FILLER_66_110 ();
 sg13g2_decap_4 FILLER_66_149 ();
 sg13g2_fill_2 FILLER_66_153 ();
 sg13g2_decap_4 FILLER_66_163 ();
 sg13g2_fill_2 FILLER_66_167 ();
 sg13g2_fill_2 FILLER_66_226 ();
 sg13g2_fill_1 FILLER_66_228 ();
 sg13g2_fill_2 FILLER_66_255 ();
 sg13g2_fill_1 FILLER_66_257 ();
 sg13g2_fill_1 FILLER_66_284 ();
 sg13g2_fill_2 FILLER_66_332 ();
 sg13g2_fill_1 FILLER_66_334 ();
 sg13g2_fill_2 FILLER_66_341 ();
 sg13g2_fill_2 FILLER_66_353 ();
 sg13g2_fill_1 FILLER_66_355 ();
 sg13g2_decap_8 FILLER_66_361 ();
 sg13g2_decap_4 FILLER_66_368 ();
 sg13g2_fill_1 FILLER_66_372 ();
 sg13g2_fill_2 FILLER_66_406 ();
 sg13g2_fill_1 FILLER_66_408 ();
 sg13g2_fill_2 FILLER_66_418 ();
 sg13g2_fill_1 FILLER_66_420 ();
 sg13g2_fill_1 FILLER_66_434 ();
 sg13g2_fill_2 FILLER_66_440 ();
 sg13g2_fill_1 FILLER_66_442 ();
 sg13g2_fill_2 FILLER_66_463 ();
 sg13g2_fill_1 FILLER_66_465 ();
 sg13g2_decap_8 FILLER_66_472 ();
 sg13g2_fill_2 FILLER_66_479 ();
 sg13g2_decap_4 FILLER_66_499 ();
 sg13g2_decap_4 FILLER_66_515 ();
 sg13g2_fill_1 FILLER_66_519 ();
 sg13g2_fill_1 FILLER_66_525 ();
 sg13g2_decap_8 FILLER_66_567 ();
 sg13g2_fill_1 FILLER_66_574 ();
 sg13g2_fill_1 FILLER_66_585 ();
 sg13g2_decap_8 FILLER_66_591 ();
 sg13g2_fill_2 FILLER_66_608 ();
 sg13g2_decap_4 FILLER_66_630 ();
 sg13g2_fill_1 FILLER_66_634 ();
 sg13g2_decap_8 FILLER_66_643 ();
 sg13g2_decap_4 FILLER_66_650 ();
 sg13g2_fill_1 FILLER_66_654 ();
 sg13g2_decap_8 FILLER_66_660 ();
 sg13g2_fill_2 FILLER_66_667 ();
 sg13g2_fill_1 FILLER_66_669 ();
 sg13g2_fill_1 FILLER_66_674 ();
 sg13g2_fill_2 FILLER_66_682 ();
 sg13g2_fill_1 FILLER_66_684 ();
 sg13g2_decap_8 FILLER_66_707 ();
 sg13g2_decap_8 FILLER_66_714 ();
 sg13g2_fill_1 FILLER_66_748 ();
 sg13g2_fill_2 FILLER_66_757 ();
 sg13g2_decap_8 FILLER_66_770 ();
 sg13g2_decap_4 FILLER_66_777 ();
 sg13g2_fill_2 FILLER_66_781 ();
 sg13g2_decap_8 FILLER_66_808 ();
 sg13g2_fill_1 FILLER_66_815 ();
 sg13g2_decap_4 FILLER_66_822 ();
 sg13g2_fill_2 FILLER_66_830 ();
 sg13g2_fill_1 FILLER_66_832 ();
 sg13g2_decap_4 FILLER_66_856 ();
 sg13g2_fill_2 FILLER_66_860 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_4 FILLER_67_7 ();
 sg13g2_decap_4 FILLER_67_37 ();
 sg13g2_fill_2 FILLER_67_41 ();
 sg13g2_decap_8 FILLER_67_59 ();
 sg13g2_decap_4 FILLER_67_66 ();
 sg13g2_fill_2 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_4 FILLER_67_89 ();
 sg13g2_fill_1 FILLER_67_93 ();
 sg13g2_decap_4 FILLER_67_100 ();
 sg13g2_fill_1 FILLER_67_104 ();
 sg13g2_fill_2 FILLER_67_110 ();
 sg13g2_fill_1 FILLER_67_112 ();
 sg13g2_fill_2 FILLER_67_126 ();
 sg13g2_fill_1 FILLER_67_128 ();
 sg13g2_decap_8 FILLER_67_141 ();
 sg13g2_decap_8 FILLER_67_148 ();
 sg13g2_decap_4 FILLER_67_155 ();
 sg13g2_fill_1 FILLER_67_184 ();
 sg13g2_fill_2 FILLER_67_211 ();
 sg13g2_decap_8 FILLER_67_239 ();
 sg13g2_decap_4 FILLER_67_246 ();
 sg13g2_fill_2 FILLER_67_284 ();
 sg13g2_fill_1 FILLER_67_286 ();
 sg13g2_decap_4 FILLER_67_332 ();
 sg13g2_fill_2 FILLER_67_352 ();
 sg13g2_decap_8 FILLER_67_385 ();
 sg13g2_fill_2 FILLER_67_392 ();
 sg13g2_decap_8 FILLER_67_403 ();
 sg13g2_decap_8 FILLER_67_410 ();
 sg13g2_fill_1 FILLER_67_417 ();
 sg13g2_fill_2 FILLER_67_441 ();
 sg13g2_fill_1 FILLER_67_443 ();
 sg13g2_fill_2 FILLER_67_453 ();
 sg13g2_fill_1 FILLER_67_455 ();
 sg13g2_fill_2 FILLER_67_466 ();
 sg13g2_fill_1 FILLER_67_504 ();
 sg13g2_fill_2 FILLER_67_537 ();
 sg13g2_fill_1 FILLER_67_544 ();
 sg13g2_decap_8 FILLER_67_552 ();
 sg13g2_fill_2 FILLER_67_559 ();
 sg13g2_fill_1 FILLER_67_561 ();
 sg13g2_fill_2 FILLER_67_572 ();
 sg13g2_fill_2 FILLER_67_578 ();
 sg13g2_fill_1 FILLER_67_580 ();
 sg13g2_fill_2 FILLER_67_608 ();
 sg13g2_fill_1 FILLER_67_610 ();
 sg13g2_fill_1 FILLER_67_625 ();
 sg13g2_decap_4 FILLER_67_632 ();
 sg13g2_fill_1 FILLER_67_661 ();
 sg13g2_decap_4 FILLER_67_681 ();
 sg13g2_fill_2 FILLER_67_685 ();
 sg13g2_fill_1 FILLER_67_697 ();
 sg13g2_fill_2 FILLER_67_704 ();
 sg13g2_decap_8 FILLER_67_714 ();
 sg13g2_decap_4 FILLER_67_721 ();
 sg13g2_fill_1 FILLER_67_725 ();
 sg13g2_fill_2 FILLER_67_731 ();
 sg13g2_fill_1 FILLER_67_733 ();
 sg13g2_decap_8 FILLER_67_742 ();
 sg13g2_fill_2 FILLER_67_765 ();
 sg13g2_fill_1 FILLER_67_767 ();
 sg13g2_decap_8 FILLER_67_785 ();
 sg13g2_fill_1 FILLER_67_792 ();
 sg13g2_decap_8 FILLER_67_809 ();
 sg13g2_fill_2 FILLER_67_831 ();
 sg13g2_fill_1 FILLER_67_833 ();
 sg13g2_fill_2 FILLER_67_859 ();
 sg13g2_fill_1 FILLER_67_861 ();
 sg13g2_decap_4 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_4 ();
 sg13g2_fill_2 FILLER_68_37 ();
 sg13g2_fill_1 FILLER_68_39 ();
 sg13g2_decap_4 FILLER_68_99 ();
 sg13g2_fill_1 FILLER_68_119 ();
 sg13g2_fill_2 FILLER_68_129 ();
 sg13g2_fill_1 FILLER_68_131 ();
 sg13g2_decap_8 FILLER_68_140 ();
 sg13g2_decap_4 FILLER_68_147 ();
 sg13g2_fill_1 FILLER_68_195 ();
 sg13g2_decap_8 FILLER_68_200 ();
 sg13g2_decap_8 FILLER_68_207 ();
 sg13g2_decap_8 FILLER_68_214 ();
 sg13g2_fill_2 FILLER_68_298 ();
 sg13g2_decap_8 FILLER_68_338 ();
 sg13g2_fill_2 FILLER_68_345 ();
 sg13g2_fill_1 FILLER_68_347 ();
 sg13g2_fill_1 FILLER_68_360 ();
 sg13g2_decap_8 FILLER_68_376 ();
 sg13g2_decap_4 FILLER_68_383 ();
 sg13g2_fill_1 FILLER_68_387 ();
 sg13g2_fill_2 FILLER_68_392 ();
 sg13g2_decap_4 FILLER_68_399 ();
 sg13g2_fill_1 FILLER_68_403 ();
 sg13g2_decap_4 FILLER_68_424 ();
 sg13g2_fill_1 FILLER_68_428 ();
 sg13g2_decap_8 FILLER_68_469 ();
 sg13g2_fill_2 FILLER_68_476 ();
 sg13g2_fill_1 FILLER_68_478 ();
 sg13g2_fill_2 FILLER_68_488 ();
 sg13g2_fill_1 FILLER_68_500 ();
 sg13g2_decap_8 FILLER_68_506 ();
 sg13g2_fill_2 FILLER_68_513 ();
 sg13g2_fill_1 FILLER_68_515 ();
 sg13g2_decap_8 FILLER_68_521 ();
 sg13g2_decap_4 FILLER_68_528 ();
 sg13g2_fill_2 FILLER_68_532 ();
 sg13g2_fill_2 FILLER_68_543 ();
 sg13g2_fill_2 FILLER_68_551 ();
 sg13g2_fill_1 FILLER_68_553 ();
 sg13g2_fill_2 FILLER_68_565 ();
 sg13g2_fill_1 FILLER_68_567 ();
 sg13g2_fill_1 FILLER_68_572 ();
 sg13g2_decap_8 FILLER_68_579 ();
 sg13g2_fill_2 FILLER_68_586 ();
 sg13g2_fill_1 FILLER_68_588 ();
 sg13g2_decap_8 FILLER_68_594 ();
 sg13g2_fill_2 FILLER_68_601 ();
 sg13g2_decap_8 FILLER_68_608 ();
 sg13g2_fill_2 FILLER_68_615 ();
 sg13g2_decap_8 FILLER_68_623 ();
 sg13g2_decap_8 FILLER_68_630 ();
 sg13g2_decap_4 FILLER_68_637 ();
 sg13g2_decap_8 FILLER_68_660 ();
 sg13g2_fill_2 FILLER_68_667 ();
 sg13g2_fill_1 FILLER_68_677 ();
 sg13g2_fill_2 FILLER_68_694 ();
 sg13g2_fill_1 FILLER_68_696 ();
 sg13g2_decap_4 FILLER_68_703 ();
 sg13g2_decap_4 FILLER_68_718 ();
 sg13g2_decap_4 FILLER_68_734 ();
 sg13g2_fill_1 FILLER_68_738 ();
 sg13g2_decap_8 FILLER_68_744 ();
 sg13g2_decap_8 FILLER_68_751 ();
 sg13g2_fill_2 FILLER_68_758 ();
 sg13g2_fill_1 FILLER_68_760 ();
 sg13g2_fill_2 FILLER_68_765 ();
 sg13g2_decap_4 FILLER_68_788 ();
 sg13g2_fill_2 FILLER_68_792 ();
 sg13g2_fill_2 FILLER_68_818 ();
 sg13g2_fill_1 FILLER_68_820 ();
 sg13g2_fill_2 FILLER_68_827 ();
 sg13g2_fill_1 FILLER_68_847 ();
 sg13g2_decap_4 FILLER_68_856 ();
 sg13g2_fill_2 FILLER_68_860 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_fill_1 FILLER_69_30 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_fill_2 FILLER_69_47 ();
 sg13g2_fill_2 FILLER_69_54 ();
 sg13g2_fill_2 FILLER_69_60 ();
 sg13g2_decap_4 FILLER_69_74 ();
 sg13g2_fill_1 FILLER_69_78 ();
 sg13g2_fill_2 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_94 ();
 sg13g2_decap_4 FILLER_69_101 ();
 sg13g2_fill_2 FILLER_69_110 ();
 sg13g2_fill_1 FILLER_69_112 ();
 sg13g2_fill_2 FILLER_69_128 ();
 sg13g2_decap_8 FILLER_69_147 ();
 sg13g2_decap_8 FILLER_69_154 ();
 sg13g2_decap_8 FILLER_69_161 ();
 sg13g2_fill_2 FILLER_69_173 ();
 sg13g2_fill_2 FILLER_69_180 ();
 sg13g2_decap_4 FILLER_69_208 ();
 sg13g2_fill_1 FILLER_69_212 ();
 sg13g2_fill_2 FILLER_69_259 ();
 sg13g2_fill_1 FILLER_69_261 ();
 sg13g2_fill_2 FILLER_69_267 ();
 sg13g2_fill_1 FILLER_69_269 ();
 sg13g2_decap_4 FILLER_69_275 ();
 sg13g2_fill_2 FILLER_69_279 ();
 sg13g2_decap_8 FILLER_69_343 ();
 sg13g2_fill_2 FILLER_69_350 ();
 sg13g2_fill_2 FILLER_69_365 ();
 sg13g2_fill_1 FILLER_69_367 ();
 sg13g2_fill_1 FILLER_69_377 ();
 sg13g2_decap_8 FILLER_69_404 ();
 sg13g2_decap_8 FILLER_69_411 ();
 sg13g2_decap_4 FILLER_69_418 ();
 sg13g2_fill_2 FILLER_69_422 ();
 sg13g2_fill_2 FILLER_69_437 ();
 sg13g2_decap_8 FILLER_69_443 ();
 sg13g2_fill_2 FILLER_69_450 ();
 sg13g2_fill_1 FILLER_69_452 ();
 sg13g2_decap_8 FILLER_69_467 ();
 sg13g2_fill_2 FILLER_69_474 ();
 sg13g2_fill_2 FILLER_69_494 ();
 sg13g2_fill_1 FILLER_69_496 ();
 sg13g2_fill_2 FILLER_69_502 ();
 sg13g2_decap_4 FILLER_69_522 ();
 sg13g2_fill_1 FILLER_69_526 ();
 sg13g2_fill_2 FILLER_69_539 ();
 sg13g2_fill_1 FILLER_69_541 ();
 sg13g2_decap_8 FILLER_69_551 ();
 sg13g2_decap_4 FILLER_69_558 ();
 sg13g2_fill_2 FILLER_69_562 ();
 sg13g2_fill_1 FILLER_69_588 ();
 sg13g2_fill_2 FILLER_69_613 ();
 sg13g2_fill_1 FILLER_69_615 ();
 sg13g2_decap_8 FILLER_69_633 ();
 sg13g2_fill_2 FILLER_69_640 ();
 sg13g2_decap_8 FILLER_69_651 ();
 sg13g2_decap_4 FILLER_69_658 ();
 sg13g2_decap_8 FILLER_69_684 ();
 sg13g2_decap_4 FILLER_69_691 ();
 sg13g2_fill_1 FILLER_69_695 ();
 sg13g2_decap_8 FILLER_69_704 ();
 sg13g2_decap_4 FILLER_69_711 ();
 sg13g2_fill_2 FILLER_69_715 ();
 sg13g2_fill_1 FILLER_69_736 ();
 sg13g2_decap_8 FILLER_69_745 ();
 sg13g2_fill_1 FILLER_69_752 ();
 sg13g2_fill_1 FILLER_69_778 ();
 sg13g2_fill_2 FILLER_69_793 ();
 sg13g2_decap_8 FILLER_69_800 ();
 sg13g2_decap_8 FILLER_69_815 ();
 sg13g2_decap_8 FILLER_69_827 ();
 sg13g2_fill_2 FILLER_69_834 ();
 sg13g2_decap_4 FILLER_69_856 ();
 sg13g2_fill_2 FILLER_69_860 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_4 FILLER_70_7 ();
 sg13g2_fill_2 FILLER_70_11 ();
 sg13g2_decap_8 FILLER_70_27 ();
 sg13g2_fill_1 FILLER_70_34 ();
 sg13g2_fill_2 FILLER_70_56 ();
 sg13g2_fill_2 FILLER_70_78 ();
 sg13g2_decap_8 FILLER_70_96 ();
 sg13g2_decap_8 FILLER_70_103 ();
 sg13g2_decap_8 FILLER_70_110 ();
 sg13g2_fill_1 FILLER_70_132 ();
 sg13g2_decap_4 FILLER_70_149 ();
 sg13g2_fill_2 FILLER_70_153 ();
 sg13g2_decap_8 FILLER_70_160 ();
 sg13g2_decap_4 FILLER_70_167 ();
 sg13g2_fill_2 FILLER_70_171 ();
 sg13g2_fill_2 FILLER_70_176 ();
 sg13g2_decap_8 FILLER_70_216 ();
 sg13g2_fill_2 FILLER_70_223 ();
 sg13g2_fill_1 FILLER_70_225 ();
 sg13g2_fill_2 FILLER_70_252 ();
 sg13g2_fill_1 FILLER_70_254 ();
 sg13g2_fill_1 FILLER_70_271 ();
 sg13g2_decap_4 FILLER_70_276 ();
 sg13g2_fill_1 FILLER_70_280 ();
 sg13g2_fill_2 FILLER_70_326 ();
 sg13g2_fill_1 FILLER_70_328 ();
 sg13g2_decap_8 FILLER_70_342 ();
 sg13g2_fill_2 FILLER_70_349 ();
 sg13g2_fill_2 FILLER_70_355 ();
 sg13g2_fill_1 FILLER_70_383 ();
 sg13g2_decap_4 FILLER_70_392 ();
 sg13g2_decap_4 FILLER_70_401 ();
 sg13g2_decap_4 FILLER_70_426 ();
 sg13g2_fill_1 FILLER_70_430 ();
 sg13g2_fill_2 FILLER_70_452 ();
 sg13g2_decap_4 FILLER_70_476 ();
 sg13g2_fill_1 FILLER_70_480 ();
 sg13g2_decap_4 FILLER_70_487 ();
 sg13g2_fill_2 FILLER_70_515 ();
 sg13g2_fill_1 FILLER_70_517 ();
 sg13g2_fill_2 FILLER_70_529 ();
 sg13g2_fill_1 FILLER_70_531 ();
 sg13g2_decap_4 FILLER_70_559 ();
 sg13g2_decap_8 FILLER_70_577 ();
 sg13g2_fill_1 FILLER_70_584 ();
 sg13g2_decap_8 FILLER_70_595 ();
 sg13g2_fill_1 FILLER_70_602 ();
 sg13g2_decap_4 FILLER_70_608 ();
 sg13g2_fill_1 FILLER_70_612 ();
 sg13g2_decap_8 FILLER_70_623 ();
 sg13g2_fill_2 FILLER_70_630 ();
 sg13g2_fill_1 FILLER_70_632 ();
 sg13g2_fill_1 FILLER_70_660 ();
 sg13g2_fill_1 FILLER_70_671 ();
 sg13g2_decap_8 FILLER_70_684 ();
 sg13g2_fill_1 FILLER_70_691 ();
 sg13g2_fill_2 FILLER_70_705 ();
 sg13g2_decap_8 FILLER_70_730 ();
 sg13g2_decap_4 FILLER_70_742 ();
 sg13g2_decap_8 FILLER_70_750 ();
 sg13g2_fill_1 FILLER_70_757 ();
 sg13g2_decap_8 FILLER_70_764 ();
 sg13g2_fill_1 FILLER_70_776 ();
 sg13g2_decap_4 FILLER_70_797 ();
 sg13g2_fill_2 FILLER_70_807 ();
 sg13g2_fill_2 FILLER_70_820 ();
 sg13g2_fill_1 FILLER_70_822 ();
 sg13g2_decap_8 FILLER_70_837 ();
 sg13g2_fill_1 FILLER_70_844 ();
 sg13g2_decap_8 FILLER_70_849 ();
 sg13g2_decap_4 FILLER_70_856 ();
 sg13g2_fill_2 FILLER_70_860 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_4 FILLER_71_37 ();
 sg13g2_decap_8 FILLER_71_48 ();
 sg13g2_decap_4 FILLER_71_55 ();
 sg13g2_decap_8 FILLER_71_76 ();
 sg13g2_fill_1 FILLER_71_83 ();
 sg13g2_decap_8 FILLER_71_101 ();
 sg13g2_fill_2 FILLER_71_108 ();
 sg13g2_fill_2 FILLER_71_119 ();
 sg13g2_fill_1 FILLER_71_136 ();
 sg13g2_decap_8 FILLER_71_143 ();
 sg13g2_fill_2 FILLER_71_150 ();
 sg13g2_decap_8 FILLER_71_191 ();
 sg13g2_fill_2 FILLER_71_198 ();
 sg13g2_fill_1 FILLER_71_200 ();
 sg13g2_decap_8 FILLER_71_205 ();
 sg13g2_decap_8 FILLER_71_212 ();
 sg13g2_decap_4 FILLER_71_219 ();
 sg13g2_fill_1 FILLER_71_249 ();
 sg13g2_fill_2 FILLER_71_260 ();
 sg13g2_decap_8 FILLER_71_272 ();
 sg13g2_fill_2 FILLER_71_374 ();
 sg13g2_decap_8 FILLER_71_407 ();
 sg13g2_decap_8 FILLER_71_414 ();
 sg13g2_decap_8 FILLER_71_421 ();
 sg13g2_decap_4 FILLER_71_428 ();
 sg13g2_decap_8 FILLER_71_445 ();
 sg13g2_decap_8 FILLER_71_452 ();
 sg13g2_fill_2 FILLER_71_471 ();
 sg13g2_decap_4 FILLER_71_478 ();
 sg13g2_decap_8 FILLER_71_487 ();
 sg13g2_decap_4 FILLER_71_494 ();
 sg13g2_fill_1 FILLER_71_498 ();
 sg13g2_decap_8 FILLER_71_504 ();
 sg13g2_fill_2 FILLER_71_511 ();
 sg13g2_fill_2 FILLER_71_534 ();
 sg13g2_fill_1 FILLER_71_536 ();
 sg13g2_decap_8 FILLER_71_543 ();
 sg13g2_decap_8 FILLER_71_550 ();
 sg13g2_decap_4 FILLER_71_557 ();
 sg13g2_fill_1 FILLER_71_561 ();
 sg13g2_decap_4 FILLER_71_580 ();
 sg13g2_fill_1 FILLER_71_584 ();
 sg13g2_fill_1 FILLER_71_603 ();
 sg13g2_decap_4 FILLER_71_633 ();
 sg13g2_fill_2 FILLER_71_637 ();
 sg13g2_decap_8 FILLER_71_643 ();
 sg13g2_decap_4 FILLER_71_650 ();
 sg13g2_fill_1 FILLER_71_654 ();
 sg13g2_fill_2 FILLER_71_659 ();
 sg13g2_decap_8 FILLER_71_678 ();
 sg13g2_decap_4 FILLER_71_685 ();
 sg13g2_fill_2 FILLER_71_689 ();
 sg13g2_decap_8 FILLER_71_708 ();
 sg13g2_fill_2 FILLER_71_715 ();
 sg13g2_fill_1 FILLER_71_717 ();
 sg13g2_decap_4 FILLER_71_727 ();
 sg13g2_fill_1 FILLER_71_731 ();
 sg13g2_fill_1 FILLER_71_738 ();
 sg13g2_decap_4 FILLER_71_770 ();
 sg13g2_fill_1 FILLER_71_774 ();
 sg13g2_fill_2 FILLER_71_790 ();
 sg13g2_decap_8 FILLER_71_797 ();
 sg13g2_decap_4 FILLER_71_804 ();
 sg13g2_fill_1 FILLER_71_808 ();
 sg13g2_fill_2 FILLER_71_819 ();
 sg13g2_decap_4 FILLER_71_826 ();
 sg13g2_fill_2 FILLER_71_838 ();
 sg13g2_fill_1 FILLER_71_840 ();
 sg13g2_fill_1 FILLER_71_847 ();
 sg13g2_decap_8 FILLER_71_853 ();
 sg13g2_fill_2 FILLER_71_860 ();
 sg13g2_decap_4 FILLER_72_0 ();
 sg13g2_fill_1 FILLER_72_4 ();
 sg13g2_decap_8 FILLER_72_29 ();
 sg13g2_decap_8 FILLER_72_36 ();
 sg13g2_decap_4 FILLER_72_43 ();
 sg13g2_fill_2 FILLER_72_47 ();
 sg13g2_fill_2 FILLER_72_54 ();
 sg13g2_fill_1 FILLER_72_56 ();
 sg13g2_fill_1 FILLER_72_62 ();
 sg13g2_decap_4 FILLER_72_73 ();
 sg13g2_decap_4 FILLER_72_84 ();
 sg13g2_fill_1 FILLER_72_88 ();
 sg13g2_decap_4 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_143 ();
 sg13g2_decap_8 FILLER_72_150 ();
 sg13g2_fill_1 FILLER_72_162 ();
 sg13g2_fill_1 FILLER_72_170 ();
 sg13g2_decap_4 FILLER_72_206 ();
 sg13g2_fill_2 FILLER_72_236 ();
 sg13g2_fill_2 FILLER_72_262 ();
 sg13g2_fill_2 FILLER_72_274 ();
 sg13g2_fill_1 FILLER_72_276 ();
 sg13g2_fill_2 FILLER_72_287 ();
 sg13g2_fill_2 FILLER_72_294 ();
 sg13g2_fill_1 FILLER_72_296 ();
 sg13g2_fill_2 FILLER_72_304 ();
 sg13g2_fill_1 FILLER_72_306 ();
 sg13g2_fill_2 FILLER_72_316 ();
 sg13g2_fill_2 FILLER_72_348 ();
 sg13g2_decap_8 FILLER_72_354 ();
 sg13g2_decap_8 FILLER_72_361 ();
 sg13g2_fill_2 FILLER_72_408 ();
 sg13g2_fill_1 FILLER_72_410 ();
 sg13g2_decap_4 FILLER_72_425 ();
 sg13g2_fill_1 FILLER_72_429 ();
 sg13g2_decap_4 FILLER_72_451 ();
 sg13g2_fill_1 FILLER_72_455 ();
 sg13g2_fill_2 FILLER_72_472 ();
 sg13g2_fill_1 FILLER_72_486 ();
 sg13g2_decap_4 FILLER_72_512 ();
 sg13g2_fill_2 FILLER_72_521 ();
 sg13g2_fill_1 FILLER_72_523 ();
 sg13g2_fill_2 FILLER_72_529 ();
 sg13g2_fill_1 FILLER_72_531 ();
 sg13g2_decap_4 FILLER_72_551 ();
 sg13g2_fill_2 FILLER_72_560 ();
 sg13g2_fill_1 FILLER_72_562 ();
 sg13g2_decap_8 FILLER_72_579 ();
 sg13g2_decap_8 FILLER_72_586 ();
 sg13g2_decap_8 FILLER_72_603 ();
 sg13g2_fill_1 FILLER_72_610 ();
 sg13g2_fill_1 FILLER_72_616 ();
 sg13g2_fill_1 FILLER_72_635 ();
 sg13g2_decap_8 FILLER_72_641 ();
 sg13g2_decap_8 FILLER_72_648 ();
 sg13g2_fill_2 FILLER_72_655 ();
 sg13g2_decap_4 FILLER_72_681 ();
 sg13g2_fill_1 FILLER_72_685 ();
 sg13g2_fill_2 FILLER_72_710 ();
 sg13g2_fill_1 FILLER_72_712 ();
 sg13g2_decap_8 FILLER_72_751 ();
 sg13g2_decap_8 FILLER_72_758 ();
 sg13g2_decap_4 FILLER_72_765 ();
 sg13g2_fill_2 FILLER_72_769 ();
 sg13g2_decap_4 FILLER_72_776 ();
 sg13g2_fill_1 FILLER_72_780 ();
 sg13g2_decap_8 FILLER_72_801 ();
 sg13g2_fill_2 FILLER_72_808 ();
 sg13g2_fill_1 FILLER_72_817 ();
 sg13g2_decap_4 FILLER_72_833 ();
 sg13g2_fill_2 FILLER_72_845 ();
 sg13g2_fill_2 FILLER_72_860 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_fill_2 FILLER_73_7 ();
 sg13g2_fill_1 FILLER_73_9 ();
 sg13g2_decap_4 FILLER_73_33 ();
 sg13g2_fill_2 FILLER_73_37 ();
 sg13g2_fill_1 FILLER_73_45 ();
 sg13g2_decap_4 FILLER_73_68 ();
 sg13g2_fill_1 FILLER_73_72 ();
 sg13g2_fill_2 FILLER_73_79 ();
 sg13g2_fill_1 FILLER_73_81 ();
 sg13g2_decap_8 FILLER_73_95 ();
 sg13g2_decap_4 FILLER_73_102 ();
 sg13g2_fill_2 FILLER_73_106 ();
 sg13g2_decap_8 FILLER_73_119 ();
 sg13g2_fill_2 FILLER_73_126 ();
 sg13g2_decap_8 FILLER_73_138 ();
 sg13g2_decap_4 FILLER_73_145 ();
 sg13g2_fill_2 FILLER_73_169 ();
 sg13g2_fill_1 FILLER_73_171 ();
 sg13g2_fill_2 FILLER_73_189 ();
 sg13g2_decap_4 FILLER_73_199 ();
 sg13g2_fill_2 FILLER_73_203 ();
 sg13g2_fill_2 FILLER_73_213 ();
 sg13g2_fill_2 FILLER_73_233 ();
 sg13g2_fill_1 FILLER_73_250 ();
 sg13g2_fill_2 FILLER_73_276 ();
 sg13g2_fill_1 FILLER_73_278 ();
 sg13g2_fill_2 FILLER_73_305 ();
 sg13g2_fill_1 FILLER_73_307 ();
 sg13g2_fill_2 FILLER_73_318 ();
 sg13g2_fill_1 FILLER_73_320 ();
 sg13g2_fill_2 FILLER_73_331 ();
 sg13g2_fill_1 FILLER_73_333 ();
 sg13g2_decap_4 FILLER_73_359 ();
 sg13g2_fill_1 FILLER_73_363 ();
 sg13g2_fill_2 FILLER_73_372 ();
 sg13g2_fill_2 FILLER_73_390 ();
 sg13g2_fill_1 FILLER_73_400 ();
 sg13g2_decap_8 FILLER_73_419 ();
 sg13g2_decap_8 FILLER_73_426 ();
 sg13g2_decap_8 FILLER_73_438 ();
 sg13g2_fill_1 FILLER_73_445 ();
 sg13g2_fill_1 FILLER_73_454 ();
 sg13g2_decap_8 FILLER_73_478 ();
 sg13g2_fill_2 FILLER_73_485 ();
 sg13g2_fill_1 FILLER_73_487 ();
 sg13g2_decap_4 FILLER_73_499 ();
 sg13g2_fill_2 FILLER_73_503 ();
 sg13g2_decap_4 FILLER_73_513 ();
 sg13g2_fill_2 FILLER_73_517 ();
 sg13g2_fill_1 FILLER_73_523 ();
 sg13g2_decap_8 FILLER_73_530 ();
 sg13g2_decap_4 FILLER_73_537 ();
 sg13g2_fill_2 FILLER_73_541 ();
 sg13g2_fill_2 FILLER_73_560 ();
 sg13g2_fill_2 FILLER_73_566 ();
 sg13g2_fill_1 FILLER_73_568 ();
 sg13g2_fill_1 FILLER_73_585 ();
 sg13g2_fill_1 FILLER_73_608 ();
 sg13g2_fill_2 FILLER_73_614 ();
 sg13g2_fill_1 FILLER_73_616 ();
 sg13g2_decap_8 FILLER_73_630 ();
 sg13g2_fill_2 FILLER_73_637 ();
 sg13g2_decap_4 FILLER_73_656 ();
 sg13g2_fill_2 FILLER_73_660 ();
 sg13g2_fill_1 FILLER_73_667 ();
 sg13g2_decap_8 FILLER_73_673 ();
 sg13g2_decap_8 FILLER_73_680 ();
 sg13g2_decap_4 FILLER_73_707 ();
 sg13g2_decap_8 FILLER_73_725 ();
 sg13g2_fill_1 FILLER_73_732 ();
 sg13g2_fill_1 FILLER_73_738 ();
 sg13g2_fill_2 FILLER_73_755 ();
 sg13g2_fill_1 FILLER_73_757 ();
 sg13g2_fill_2 FILLER_73_772 ();
 sg13g2_fill_2 FILLER_73_788 ();
 sg13g2_fill_1 FILLER_73_790 ();
 sg13g2_fill_2 FILLER_73_801 ();
 sg13g2_fill_1 FILLER_73_803 ();
 sg13g2_decap_4 FILLER_73_808 ();
 sg13g2_decap_8 FILLER_73_829 ();
 sg13g2_decap_4 FILLER_73_836 ();
 sg13g2_decap_4 FILLER_73_856 ();
 sg13g2_fill_2 FILLER_73_860 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_fill_2 FILLER_74_7 ();
 sg13g2_fill_2 FILLER_74_33 ();
 sg13g2_fill_2 FILLER_74_54 ();
 sg13g2_fill_1 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_62 ();
 sg13g2_decap_4 FILLER_74_69 ();
 sg13g2_fill_1 FILLER_74_73 ();
 sg13g2_decap_4 FILLER_74_94 ();
 sg13g2_fill_2 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_128 ();
 sg13g2_decap_8 FILLER_74_139 ();
 sg13g2_fill_2 FILLER_74_146 ();
 sg13g2_decap_4 FILLER_74_152 ();
 sg13g2_decap_4 FILLER_74_160 ();
 sg13g2_fill_2 FILLER_74_164 ();
 sg13g2_decap_4 FILLER_74_171 ();
 sg13g2_fill_1 FILLER_74_175 ();
 sg13g2_fill_2 FILLER_74_278 ();
 sg13g2_fill_2 FILLER_74_289 ();
 sg13g2_fill_1 FILLER_74_291 ();
 sg13g2_fill_1 FILLER_74_318 ();
 sg13g2_fill_2 FILLER_74_338 ();
 sg13g2_decap_4 FILLER_74_366 ();
 sg13g2_fill_2 FILLER_74_370 ();
 sg13g2_fill_2 FILLER_74_387 ();
 sg13g2_fill_1 FILLER_74_389 ();
 sg13g2_fill_1 FILLER_74_396 ();
 sg13g2_decap_8 FILLER_74_413 ();
 sg13g2_decap_4 FILLER_74_420 ();
 sg13g2_fill_2 FILLER_74_445 ();
 sg13g2_fill_1 FILLER_74_447 ();
 sg13g2_decap_8 FILLER_74_454 ();
 sg13g2_decap_4 FILLER_74_461 ();
 sg13g2_fill_2 FILLER_74_476 ();
 sg13g2_fill_1 FILLER_74_478 ();
 sg13g2_fill_2 FILLER_74_508 ();
 sg13g2_fill_1 FILLER_74_528 ();
 sg13g2_decap_4 FILLER_74_542 ();
 sg13g2_decap_8 FILLER_74_560 ();
 sg13g2_fill_1 FILLER_74_567 ();
 sg13g2_decap_8 FILLER_74_583 ();
 sg13g2_fill_2 FILLER_74_590 ();
 sg13g2_fill_1 FILLER_74_592 ();
 sg13g2_decap_8 FILLER_74_608 ();
 sg13g2_fill_2 FILLER_74_620 ();
 sg13g2_decap_4 FILLER_74_642 ();
 sg13g2_fill_1 FILLER_74_646 ();
 sg13g2_fill_2 FILLER_74_652 ();
 sg13g2_fill_1 FILLER_74_654 ();
 sg13g2_decap_8 FILLER_74_680 ();
 sg13g2_decap_4 FILLER_74_687 ();
 sg13g2_fill_2 FILLER_74_696 ();
 sg13g2_fill_1 FILLER_74_698 ();
 sg13g2_fill_1 FILLER_74_712 ();
 sg13g2_decap_8 FILLER_74_737 ();
 sg13g2_fill_2 FILLER_74_744 ();
 sg13g2_fill_1 FILLER_74_746 ();
 sg13g2_decap_4 FILLER_74_753 ();
 sg13g2_fill_1 FILLER_74_757 ();
 sg13g2_decap_8 FILLER_74_780 ();
 sg13g2_decap_8 FILLER_74_787 ();
 sg13g2_fill_2 FILLER_74_794 ();
 sg13g2_fill_2 FILLER_74_811 ();
 sg13g2_fill_1 FILLER_74_832 ();
 sg13g2_fill_2 FILLER_74_859 ();
 sg13g2_fill_1 FILLER_74_861 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_fill_1 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_33 ();
 sg13g2_decap_8 FILLER_75_40 ();
 sg13g2_fill_2 FILLER_75_47 ();
 sg13g2_fill_2 FILLER_75_58 ();
 sg13g2_fill_2 FILLER_75_80 ();
 sg13g2_decap_8 FILLER_75_113 ();
 sg13g2_decap_4 FILLER_75_120 ();
 sg13g2_decap_4 FILLER_75_155 ();
 sg13g2_fill_2 FILLER_75_190 ();
 sg13g2_fill_1 FILLER_75_245 ();
 sg13g2_fill_2 FILLER_75_260 ();
 sg13g2_fill_2 FILLER_75_276 ();
 sg13g2_fill_2 FILLER_75_299 ();
 sg13g2_fill_1 FILLER_75_301 ();
 sg13g2_fill_2 FILLER_75_306 ();
 sg13g2_fill_1 FILLER_75_308 ();
 sg13g2_fill_2 FILLER_75_323 ();
 sg13g2_fill_2 FILLER_75_343 ();
 sg13g2_decap_8 FILLER_75_406 ();
 sg13g2_decap_8 FILLER_75_413 ();
 sg13g2_decap_8 FILLER_75_420 ();
 sg13g2_decap_4 FILLER_75_427 ();
 sg13g2_decap_8 FILLER_75_436 ();
 sg13g2_fill_1 FILLER_75_443 ();
 sg13g2_fill_2 FILLER_75_460 ();
 sg13g2_fill_1 FILLER_75_462 ();
 sg13g2_decap_4 FILLER_75_472 ();
 sg13g2_fill_2 FILLER_75_476 ();
 sg13g2_fill_2 FILLER_75_483 ();
 sg13g2_fill_1 FILLER_75_485 ();
 sg13g2_decap_4 FILLER_75_494 ();
 sg13g2_fill_1 FILLER_75_498 ();
 sg13g2_fill_1 FILLER_75_505 ();
 sg13g2_decap_8 FILLER_75_510 ();
 sg13g2_fill_2 FILLER_75_517 ();
 sg13g2_fill_1 FILLER_75_519 ();
 sg13g2_decap_8 FILLER_75_524 ();
 sg13g2_fill_1 FILLER_75_531 ();
 sg13g2_decap_8 FILLER_75_542 ();
 sg13g2_fill_2 FILLER_75_549 ();
 sg13g2_fill_1 FILLER_75_551 ();
 sg13g2_decap_8 FILLER_75_557 ();
 sg13g2_decap_8 FILLER_75_569 ();
 sg13g2_fill_1 FILLER_75_576 ();
 sg13g2_fill_2 FILLER_75_598 ();
 sg13g2_decap_8 FILLER_75_605 ();
 sg13g2_fill_2 FILLER_75_612 ();
 sg13g2_fill_1 FILLER_75_619 ();
 sg13g2_fill_1 FILLER_75_625 ();
 sg13g2_decap_8 FILLER_75_630 ();
 sg13g2_decap_8 FILLER_75_659 ();
 sg13g2_fill_1 FILLER_75_666 ();
 sg13g2_fill_2 FILLER_75_681 ();
 sg13g2_fill_1 FILLER_75_689 ();
 sg13g2_decap_8 FILLER_75_712 ();
 sg13g2_decap_4 FILLER_75_719 ();
 sg13g2_decap_4 FILLER_75_727 ();
 sg13g2_fill_2 FILLER_75_731 ();
 sg13g2_decap_8 FILLER_75_746 ();
 sg13g2_fill_2 FILLER_75_759 ();
 sg13g2_fill_1 FILLER_75_761 ();
 sg13g2_fill_2 FILLER_75_768 ();
 sg13g2_fill_1 FILLER_75_770 ();
 sg13g2_fill_1 FILLER_75_782 ();
 sg13g2_fill_2 FILLER_75_796 ();
 sg13g2_fill_1 FILLER_75_798 ();
 sg13g2_decap_8 FILLER_75_815 ();
 sg13g2_decap_8 FILLER_75_822 ();
 sg13g2_fill_1 FILLER_75_829 ();
 sg13g2_decap_4 FILLER_75_846 ();
 sg13g2_decap_4 FILLER_75_858 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_4 FILLER_76_7 ();
 sg13g2_fill_1 FILLER_76_11 ();
 sg13g2_fill_2 FILLER_76_39 ();
 sg13g2_fill_1 FILLER_76_45 ();
 sg13g2_fill_2 FILLER_76_55 ();
 sg13g2_fill_1 FILLER_76_57 ();
 sg13g2_decap_8 FILLER_76_66 ();
 sg13g2_fill_1 FILLER_76_73 ();
 sg13g2_fill_2 FILLER_76_87 ();
 sg13g2_decap_8 FILLER_76_118 ();
 sg13g2_decap_8 FILLER_76_125 ();
 sg13g2_decap_4 FILLER_76_132 ();
 sg13g2_fill_2 FILLER_76_136 ();
 sg13g2_fill_1 FILLER_76_147 ();
 sg13g2_fill_1 FILLER_76_189 ();
 sg13g2_decap_8 FILLER_76_195 ();
 sg13g2_decap_8 FILLER_76_202 ();
 sg13g2_fill_1 FILLER_76_227 ();
 sg13g2_fill_1 FILLER_76_237 ();
 sg13g2_fill_2 FILLER_76_252 ();
 sg13g2_fill_1 FILLER_76_254 ();
 sg13g2_fill_2 FILLER_76_280 ();
 sg13g2_fill_1 FILLER_76_282 ();
 sg13g2_fill_2 FILLER_76_309 ();
 sg13g2_fill_1 FILLER_76_361 ();
 sg13g2_fill_2 FILLER_76_391 ();
 sg13g2_decap_8 FILLER_76_399 ();
 sg13g2_fill_1 FILLER_76_406 ();
 sg13g2_decap_4 FILLER_76_414 ();
 sg13g2_fill_2 FILLER_76_418 ();
 sg13g2_decap_4 FILLER_76_442 ();
 sg13g2_fill_1 FILLER_76_446 ();
 sg13g2_fill_2 FILLER_76_464 ();
 sg13g2_decap_8 FILLER_76_484 ();
 sg13g2_fill_2 FILLER_76_491 ();
 sg13g2_fill_2 FILLER_76_501 ();
 sg13g2_fill_1 FILLER_76_503 ();
 sg13g2_fill_2 FILLER_76_524 ();
 sg13g2_fill_1 FILLER_76_526 ();
 sg13g2_fill_1 FILLER_76_540 ();
 sg13g2_fill_2 FILLER_76_577 ();
 sg13g2_fill_1 FILLER_76_579 ();
 sg13g2_decap_4 FILLER_76_585 ();
 sg13g2_fill_2 FILLER_76_589 ();
 sg13g2_fill_2 FILLER_76_609 ();
 sg13g2_fill_1 FILLER_76_611 ();
 sg13g2_decap_8 FILLER_76_630 ();
 sg13g2_fill_2 FILLER_76_637 ();
 sg13g2_fill_1 FILLER_76_639 ();
 sg13g2_decap_8 FILLER_76_650 ();
 sg13g2_decap_4 FILLER_76_657 ();
 sg13g2_fill_1 FILLER_76_689 ();
 sg13g2_fill_2 FILLER_76_696 ();
 sg13g2_decap_4 FILLER_76_709 ();
 sg13g2_fill_1 FILLER_76_713 ();
 sg13g2_decap_4 FILLER_76_740 ();
 sg13g2_fill_2 FILLER_76_744 ();
 sg13g2_fill_2 FILLER_76_773 ();
 sg13g2_fill_1 FILLER_76_775 ();
 sg13g2_fill_2 FILLER_76_781 ();
 sg13g2_fill_1 FILLER_76_783 ();
 sg13g2_fill_2 FILLER_76_809 ();
 sg13g2_fill_1 FILLER_76_811 ();
 sg13g2_fill_2 FILLER_76_820 ();
 sg13g2_fill_1 FILLER_76_822 ();
 sg13g2_decap_8 FILLER_76_831 ();
 sg13g2_fill_2 FILLER_76_838 ();
 sg13g2_decap_8 FILLER_76_853 ();
 sg13g2_fill_2 FILLER_76_860 ();
 sg13g2_fill_2 FILLER_77_0 ();
 sg13g2_fill_2 FILLER_77_30 ();
 sg13g2_fill_2 FILLER_77_37 ();
 sg13g2_fill_1 FILLER_77_39 ();
 sg13g2_fill_2 FILLER_77_48 ();
 sg13g2_fill_1 FILLER_77_50 ();
 sg13g2_fill_1 FILLER_77_67 ();
 sg13g2_fill_2 FILLER_77_80 ();
 sg13g2_decap_8 FILLER_77_94 ();
 sg13g2_decap_8 FILLER_77_101 ();
 sg13g2_fill_2 FILLER_77_108 ();
 sg13g2_fill_2 FILLER_77_119 ();
 sg13g2_decap_4 FILLER_77_156 ();
 sg13g2_decap_8 FILLER_77_168 ();
 sg13g2_fill_2 FILLER_77_183 ();
 sg13g2_fill_1 FILLER_77_185 ();
 sg13g2_fill_2 FILLER_77_200 ();
 sg13g2_fill_1 FILLER_77_254 ();
 sg13g2_fill_2 FILLER_77_290 ();
 sg13g2_fill_1 FILLER_77_336 ();
 sg13g2_fill_1 FILLER_77_372 ();
 sg13g2_fill_2 FILLER_77_377 ();
 sg13g2_decap_4 FILLER_77_447 ();
 sg13g2_fill_2 FILLER_77_451 ();
 sg13g2_decap_8 FILLER_77_461 ();
 sg13g2_decap_8 FILLER_77_468 ();
 sg13g2_decap_8 FILLER_77_491 ();
 sg13g2_decap_8 FILLER_77_498 ();
 sg13g2_fill_1 FILLER_77_505 ();
 sg13g2_fill_1 FILLER_77_512 ();
 sg13g2_fill_1 FILLER_77_519 ();
 sg13g2_fill_2 FILLER_77_526 ();
 sg13g2_fill_2 FILLER_77_533 ();
 sg13g2_decap_8 FILLER_77_540 ();
 sg13g2_decap_8 FILLER_77_547 ();
 sg13g2_fill_2 FILLER_77_554 ();
 sg13g2_decap_8 FILLER_77_567 ();
 sg13g2_fill_1 FILLER_77_574 ();
 sg13g2_fill_1 FILLER_77_587 ();
 sg13g2_fill_2 FILLER_77_601 ();
 sg13g2_fill_2 FILLER_77_611 ();
 sg13g2_decap_8 FILLER_77_618 ();
 sg13g2_fill_2 FILLER_77_625 ();
 sg13g2_fill_2 FILLER_77_645 ();
 sg13g2_fill_2 FILLER_77_665 ();
 sg13g2_fill_1 FILLER_77_667 ();
 sg13g2_fill_2 FILLER_77_673 ();
 sg13g2_decap_8 FILLER_77_681 ();
 sg13g2_decap_4 FILLER_77_688 ();
 sg13g2_fill_1 FILLER_77_692 ();
 sg13g2_decap_8 FILLER_77_705 ();
 sg13g2_decap_8 FILLER_77_712 ();
 sg13g2_decap_4 FILLER_77_719 ();
 sg13g2_fill_1 FILLER_77_723 ();
 sg13g2_fill_1 FILLER_77_738 ();
 sg13g2_fill_2 FILLER_77_751 ();
 sg13g2_fill_1 FILLER_77_753 ();
 sg13g2_decap_8 FILLER_77_760 ();
 sg13g2_decap_4 FILLER_77_767 ();
 sg13g2_fill_2 FILLER_77_771 ();
 sg13g2_fill_2 FILLER_77_786 ();
 sg13g2_decap_8 FILLER_77_793 ();
 sg13g2_fill_2 FILLER_77_800 ();
 sg13g2_fill_1 FILLER_77_802 ();
 sg13g2_decap_4 FILLER_77_811 ();
 sg13g2_fill_2 FILLER_77_815 ();
 sg13g2_fill_1 FILLER_77_825 ();
 sg13g2_decap_8 FILLER_77_847 ();
 sg13g2_decap_8 FILLER_77_854 ();
 sg13g2_fill_1 FILLER_77_861 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_4 FILLER_78_7 ();
 sg13g2_fill_1 FILLER_78_11 ();
 sg13g2_decap_8 FILLER_78_30 ();
 sg13g2_decap_4 FILLER_78_37 ();
 sg13g2_fill_2 FILLER_78_41 ();
 sg13g2_decap_4 FILLER_78_65 ();
 sg13g2_decap_8 FILLER_78_74 ();
 sg13g2_decap_8 FILLER_78_81 ();
 sg13g2_decap_8 FILLER_78_88 ();
 sg13g2_fill_1 FILLER_78_95 ();
 sg13g2_fill_1 FILLER_78_144 ();
 sg13g2_fill_1 FILLER_78_153 ();
 sg13g2_decap_8 FILLER_78_167 ();
 sg13g2_fill_1 FILLER_78_174 ();
 sg13g2_fill_1 FILLER_78_293 ();
 sg13g2_fill_1 FILLER_78_354 ();
 sg13g2_fill_2 FILLER_78_373 ();
 sg13g2_fill_2 FILLER_78_387 ();
 sg13g2_fill_1 FILLER_78_398 ();
 sg13g2_decap_8 FILLER_78_425 ();
 sg13g2_fill_1 FILLER_78_432 ();
 sg13g2_decap_8 FILLER_78_446 ();
 sg13g2_fill_1 FILLER_78_453 ();
 sg13g2_decap_8 FILLER_78_480 ();
 sg13g2_fill_2 FILLER_78_487 ();
 sg13g2_decap_8 FILLER_78_505 ();
 sg13g2_fill_2 FILLER_78_512 ();
 sg13g2_decap_8 FILLER_78_519 ();
 sg13g2_decap_4 FILLER_78_526 ();
 sg13g2_decap_4 FILLER_78_546 ();
 sg13g2_fill_2 FILLER_78_550 ();
 sg13g2_fill_2 FILLER_78_568 ();
 sg13g2_fill_1 FILLER_78_570 ();
 sg13g2_fill_1 FILLER_78_587 ();
 sg13g2_decap_4 FILLER_78_596 ();
 sg13g2_fill_2 FILLER_78_612 ();
 sg13g2_fill_1 FILLER_78_642 ();
 sg13g2_fill_2 FILLER_78_651 ();
 sg13g2_fill_1 FILLER_78_653 ();
 sg13g2_decap_8 FILLER_78_660 ();
 sg13g2_fill_2 FILLER_78_667 ();
 sg13g2_fill_1 FILLER_78_669 ();
 sg13g2_fill_2 FILLER_78_686 ();
 sg13g2_decap_8 FILLER_78_708 ();
 sg13g2_fill_1 FILLER_78_715 ();
 sg13g2_fill_2 FILLER_78_724 ();
 sg13g2_fill_1 FILLER_78_726 ();
 sg13g2_decap_4 FILLER_78_735 ();
 sg13g2_fill_1 FILLER_78_739 ();
 sg13g2_fill_1 FILLER_78_764 ();
 sg13g2_decap_8 FILLER_78_770 ();
 sg13g2_fill_2 FILLER_78_777 ();
 sg13g2_decap_4 FILLER_78_783 ();
 sg13g2_decap_8 FILLER_78_801 ();
 sg13g2_fill_1 FILLER_78_808 ();
 sg13g2_fill_1 FILLER_78_829 ();
 sg13g2_decap_8 FILLER_78_835 ();
 sg13g2_decap_8 FILLER_78_842 ();
 sg13g2_decap_8 FILLER_78_849 ();
 sg13g2_decap_4 FILLER_78_856 ();
 sg13g2_fill_2 FILLER_78_860 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_fill_1 FILLER_79_14 ();
 sg13g2_fill_1 FILLER_79_30 ();
 sg13g2_fill_2 FILLER_79_46 ();
 sg13g2_fill_2 FILLER_79_65 ();
 sg13g2_fill_1 FILLER_79_67 ();
 sg13g2_decap_8 FILLER_79_76 ();
 sg13g2_decap_4 FILLER_79_83 ();
 sg13g2_fill_1 FILLER_79_87 ();
 sg13g2_fill_2 FILLER_79_150 ();
 sg13g2_fill_1 FILLER_79_152 ();
 sg13g2_decap_4 FILLER_79_204 ();
 sg13g2_fill_1 FILLER_79_208 ();
 sg13g2_fill_1 FILLER_79_240 ();
 sg13g2_decap_4 FILLER_79_245 ();
 sg13g2_fill_2 FILLER_79_249 ();
 sg13g2_decap_4 FILLER_79_277 ();
 sg13g2_fill_2 FILLER_79_281 ();
 sg13g2_fill_2 FILLER_79_461 ();
 sg13g2_fill_2 FILLER_79_508 ();
 sg13g2_fill_1 FILLER_79_510 ();
 sg13g2_decap_8 FILLER_79_524 ();
 sg13g2_decap_8 FILLER_79_531 ();
 sg13g2_decap_8 FILLER_79_538 ();
 sg13g2_decap_4 FILLER_79_545 ();
 sg13g2_fill_1 FILLER_79_549 ();
 sg13g2_decap_4 FILLER_79_554 ();
 sg13g2_fill_1 FILLER_79_558 ();
 sg13g2_decap_8 FILLER_79_564 ();
 sg13g2_decap_8 FILLER_79_571 ();
 sg13g2_fill_2 FILLER_79_578 ();
 sg13g2_fill_1 FILLER_79_580 ();
 sg13g2_decap_8 FILLER_79_585 ();
 sg13g2_fill_2 FILLER_79_592 ();
 sg13g2_fill_1 FILLER_79_594 ();
 sg13g2_decap_4 FILLER_79_603 ();
 sg13g2_fill_2 FILLER_79_607 ();
 sg13g2_decap_8 FILLER_79_615 ();
 sg13g2_decap_8 FILLER_79_622 ();
 sg13g2_decap_8 FILLER_79_629 ();
 sg13g2_decap_8 FILLER_79_658 ();
 sg13g2_fill_2 FILLER_79_665 ();
 sg13g2_fill_1 FILLER_79_667 ();
 sg13g2_decap_4 FILLER_79_672 ();
 sg13g2_decap_8 FILLER_79_681 ();
 sg13g2_fill_1 FILLER_79_700 ();
 sg13g2_fill_2 FILLER_79_720 ();
 sg13g2_fill_2 FILLER_79_738 ();
 sg13g2_fill_1 FILLER_79_740 ();
 sg13g2_fill_1 FILLER_79_749 ();
 sg13g2_decap_4 FILLER_79_758 ();
 sg13g2_fill_1 FILLER_79_782 ();
 sg13g2_decap_8 FILLER_79_803 ();
 sg13g2_decap_8 FILLER_79_810 ();
 sg13g2_fill_2 FILLER_79_817 ();
 sg13g2_fill_1 FILLER_79_819 ();
 sg13g2_decap_8 FILLER_79_825 ();
 sg13g2_decap_8 FILLER_79_832 ();
 sg13g2_decap_8 FILLER_79_839 ();
 sg13g2_decap_8 FILLER_79_846 ();
 sg13g2_decap_8 FILLER_79_853 ();
 sg13g2_fill_2 FILLER_79_860 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_4 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_29 ();
 sg13g2_decap_8 FILLER_80_36 ();
 sg13g2_decap_8 FILLER_80_43 ();
 sg13g2_decap_8 FILLER_80_58 ();
 sg13g2_decap_8 FILLER_80_65 ();
 sg13g2_decap_8 FILLER_80_72 ();
 sg13g2_fill_2 FILLER_80_79 ();
 sg13g2_fill_1 FILLER_80_81 ();
 sg13g2_fill_1 FILLER_80_112 ();
 sg13g2_decap_4 FILLER_80_125 ();
 sg13g2_fill_1 FILLER_80_129 ();
 sg13g2_decap_8 FILLER_80_134 ();
 sg13g2_fill_2 FILLER_80_149 ();
 sg13g2_decap_8 FILLER_80_211 ();
 sg13g2_decap_8 FILLER_80_218 ();
 sg13g2_decap_8 FILLER_80_229 ();
 sg13g2_decap_8 FILLER_80_236 ();
 sg13g2_fill_1 FILLER_80_243 ();
 sg13g2_fill_2 FILLER_80_261 ();
 sg13g2_fill_1 FILLER_80_263 ();
 sg13g2_fill_1 FILLER_80_301 ();
 sg13g2_fill_2 FILLER_80_326 ();
 sg13g2_fill_2 FILLER_80_396 ();
 sg13g2_decap_8 FILLER_80_411 ();
 sg13g2_decap_4 FILLER_80_418 ();
 sg13g2_fill_1 FILLER_80_422 ();
 sg13g2_decap_8 FILLER_80_427 ();
 sg13g2_decap_8 FILLER_80_434 ();
 sg13g2_decap_4 FILLER_80_441 ();
 sg13g2_decap_8 FILLER_80_449 ();
 sg13g2_fill_1 FILLER_80_456 ();
 sg13g2_decap_8 FILLER_80_465 ();
 sg13g2_fill_1 FILLER_80_472 ();
 sg13g2_decap_8 FILLER_80_486 ();
 sg13g2_decap_8 FILLER_80_493 ();
 sg13g2_fill_2 FILLER_80_500 ();
 sg13g2_fill_1 FILLER_80_502 ();
 sg13g2_decap_4 FILLER_80_529 ();
 sg13g2_fill_1 FILLER_80_533 ();
 sg13g2_decap_4 FILLER_80_565 ();
 sg13g2_fill_1 FILLER_80_569 ();
 sg13g2_decap_8 FILLER_80_596 ();
 sg13g2_decap_4 FILLER_80_603 ();
 sg13g2_fill_2 FILLER_80_607 ();
 sg13g2_decap_4 FILLER_80_617 ();
 sg13g2_fill_1 FILLER_80_621 ();
 sg13g2_decap_8 FILLER_80_630 ();
 sg13g2_decap_4 FILLER_80_637 ();
 sg13g2_fill_2 FILLER_80_657 ();
 sg13g2_fill_1 FILLER_80_659 ();
 sg13g2_decap_8 FILLER_80_681 ();
 sg13g2_fill_2 FILLER_80_688 ();
 sg13g2_decap_8 FILLER_80_708 ();
 sg13g2_decap_8 FILLER_80_715 ();
 sg13g2_decap_4 FILLER_80_722 ();
 sg13g2_fill_1 FILLER_80_726 ();
 sg13g2_decap_8 FILLER_80_736 ();
 sg13g2_decap_8 FILLER_80_743 ();
 sg13g2_decap_4 FILLER_80_750 ();
 sg13g2_fill_2 FILLER_80_765 ();
 sg13g2_decap_8 FILLER_80_775 ();
 sg13g2_decap_8 FILLER_80_782 ();
 sg13g2_decap_8 FILLER_80_789 ();
 sg13g2_decap_8 FILLER_80_796 ();
 sg13g2_decap_8 FILLER_80_803 ();
 sg13g2_decap_8 FILLER_80_810 ();
 sg13g2_decap_8 FILLER_80_817 ();
 sg13g2_decap_8 FILLER_80_824 ();
 sg13g2_decap_8 FILLER_80_831 ();
 sg13g2_decap_8 FILLER_80_838 ();
 sg13g2_decap_8 FILLER_80_845 ();
 sg13g2_decap_8 FILLER_80_852 ();
 sg13g2_fill_2 FILLER_80_859 ();
 sg13g2_fill_1 FILLER_80_861 ();
 assign uio_oe[0] = net17;
 assign uio_oe[1] = net18;
 assign uio_oe[2] = net19;
 assign uio_oe[3] = net20;
 assign uio_out[0] = net21;
 assign uio_out[1] = net22;
 assign uio_out[2] = net23;
 assign uio_out[3] = net24;
endmodule
